VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_tholin_riscv
  CLASS BLOCK ;
  FOREIGN wrapped_tholin_riscv ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 550.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END custom_settings[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 4.000 506.560 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END io_in[32]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 9.290 546.000 9.570 550.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 170.290 546.000 170.570 550.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 186.390 546.000 186.670 550.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 202.490 546.000 202.770 550.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 218.590 546.000 218.870 550.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 234.690 546.000 234.970 550.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 250.790 546.000 251.070 550.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 546.000 267.170 550.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 546.000 283.270 550.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 546.000 299.370 550.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 546.000 315.470 550.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 25.390 546.000 25.670 550.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 546.000 331.570 550.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 546.000 347.670 550.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 546.000 363.770 550.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 546.000 379.870 550.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 546.000 395.970 550.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 546.000 412.070 550.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 546.000 428.170 550.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 443.990 546.000 444.270 550.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 460.090 546.000 460.370 550.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 476.190 546.000 476.470 550.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 41.490 546.000 41.770 550.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 492.290 546.000 492.570 550.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 508.390 546.000 508.670 550.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 524.490 546.000 524.770 550.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 546.000 540.870 550.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 57.590 546.000 57.870 550.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 73.690 546.000 73.970 550.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 89.790 546.000 90.070 550.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 105.890 546.000 106.170 550.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 121.990 546.000 122.270 550.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 138.090 546.000 138.370 550.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 154.190 546.000 154.470 550.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439350 ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439350 ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 456.870 0.000 457.150 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 489.990 0.000 490.270 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 523.110 0.000 523.390 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END io_out[32]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.778900 ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.227250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END rst_n
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 538.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 538.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.855000 ;
    ANTENNADIFFAREA 0.406350 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 544.180 538.645 ;
      LAYER met1 ;
        RECT 5.130 10.240 544.180 538.800 ;
      LAYER met2 ;
        RECT 5.150 545.720 9.010 546.450 ;
        RECT 9.850 545.720 25.110 546.450 ;
        RECT 25.950 545.720 41.210 546.450 ;
        RECT 42.050 545.720 57.310 546.450 ;
        RECT 58.150 545.720 73.410 546.450 ;
        RECT 74.250 545.720 89.510 546.450 ;
        RECT 90.350 545.720 105.610 546.450 ;
        RECT 106.450 545.720 121.710 546.450 ;
        RECT 122.550 545.720 137.810 546.450 ;
        RECT 138.650 545.720 153.910 546.450 ;
        RECT 154.750 545.720 170.010 546.450 ;
        RECT 170.850 545.720 186.110 546.450 ;
        RECT 186.950 545.720 202.210 546.450 ;
        RECT 203.050 545.720 218.310 546.450 ;
        RECT 219.150 545.720 234.410 546.450 ;
        RECT 235.250 545.720 250.510 546.450 ;
        RECT 251.350 545.720 266.610 546.450 ;
        RECT 267.450 545.720 282.710 546.450 ;
        RECT 283.550 545.720 298.810 546.450 ;
        RECT 299.650 545.720 314.910 546.450 ;
        RECT 315.750 545.720 331.010 546.450 ;
        RECT 331.850 545.720 347.110 546.450 ;
        RECT 347.950 545.720 363.210 546.450 ;
        RECT 364.050 545.720 379.310 546.450 ;
        RECT 380.150 545.720 395.410 546.450 ;
        RECT 396.250 545.720 411.510 546.450 ;
        RECT 412.350 545.720 427.610 546.450 ;
        RECT 428.450 545.720 443.710 546.450 ;
        RECT 444.550 545.720 459.810 546.450 ;
        RECT 460.650 545.720 475.910 546.450 ;
        RECT 476.750 545.720 492.010 546.450 ;
        RECT 492.850 545.720 508.110 546.450 ;
        RECT 508.950 545.720 524.210 546.450 ;
        RECT 525.050 545.720 540.310 546.450 ;
        RECT 5.150 4.280 540.860 545.720 ;
        RECT 5.150 3.670 9.470 4.280 ;
        RECT 10.310 3.670 26.030 4.280 ;
        RECT 26.870 3.670 42.590 4.280 ;
        RECT 43.430 3.670 59.150 4.280 ;
        RECT 59.990 3.670 75.710 4.280 ;
        RECT 76.550 3.670 92.270 4.280 ;
        RECT 93.110 3.670 108.830 4.280 ;
        RECT 109.670 3.670 125.390 4.280 ;
        RECT 126.230 3.670 141.950 4.280 ;
        RECT 142.790 3.670 158.510 4.280 ;
        RECT 159.350 3.670 175.070 4.280 ;
        RECT 175.910 3.670 191.630 4.280 ;
        RECT 192.470 3.670 208.190 4.280 ;
        RECT 209.030 3.670 224.750 4.280 ;
        RECT 225.590 3.670 241.310 4.280 ;
        RECT 242.150 3.670 257.870 4.280 ;
        RECT 258.710 3.670 274.430 4.280 ;
        RECT 275.270 3.670 290.990 4.280 ;
        RECT 291.830 3.670 307.550 4.280 ;
        RECT 308.390 3.670 324.110 4.280 ;
        RECT 324.950 3.670 340.670 4.280 ;
        RECT 341.510 3.670 357.230 4.280 ;
        RECT 358.070 3.670 373.790 4.280 ;
        RECT 374.630 3.670 390.350 4.280 ;
        RECT 391.190 3.670 406.910 4.280 ;
        RECT 407.750 3.670 423.470 4.280 ;
        RECT 424.310 3.670 440.030 4.280 ;
        RECT 440.870 3.670 456.590 4.280 ;
        RECT 457.430 3.670 473.150 4.280 ;
        RECT 473.990 3.670 489.710 4.280 ;
        RECT 490.550 3.670 506.270 4.280 ;
        RECT 507.110 3.670 522.830 4.280 ;
        RECT 523.670 3.670 539.390 4.280 ;
        RECT 540.230 3.670 540.860 4.280 ;
      LAYER met3 ;
        RECT 3.990 520.560 517.895 538.725 ;
        RECT 4.400 519.160 517.895 520.560 ;
        RECT 3.990 506.960 517.895 519.160 ;
        RECT 4.400 505.560 517.895 506.960 ;
        RECT 3.990 493.360 517.895 505.560 ;
        RECT 4.400 491.960 517.895 493.360 ;
        RECT 3.990 479.760 517.895 491.960 ;
        RECT 4.400 478.360 517.895 479.760 ;
        RECT 3.990 466.160 517.895 478.360 ;
        RECT 4.400 464.760 517.895 466.160 ;
        RECT 3.990 452.560 517.895 464.760 ;
        RECT 4.400 451.160 517.895 452.560 ;
        RECT 3.990 438.960 517.895 451.160 ;
        RECT 4.400 437.560 517.895 438.960 ;
        RECT 3.990 425.360 517.895 437.560 ;
        RECT 4.400 423.960 517.895 425.360 ;
        RECT 3.990 411.760 517.895 423.960 ;
        RECT 4.400 410.360 517.895 411.760 ;
        RECT 3.990 398.160 517.895 410.360 ;
        RECT 4.400 396.760 517.895 398.160 ;
        RECT 3.990 384.560 517.895 396.760 ;
        RECT 4.400 383.160 517.895 384.560 ;
        RECT 3.990 370.960 517.895 383.160 ;
        RECT 4.400 369.560 517.895 370.960 ;
        RECT 3.990 357.360 517.895 369.560 ;
        RECT 4.400 355.960 517.895 357.360 ;
        RECT 3.990 343.760 517.895 355.960 ;
        RECT 4.400 342.360 517.895 343.760 ;
        RECT 3.990 330.160 517.895 342.360 ;
        RECT 4.400 328.760 517.895 330.160 ;
        RECT 3.990 316.560 517.895 328.760 ;
        RECT 4.400 315.160 517.895 316.560 ;
        RECT 3.990 302.960 517.895 315.160 ;
        RECT 4.400 301.560 517.895 302.960 ;
        RECT 3.990 289.360 517.895 301.560 ;
        RECT 4.400 287.960 517.895 289.360 ;
        RECT 3.990 275.760 517.895 287.960 ;
        RECT 4.400 274.360 517.895 275.760 ;
        RECT 3.990 262.160 517.895 274.360 ;
        RECT 4.400 260.760 517.895 262.160 ;
        RECT 3.990 248.560 517.895 260.760 ;
        RECT 4.400 247.160 517.895 248.560 ;
        RECT 3.990 234.960 517.895 247.160 ;
        RECT 4.400 233.560 517.895 234.960 ;
        RECT 3.990 221.360 517.895 233.560 ;
        RECT 4.400 219.960 517.895 221.360 ;
        RECT 3.990 207.760 517.895 219.960 ;
        RECT 4.400 206.360 517.895 207.760 ;
        RECT 3.990 194.160 517.895 206.360 ;
        RECT 4.400 192.760 517.895 194.160 ;
        RECT 3.990 180.560 517.895 192.760 ;
        RECT 4.400 179.160 517.895 180.560 ;
        RECT 3.990 166.960 517.895 179.160 ;
        RECT 4.400 165.560 517.895 166.960 ;
        RECT 3.990 153.360 517.895 165.560 ;
        RECT 4.400 151.960 517.895 153.360 ;
        RECT 3.990 139.760 517.895 151.960 ;
        RECT 4.400 138.360 517.895 139.760 ;
        RECT 3.990 126.160 517.895 138.360 ;
        RECT 4.400 124.760 517.895 126.160 ;
        RECT 3.990 112.560 517.895 124.760 ;
        RECT 4.400 111.160 517.895 112.560 ;
        RECT 3.990 98.960 517.895 111.160 ;
        RECT 4.400 97.560 517.895 98.960 ;
        RECT 3.990 85.360 517.895 97.560 ;
        RECT 4.400 83.960 517.895 85.360 ;
        RECT 3.990 71.760 517.895 83.960 ;
        RECT 4.400 70.360 517.895 71.760 ;
        RECT 3.990 58.160 517.895 70.360 ;
        RECT 4.400 56.760 517.895 58.160 ;
        RECT 3.990 44.560 517.895 56.760 ;
        RECT 4.400 43.160 517.895 44.560 ;
        RECT 3.990 30.960 517.895 43.160 ;
        RECT 4.400 29.560 517.895 30.960 ;
        RECT 3.990 10.715 517.895 29.560 ;
      LAYER met4 ;
        RECT 47.215 13.775 97.440 531.585 ;
        RECT 99.840 13.775 174.240 531.585 ;
        RECT 176.640 13.775 251.040 531.585 ;
        RECT 253.440 13.775 327.840 531.585 ;
        RECT 330.240 13.775 404.640 531.585 ;
        RECT 407.040 13.775 481.440 531.585 ;
        RECT 483.840 13.775 487.305 531.585 ;
  END
END wrapped_tholin_riscv
END LIBRARY

