magic
tech sky130A
magscale 1 2
timestamp 1737407066
<< obsli1 >>
rect 1104 2159 108836 107729
<< obsm1 >>
rect 1026 2048 108836 107760
<< metal2 >>
rect 1858 109200 1914 110000
rect 5078 109200 5134 110000
rect 8298 109200 8354 110000
rect 11518 109200 11574 110000
rect 14738 109200 14794 110000
rect 17958 109200 18014 110000
rect 21178 109200 21234 110000
rect 24398 109200 24454 110000
rect 27618 109200 27674 110000
rect 30838 109200 30894 110000
rect 34058 109200 34114 110000
rect 37278 109200 37334 110000
rect 40498 109200 40554 110000
rect 43718 109200 43774 110000
rect 46938 109200 46994 110000
rect 50158 109200 50214 110000
rect 53378 109200 53434 110000
rect 56598 109200 56654 110000
rect 59818 109200 59874 110000
rect 63038 109200 63094 110000
rect 66258 109200 66314 110000
rect 69478 109200 69534 110000
rect 72698 109200 72754 110000
rect 75918 109200 75974 110000
rect 79138 109200 79194 110000
rect 82358 109200 82414 110000
rect 85578 109200 85634 110000
rect 88798 109200 88854 110000
rect 92018 109200 92074 110000
rect 95238 109200 95294 110000
rect 98458 109200 98514 110000
rect 101678 109200 101734 110000
rect 104898 109200 104954 110000
rect 108118 109200 108174 110000
rect 1950 0 2006 800
rect 5262 0 5318 800
rect 8574 0 8630 800
rect 11886 0 11942 800
rect 15198 0 15254 800
rect 18510 0 18566 800
rect 21822 0 21878 800
rect 25134 0 25190 800
rect 28446 0 28502 800
rect 31758 0 31814 800
rect 35070 0 35126 800
rect 38382 0 38438 800
rect 41694 0 41750 800
rect 45006 0 45062 800
rect 48318 0 48374 800
rect 51630 0 51686 800
rect 54942 0 54998 800
rect 58254 0 58310 800
rect 61566 0 61622 800
rect 64878 0 64934 800
rect 68190 0 68246 800
rect 71502 0 71558 800
rect 74814 0 74870 800
rect 78126 0 78182 800
rect 81438 0 81494 800
rect 84750 0 84806 800
rect 88062 0 88118 800
rect 91374 0 91430 800
rect 94686 0 94742 800
rect 97998 0 98054 800
rect 101310 0 101366 800
rect 104622 0 104678 800
rect 107934 0 107990 800
<< obsm2 >>
rect 1030 109144 1802 109290
rect 1970 109144 5022 109290
rect 5190 109144 8242 109290
rect 8410 109144 11462 109290
rect 11630 109144 14682 109290
rect 14850 109144 17902 109290
rect 18070 109144 21122 109290
rect 21290 109144 24342 109290
rect 24510 109144 27562 109290
rect 27730 109144 30782 109290
rect 30950 109144 34002 109290
rect 34170 109144 37222 109290
rect 37390 109144 40442 109290
rect 40610 109144 43662 109290
rect 43830 109144 46882 109290
rect 47050 109144 50102 109290
rect 50270 109144 53322 109290
rect 53490 109144 56542 109290
rect 56710 109144 59762 109290
rect 59930 109144 62982 109290
rect 63150 109144 66202 109290
rect 66370 109144 69422 109290
rect 69590 109144 72642 109290
rect 72810 109144 75862 109290
rect 76030 109144 79082 109290
rect 79250 109144 82302 109290
rect 82470 109144 85522 109290
rect 85690 109144 88742 109290
rect 88910 109144 91962 109290
rect 92130 109144 95182 109290
rect 95350 109144 98402 109290
rect 98570 109144 101622 109290
rect 101790 109144 104842 109290
rect 105010 109144 108062 109290
rect 1030 856 108172 109144
rect 1030 734 1894 856
rect 2062 734 5206 856
rect 5374 734 8518 856
rect 8686 734 11830 856
rect 11998 734 15142 856
rect 15310 734 18454 856
rect 18622 734 21766 856
rect 21934 734 25078 856
rect 25246 734 28390 856
rect 28558 734 31702 856
rect 31870 734 35014 856
rect 35182 734 38326 856
rect 38494 734 41638 856
rect 41806 734 44950 856
rect 45118 734 48262 856
rect 48430 734 51574 856
rect 51742 734 54886 856
rect 55054 734 58198 856
rect 58366 734 61510 856
rect 61678 734 64822 856
rect 64990 734 68134 856
rect 68302 734 71446 856
rect 71614 734 74758 856
rect 74926 734 78070 856
rect 78238 734 81382 856
rect 81550 734 84694 856
rect 84862 734 88006 856
rect 88174 734 91318 856
rect 91486 734 94630 856
rect 94798 734 97942 856
rect 98110 734 101254 856
rect 101422 734 104566 856
rect 104734 734 107878 856
rect 108046 734 108172 856
<< metal3 >>
rect 0 103912 800 104032
rect 0 101192 800 101312
rect 0 98472 800 98592
rect 0 95752 800 95872
rect 0 93032 800 93152
rect 0 90312 800 90432
rect 0 87592 800 87712
rect 0 84872 800 84992
rect 0 82152 800 82272
rect 0 79432 800 79552
rect 0 76712 800 76832
rect 0 73992 800 74112
rect 0 71272 800 71392
rect 0 68552 800 68672
rect 0 65832 800 65952
rect 0 63112 800 63232
rect 0 60392 800 60512
rect 0 57672 800 57792
rect 0 54952 800 55072
rect 0 52232 800 52352
rect 0 49512 800 49632
rect 0 46792 800 46912
rect 0 44072 800 44192
rect 0 41352 800 41472
rect 0 38632 800 38752
rect 0 35912 800 36032
rect 0 33192 800 33312
rect 0 30472 800 30592
rect 0 27752 800 27872
rect 0 25032 800 25152
rect 0 22312 800 22432
rect 0 19592 800 19712
rect 0 16872 800 16992
rect 0 14152 800 14272
rect 0 11432 800 11552
rect 0 8712 800 8832
rect 0 5992 800 6112
<< obsm3 >>
rect 798 104112 103579 107745
rect 880 103832 103579 104112
rect 798 101392 103579 103832
rect 880 101112 103579 101392
rect 798 98672 103579 101112
rect 880 98392 103579 98672
rect 798 95952 103579 98392
rect 880 95672 103579 95952
rect 798 93232 103579 95672
rect 880 92952 103579 93232
rect 798 90512 103579 92952
rect 880 90232 103579 90512
rect 798 87792 103579 90232
rect 880 87512 103579 87792
rect 798 85072 103579 87512
rect 880 84792 103579 85072
rect 798 82352 103579 84792
rect 880 82072 103579 82352
rect 798 79632 103579 82072
rect 880 79352 103579 79632
rect 798 76912 103579 79352
rect 880 76632 103579 76912
rect 798 74192 103579 76632
rect 880 73912 103579 74192
rect 798 71472 103579 73912
rect 880 71192 103579 71472
rect 798 68752 103579 71192
rect 880 68472 103579 68752
rect 798 66032 103579 68472
rect 880 65752 103579 66032
rect 798 63312 103579 65752
rect 880 63032 103579 63312
rect 798 60592 103579 63032
rect 880 60312 103579 60592
rect 798 57872 103579 60312
rect 880 57592 103579 57872
rect 798 55152 103579 57592
rect 880 54872 103579 55152
rect 798 52432 103579 54872
rect 880 52152 103579 52432
rect 798 49712 103579 52152
rect 880 49432 103579 49712
rect 798 46992 103579 49432
rect 880 46712 103579 46992
rect 798 44272 103579 46712
rect 880 43992 103579 44272
rect 798 41552 103579 43992
rect 880 41272 103579 41552
rect 798 38832 103579 41272
rect 880 38552 103579 38832
rect 798 36112 103579 38552
rect 880 35832 103579 36112
rect 798 33392 103579 35832
rect 880 33112 103579 33392
rect 798 30672 103579 33112
rect 880 30392 103579 30672
rect 798 27952 103579 30392
rect 880 27672 103579 27952
rect 798 25232 103579 27672
rect 880 24952 103579 25232
rect 798 22512 103579 24952
rect 880 22232 103579 22512
rect 798 19792 103579 22232
rect 880 19512 103579 19792
rect 798 17072 103579 19512
rect 880 16792 103579 17072
rect 798 14352 103579 16792
rect 880 14072 103579 14352
rect 798 11632 103579 14072
rect 880 11352 103579 11632
rect 798 8912 103579 11352
rect 880 8632 103579 8912
rect 798 6192 103579 8632
rect 880 5912 103579 6192
rect 798 2143 103579 5912
<< metal4 >>
rect 4208 2128 4528 107760
rect 19568 2128 19888 107760
rect 34928 2128 35248 107760
rect 50288 2128 50608 107760
rect 65648 2128 65968 107760
rect 81008 2128 81328 107760
rect 96368 2128 96688 107760
<< obsm4 >>
rect 9443 2755 19488 106317
rect 19968 2755 34848 106317
rect 35328 2755 50208 106317
rect 50688 2755 65568 106317
rect 66048 2755 80928 106317
rect 81408 2755 96288 106317
rect 96768 2755 97461 106317
<< labels >>
rlabel metal3 s 0 11432 800 11552 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 io_in[0]
port 3 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 io_in[10]
port 4 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 io_in[11]
port 5 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 io_in[12]
port 6 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 io_in[13]
port 7 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 io_in[14]
port 8 nsew signal input
rlabel metal3 s 0 57672 800 57792 6 io_in[15]
port 9 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 io_in[16]
port 10 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 io_in[17]
port 11 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 io_in[18]
port 12 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 io_in[19]
port 13 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 io_in[1]
port 14 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 io_in[20]
port 15 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 io_in[21]
port 16 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 io_in[22]
port 17 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 io_in[23]
port 18 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 io_in[24]
port 19 nsew signal input
rlabel metal3 s 0 84872 800 84992 6 io_in[25]
port 20 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 io_in[26]
port 21 nsew signal input
rlabel metal3 s 0 90312 800 90432 6 io_in[27]
port 22 nsew signal input
rlabel metal3 s 0 93032 800 93152 6 io_in[28]
port 23 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 io_in[29]
port 24 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 io_in[2]
port 25 nsew signal input
rlabel metal3 s 0 98472 800 98592 6 io_in[30]
port 26 nsew signal input
rlabel metal3 s 0 101192 800 101312 6 io_in[31]
port 27 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 io_in[32]
port 28 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 io_in[3]
port 29 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 io_in[4]
port 30 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 io_in[5]
port 31 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 io_in[6]
port 32 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 io_in[7]
port 33 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 io_in[8]
port 34 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 io_in[9]
port 35 nsew signal input
rlabel metal2 s 1858 109200 1914 110000 6 io_oeb[0]
port 36 nsew signal output
rlabel metal2 s 34058 109200 34114 110000 6 io_oeb[10]
port 37 nsew signal output
rlabel metal2 s 37278 109200 37334 110000 6 io_oeb[11]
port 38 nsew signal output
rlabel metal2 s 40498 109200 40554 110000 6 io_oeb[12]
port 39 nsew signal output
rlabel metal2 s 43718 109200 43774 110000 6 io_oeb[13]
port 40 nsew signal output
rlabel metal2 s 46938 109200 46994 110000 6 io_oeb[14]
port 41 nsew signal output
rlabel metal2 s 50158 109200 50214 110000 6 io_oeb[15]
port 42 nsew signal output
rlabel metal2 s 53378 109200 53434 110000 6 io_oeb[16]
port 43 nsew signal output
rlabel metal2 s 56598 109200 56654 110000 6 io_oeb[17]
port 44 nsew signal output
rlabel metal2 s 59818 109200 59874 110000 6 io_oeb[18]
port 45 nsew signal output
rlabel metal2 s 63038 109200 63094 110000 6 io_oeb[19]
port 46 nsew signal output
rlabel metal2 s 5078 109200 5134 110000 6 io_oeb[1]
port 47 nsew signal output
rlabel metal2 s 66258 109200 66314 110000 6 io_oeb[20]
port 48 nsew signal output
rlabel metal2 s 69478 109200 69534 110000 6 io_oeb[21]
port 49 nsew signal output
rlabel metal2 s 72698 109200 72754 110000 6 io_oeb[22]
port 50 nsew signal output
rlabel metal2 s 75918 109200 75974 110000 6 io_oeb[23]
port 51 nsew signal output
rlabel metal2 s 79138 109200 79194 110000 6 io_oeb[24]
port 52 nsew signal output
rlabel metal2 s 82358 109200 82414 110000 6 io_oeb[25]
port 53 nsew signal output
rlabel metal2 s 85578 109200 85634 110000 6 io_oeb[26]
port 54 nsew signal output
rlabel metal2 s 88798 109200 88854 110000 6 io_oeb[27]
port 55 nsew signal output
rlabel metal2 s 92018 109200 92074 110000 6 io_oeb[28]
port 56 nsew signal output
rlabel metal2 s 95238 109200 95294 110000 6 io_oeb[29]
port 57 nsew signal output
rlabel metal2 s 8298 109200 8354 110000 6 io_oeb[2]
port 58 nsew signal output
rlabel metal2 s 98458 109200 98514 110000 6 io_oeb[30]
port 59 nsew signal output
rlabel metal2 s 101678 109200 101734 110000 6 io_oeb[31]
port 60 nsew signal output
rlabel metal2 s 104898 109200 104954 110000 6 io_oeb[32]
port 61 nsew signal output
rlabel metal2 s 108118 109200 108174 110000 6 io_oeb[33]
port 62 nsew signal output
rlabel metal2 s 11518 109200 11574 110000 6 io_oeb[3]
port 63 nsew signal output
rlabel metal2 s 14738 109200 14794 110000 6 io_oeb[4]
port 64 nsew signal output
rlabel metal2 s 17958 109200 18014 110000 6 io_oeb[5]
port 65 nsew signal output
rlabel metal2 s 21178 109200 21234 110000 6 io_oeb[6]
port 66 nsew signal output
rlabel metal2 s 24398 109200 24454 110000 6 io_oeb[7]
port 67 nsew signal output
rlabel metal2 s 27618 109200 27674 110000 6 io_oeb[8]
port 68 nsew signal output
rlabel metal2 s 30838 109200 30894 110000 6 io_oeb[9]
port 69 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 io_out[0]
port 70 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 io_out[10]
port 71 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 io_out[11]
port 72 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 io_out[12]
port 73 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 io_out[13]
port 74 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 io_out[14]
port 75 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 io_out[15]
port 76 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 io_out[16]
port 77 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 io_out[17]
port 78 nsew signal output
rlabel metal2 s 61566 0 61622 800 6 io_out[18]
port 79 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 io_out[19]
port 80 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 io_out[1]
port 81 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 io_out[20]
port 82 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 io_out[21]
port 83 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 io_out[22]
port 84 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 io_out[23]
port 85 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 io_out[24]
port 86 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 io_out[25]
port 87 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 io_out[26]
port 88 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 io_out[27]
port 89 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 io_out[28]
port 90 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 io_out[29]
port 91 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 io_out[2]
port 92 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 io_out[30]
port 93 nsew signal output
rlabel metal2 s 104622 0 104678 800 6 io_out[31]
port 94 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 io_out[32]
port 95 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 io_out[3]
port 96 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 io_out[4]
port 97 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 io_out[5]
port 98 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 io_out[6]
port 99 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 io_out[7]
port 100 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 io_out[8]
port 101 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 io_out[9]
port 102 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 rst_n
port 103 nsew signal input
rlabel metal4 s 4208 2128 4528 107760 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 107760 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 107760 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 107760 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 107760 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 107760 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 107760 6 vssd1
port 105 nsew ground bidirectional
rlabel metal3 s 0 5992 800 6112 6 wb_clk_i
port 106 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 110000 110000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 36732996
string GDS_FILE /home/tholin/example_as_sc_hs/openlane/wrapped_tholin_riscv/runs/25_01_20_21_35/results/signoff/wrapped_tholin_riscv.magic.gds
string GDS_START 152790
<< end >>

