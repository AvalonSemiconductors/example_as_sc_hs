magic
tech sky130A
magscale 1 2
timestamp 1736541966
<< obsli1 >>
rect 1104 2159 118864 117521
<< obsm1 >>
rect 842 1980 118864 117552
<< metal2 >>
rect 2226 119200 2282 120000
rect 5722 119200 5778 120000
rect 9218 119200 9274 120000
rect 12714 119200 12770 120000
rect 16210 119200 16266 120000
rect 19706 119200 19762 120000
rect 23202 119200 23258 120000
rect 26698 119200 26754 120000
rect 30194 119200 30250 120000
rect 33690 119200 33746 120000
rect 37186 119200 37242 120000
rect 40682 119200 40738 120000
rect 44178 119200 44234 120000
rect 47674 119200 47730 120000
rect 51170 119200 51226 120000
rect 54666 119200 54722 120000
rect 58162 119200 58218 120000
rect 61658 119200 61714 120000
rect 65154 119200 65210 120000
rect 68650 119200 68706 120000
rect 72146 119200 72202 120000
rect 75642 119200 75698 120000
rect 79138 119200 79194 120000
rect 82634 119200 82690 120000
rect 86130 119200 86186 120000
rect 89626 119200 89682 120000
rect 93122 119200 93178 120000
rect 96618 119200 96674 120000
rect 100114 119200 100170 120000
rect 103610 119200 103666 120000
rect 107106 119200 107162 120000
rect 110602 119200 110658 120000
rect 114098 119200 114154 120000
rect 117594 119200 117650 120000
rect 2502 0 2558 800
rect 6090 0 6146 800
rect 9678 0 9734 800
rect 13266 0 13322 800
rect 16854 0 16910 800
rect 20442 0 20498 800
rect 24030 0 24086 800
rect 27618 0 27674 800
rect 31206 0 31262 800
rect 34794 0 34850 800
rect 38382 0 38438 800
rect 41970 0 42026 800
rect 45558 0 45614 800
rect 49146 0 49202 800
rect 52734 0 52790 800
rect 56322 0 56378 800
rect 59910 0 59966 800
rect 63498 0 63554 800
rect 67086 0 67142 800
rect 70674 0 70730 800
rect 74262 0 74318 800
rect 77850 0 77906 800
rect 81438 0 81494 800
rect 85026 0 85082 800
rect 88614 0 88670 800
rect 92202 0 92258 800
rect 95790 0 95846 800
rect 99378 0 99434 800
rect 102966 0 103022 800
rect 106554 0 106610 800
rect 110142 0 110198 800
rect 113730 0 113786 800
rect 117318 0 117374 800
<< obsm2 >>
rect 848 119144 2170 119354
rect 2338 119144 5666 119354
rect 5834 119144 9162 119354
rect 9330 119144 12658 119354
rect 12826 119144 16154 119354
rect 16322 119144 19650 119354
rect 19818 119144 23146 119354
rect 23314 119144 26642 119354
rect 26810 119144 30138 119354
rect 30306 119144 33634 119354
rect 33802 119144 37130 119354
rect 37298 119144 40626 119354
rect 40794 119144 44122 119354
rect 44290 119144 47618 119354
rect 47786 119144 51114 119354
rect 51282 119144 54610 119354
rect 54778 119144 58106 119354
rect 58274 119144 61602 119354
rect 61770 119144 65098 119354
rect 65266 119144 68594 119354
rect 68762 119144 72090 119354
rect 72258 119144 75586 119354
rect 75754 119144 79082 119354
rect 79250 119144 82578 119354
rect 82746 119144 86074 119354
rect 86242 119144 89570 119354
rect 89738 119144 93066 119354
rect 93234 119144 96562 119354
rect 96730 119144 100058 119354
rect 100226 119144 103554 119354
rect 103722 119144 107050 119354
rect 107218 119144 110546 119354
rect 110714 119144 114042 119354
rect 114210 119144 117538 119354
rect 117706 119144 118292 119354
rect 848 856 118292 119144
rect 848 734 2446 856
rect 2614 734 6034 856
rect 6202 734 9622 856
rect 9790 734 13210 856
rect 13378 734 16798 856
rect 16966 734 20386 856
rect 20554 734 23974 856
rect 24142 734 27562 856
rect 27730 734 31150 856
rect 31318 734 34738 856
rect 34906 734 38326 856
rect 38494 734 41914 856
rect 42082 734 45502 856
rect 45670 734 49090 856
rect 49258 734 52678 856
rect 52846 734 56266 856
rect 56434 734 59854 856
rect 60022 734 63442 856
rect 63610 734 67030 856
rect 67198 734 70618 856
rect 70786 734 74206 856
rect 74374 734 77794 856
rect 77962 734 81382 856
rect 81550 734 84970 856
rect 85138 734 88558 856
rect 88726 734 92146 856
rect 92314 734 95734 856
rect 95902 734 99322 856
rect 99490 734 102910 856
rect 103078 734 106498 856
rect 106666 734 110086 856
rect 110254 734 113674 856
rect 113842 734 117262 856
rect 117430 734 118292 856
<< metal3 >>
rect 0 113704 800 113824
rect 0 110712 800 110832
rect 0 107720 800 107840
rect 0 104728 800 104848
rect 0 101736 800 101856
rect 0 98744 800 98864
rect 0 95752 800 95872
rect 0 92760 800 92880
rect 0 89768 800 89888
rect 0 86776 800 86896
rect 0 83784 800 83904
rect 0 80792 800 80912
rect 0 77800 800 77920
rect 0 74808 800 74928
rect 0 71816 800 71936
rect 0 68824 800 68944
rect 0 65832 800 65952
rect 0 62840 800 62960
rect 0 59848 800 59968
rect 0 56856 800 56976
rect 0 53864 800 53984
rect 0 50872 800 50992
rect 0 47880 800 48000
rect 0 44888 800 45008
rect 0 41896 800 42016
rect 0 38904 800 39024
rect 0 35912 800 36032
rect 0 32920 800 33040
rect 0 29928 800 30048
rect 0 26936 800 27056
rect 0 23944 800 24064
rect 0 20952 800 21072
rect 0 17960 800 18080
rect 0 14968 800 15088
rect 0 11976 800 12096
rect 0 8984 800 9104
rect 0 5992 800 6112
<< obsm3 >>
rect 798 113904 112046 117537
rect 880 113624 112046 113904
rect 798 110912 112046 113624
rect 880 110632 112046 110912
rect 798 107920 112046 110632
rect 880 107640 112046 107920
rect 798 104928 112046 107640
rect 880 104648 112046 104928
rect 798 101936 112046 104648
rect 880 101656 112046 101936
rect 798 98944 112046 101656
rect 880 98664 112046 98944
rect 798 95952 112046 98664
rect 880 95672 112046 95952
rect 798 92960 112046 95672
rect 880 92680 112046 92960
rect 798 89968 112046 92680
rect 880 89688 112046 89968
rect 798 86976 112046 89688
rect 880 86696 112046 86976
rect 798 83984 112046 86696
rect 880 83704 112046 83984
rect 798 80992 112046 83704
rect 880 80712 112046 80992
rect 798 78000 112046 80712
rect 880 77720 112046 78000
rect 798 75008 112046 77720
rect 880 74728 112046 75008
rect 798 72016 112046 74728
rect 880 71736 112046 72016
rect 798 69024 112046 71736
rect 880 68744 112046 69024
rect 798 66032 112046 68744
rect 880 65752 112046 66032
rect 798 63040 112046 65752
rect 880 62760 112046 63040
rect 798 60048 112046 62760
rect 880 59768 112046 60048
rect 798 57056 112046 59768
rect 880 56776 112046 57056
rect 798 54064 112046 56776
rect 880 53784 112046 54064
rect 798 51072 112046 53784
rect 880 50792 112046 51072
rect 798 48080 112046 50792
rect 880 47800 112046 48080
rect 798 45088 112046 47800
rect 880 44808 112046 45088
rect 798 42096 112046 44808
rect 880 41816 112046 42096
rect 798 39104 112046 41816
rect 880 38824 112046 39104
rect 798 36112 112046 38824
rect 880 35832 112046 36112
rect 798 33120 112046 35832
rect 880 32840 112046 33120
rect 798 30128 112046 32840
rect 880 29848 112046 30128
rect 798 27136 112046 29848
rect 880 26856 112046 27136
rect 798 24144 112046 26856
rect 880 23864 112046 24144
rect 798 21152 112046 23864
rect 880 20872 112046 21152
rect 798 18160 112046 20872
rect 880 17880 112046 18160
rect 798 15168 112046 17880
rect 880 14888 112046 15168
rect 798 12176 112046 14888
rect 880 11896 112046 12176
rect 798 9184 112046 11896
rect 880 8904 112046 9184
rect 798 6192 112046 8904
rect 880 5912 112046 6192
rect 798 2143 112046 5912
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
<< obsm4 >>
rect 1715 3979 4128 116789
rect 4608 3979 19488 116789
rect 19968 3979 34848 116789
rect 35328 3979 50208 116789
rect 50688 3979 65568 116789
rect 66048 3979 80928 116789
rect 81408 3979 90285 116789
<< labels >>
rlabel metal3 s 0 11976 800 12096 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 io_in[0]
port 3 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 io_in[10]
port 4 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 io_in[11]
port 5 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 io_in[12]
port 6 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 io_in[13]
port 7 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 io_in[14]
port 8 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 io_in[15]
port 9 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 io_in[16]
port 10 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 io_in[17]
port 11 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 io_in[18]
port 12 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 io_in[19]
port 13 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 io_in[1]
port 14 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 io_in[20]
port 15 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 io_in[21]
port 16 nsew signal input
rlabel metal3 s 0 83784 800 83904 6 io_in[22]
port 17 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 io_in[23]
port 18 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 io_in[24]
port 19 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 io_in[25]
port 20 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 io_in[26]
port 21 nsew signal input
rlabel metal3 s 0 98744 800 98864 6 io_in[27]
port 22 nsew signal input
rlabel metal3 s 0 101736 800 101856 6 io_in[28]
port 23 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 io_in[29]
port 24 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 io_in[2]
port 25 nsew signal input
rlabel metal3 s 0 107720 800 107840 6 io_in[30]
port 26 nsew signal input
rlabel metal3 s 0 110712 800 110832 6 io_in[31]
port 27 nsew signal input
rlabel metal3 s 0 113704 800 113824 6 io_in[32]
port 28 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 io_in[3]
port 29 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 io_in[4]
port 30 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 io_in[5]
port 31 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 io_in[6]
port 32 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 io_in[7]
port 33 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 io_in[8]
port 34 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 io_in[9]
port 35 nsew signal input
rlabel metal2 s 2226 119200 2282 120000 6 io_oeb[0]
port 36 nsew signal output
rlabel metal2 s 37186 119200 37242 120000 6 io_oeb[10]
port 37 nsew signal output
rlabel metal2 s 40682 119200 40738 120000 6 io_oeb[11]
port 38 nsew signal output
rlabel metal2 s 44178 119200 44234 120000 6 io_oeb[12]
port 39 nsew signal output
rlabel metal2 s 47674 119200 47730 120000 6 io_oeb[13]
port 40 nsew signal output
rlabel metal2 s 51170 119200 51226 120000 6 io_oeb[14]
port 41 nsew signal output
rlabel metal2 s 54666 119200 54722 120000 6 io_oeb[15]
port 42 nsew signal output
rlabel metal2 s 58162 119200 58218 120000 6 io_oeb[16]
port 43 nsew signal output
rlabel metal2 s 61658 119200 61714 120000 6 io_oeb[17]
port 44 nsew signal output
rlabel metal2 s 65154 119200 65210 120000 6 io_oeb[18]
port 45 nsew signal output
rlabel metal2 s 68650 119200 68706 120000 6 io_oeb[19]
port 46 nsew signal output
rlabel metal2 s 5722 119200 5778 120000 6 io_oeb[1]
port 47 nsew signal output
rlabel metal2 s 72146 119200 72202 120000 6 io_oeb[20]
port 48 nsew signal output
rlabel metal2 s 75642 119200 75698 120000 6 io_oeb[21]
port 49 nsew signal output
rlabel metal2 s 79138 119200 79194 120000 6 io_oeb[22]
port 50 nsew signal output
rlabel metal2 s 82634 119200 82690 120000 6 io_oeb[23]
port 51 nsew signal output
rlabel metal2 s 86130 119200 86186 120000 6 io_oeb[24]
port 52 nsew signal output
rlabel metal2 s 89626 119200 89682 120000 6 io_oeb[25]
port 53 nsew signal output
rlabel metal2 s 93122 119200 93178 120000 6 io_oeb[26]
port 54 nsew signal output
rlabel metal2 s 96618 119200 96674 120000 6 io_oeb[27]
port 55 nsew signal output
rlabel metal2 s 100114 119200 100170 120000 6 io_oeb[28]
port 56 nsew signal output
rlabel metal2 s 103610 119200 103666 120000 6 io_oeb[29]
port 57 nsew signal output
rlabel metal2 s 9218 119200 9274 120000 6 io_oeb[2]
port 58 nsew signal output
rlabel metal2 s 107106 119200 107162 120000 6 io_oeb[30]
port 59 nsew signal output
rlabel metal2 s 110602 119200 110658 120000 6 io_oeb[31]
port 60 nsew signal output
rlabel metal2 s 114098 119200 114154 120000 6 io_oeb[32]
port 61 nsew signal output
rlabel metal2 s 117594 119200 117650 120000 6 io_oeb[33]
port 62 nsew signal output
rlabel metal2 s 12714 119200 12770 120000 6 io_oeb[3]
port 63 nsew signal output
rlabel metal2 s 16210 119200 16266 120000 6 io_oeb[4]
port 64 nsew signal output
rlabel metal2 s 19706 119200 19762 120000 6 io_oeb[5]
port 65 nsew signal output
rlabel metal2 s 23202 119200 23258 120000 6 io_oeb[6]
port 66 nsew signal output
rlabel metal2 s 26698 119200 26754 120000 6 io_oeb[7]
port 67 nsew signal output
rlabel metal2 s 30194 119200 30250 120000 6 io_oeb[8]
port 68 nsew signal output
rlabel metal2 s 33690 119200 33746 120000 6 io_oeb[9]
port 69 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 io_out[0]
port 70 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 io_out[10]
port 71 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 io_out[11]
port 72 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 io_out[12]
port 73 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 io_out[13]
port 74 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 io_out[14]
port 75 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 io_out[15]
port 76 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 io_out[16]
port 77 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 io_out[17]
port 78 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 io_out[18]
port 79 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 io_out[19]
port 80 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 io_out[1]
port 81 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 io_out[20]
port 82 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 io_out[21]
port 83 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 io_out[22]
port 84 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 io_out[23]
port 85 nsew signal output
rlabel metal2 s 88614 0 88670 800 6 io_out[24]
port 86 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 io_out[25]
port 87 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 io_out[26]
port 88 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 io_out[27]
port 89 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 io_out[28]
port 90 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 io_out[29]
port 91 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 io_out[2]
port 92 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 io_out[30]
port 93 nsew signal output
rlabel metal2 s 113730 0 113786 800 6 io_out[31]
port 94 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 io_out[32]
port 95 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 io_out[3]
port 96 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 io_out[4]
port 97 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 io_out[5]
port 98 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 io_out[6]
port 99 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 io_out[7]
port 100 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 io_out[8]
port 101 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 io_out[9]
port 102 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 rst_n
port 103 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 105 nsew ground bidirectional
rlabel metal3 s 0 5992 800 6112 6 wb_clk_i
port 106 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 38374814
string GDS_FILE /home/tholin/caravel_user_project/openlane/wrapped_tholin_riscv/runs/25_01_10_21_01/results/signoff/wrapped_tholin_riscv.magic.gds
string GDS_START 152726
<< end >>

