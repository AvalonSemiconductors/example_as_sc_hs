VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_tholin_riscv
  CLASS BLOCK ;
  FOREIGN wrapped_tholin_riscv ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 600.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END custom_settings[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213750 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213750 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213750 ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.427500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.427500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END io_in[32]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 11.130 596.000 11.410 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 185.930 596.000 186.210 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 203.410 596.000 203.690 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 220.890 596.000 221.170 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 238.370 596.000 238.650 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 255.850 596.000 256.130 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 273.330 596.000 273.610 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 596.000 291.090 600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 596.000 308.570 600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 596.000 326.050 600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 596.000 343.530 600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 28.610 596.000 28.890 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 596.000 361.010 600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 596.000 378.490 600.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 596.000 395.970 600.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 596.000 413.450 600.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 596.000 430.930 600.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 596.000 448.410 600.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 596.000 465.890 600.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 483.090 596.000 483.370 600.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 500.570 596.000 500.850 600.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 518.050 596.000 518.330 600.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 46.090 596.000 46.370 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 535.530 596.000 535.810 600.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 553.010 596.000 553.290 600.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 570.490 596.000 570.770 600.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 596.000 588.250 600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 63.570 596.000 63.850 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 81.050 596.000 81.330 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 98.530 596.000 98.810 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 116.010 596.000 116.290 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 133.490 596.000 133.770 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 150.970 596.000 151.250 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 168.450 596.000 168.730 600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.433550 ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.433550 ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 532.770 0.000 533.050 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END io_out[32]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.909000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END rst_n
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.855000 ;
    ANTENNADIFFAREA 0.441000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 587.605 ;
      LAYER met1 ;
        RECT 4.210 9.900 594.320 587.760 ;
      LAYER met2 ;
        RECT 4.240 595.720 10.850 596.770 ;
        RECT 11.690 595.720 28.330 596.770 ;
        RECT 29.170 595.720 45.810 596.770 ;
        RECT 46.650 595.720 63.290 596.770 ;
        RECT 64.130 595.720 80.770 596.770 ;
        RECT 81.610 595.720 98.250 596.770 ;
        RECT 99.090 595.720 115.730 596.770 ;
        RECT 116.570 595.720 133.210 596.770 ;
        RECT 134.050 595.720 150.690 596.770 ;
        RECT 151.530 595.720 168.170 596.770 ;
        RECT 169.010 595.720 185.650 596.770 ;
        RECT 186.490 595.720 203.130 596.770 ;
        RECT 203.970 595.720 220.610 596.770 ;
        RECT 221.450 595.720 238.090 596.770 ;
        RECT 238.930 595.720 255.570 596.770 ;
        RECT 256.410 595.720 273.050 596.770 ;
        RECT 273.890 595.720 290.530 596.770 ;
        RECT 291.370 595.720 308.010 596.770 ;
        RECT 308.850 595.720 325.490 596.770 ;
        RECT 326.330 595.720 342.970 596.770 ;
        RECT 343.810 595.720 360.450 596.770 ;
        RECT 361.290 595.720 377.930 596.770 ;
        RECT 378.770 595.720 395.410 596.770 ;
        RECT 396.250 595.720 412.890 596.770 ;
        RECT 413.730 595.720 430.370 596.770 ;
        RECT 431.210 595.720 447.850 596.770 ;
        RECT 448.690 595.720 465.330 596.770 ;
        RECT 466.170 595.720 482.810 596.770 ;
        RECT 483.650 595.720 500.290 596.770 ;
        RECT 501.130 595.720 517.770 596.770 ;
        RECT 518.610 595.720 535.250 596.770 ;
        RECT 536.090 595.720 552.730 596.770 ;
        RECT 553.570 595.720 570.210 596.770 ;
        RECT 571.050 595.720 587.690 596.770 ;
        RECT 588.530 595.720 591.460 596.770 ;
        RECT 4.240 4.280 591.460 595.720 ;
        RECT 4.240 3.670 12.230 4.280 ;
        RECT 13.070 3.670 30.170 4.280 ;
        RECT 31.010 3.670 48.110 4.280 ;
        RECT 48.950 3.670 66.050 4.280 ;
        RECT 66.890 3.670 83.990 4.280 ;
        RECT 84.830 3.670 101.930 4.280 ;
        RECT 102.770 3.670 119.870 4.280 ;
        RECT 120.710 3.670 137.810 4.280 ;
        RECT 138.650 3.670 155.750 4.280 ;
        RECT 156.590 3.670 173.690 4.280 ;
        RECT 174.530 3.670 191.630 4.280 ;
        RECT 192.470 3.670 209.570 4.280 ;
        RECT 210.410 3.670 227.510 4.280 ;
        RECT 228.350 3.670 245.450 4.280 ;
        RECT 246.290 3.670 263.390 4.280 ;
        RECT 264.230 3.670 281.330 4.280 ;
        RECT 282.170 3.670 299.270 4.280 ;
        RECT 300.110 3.670 317.210 4.280 ;
        RECT 318.050 3.670 335.150 4.280 ;
        RECT 335.990 3.670 353.090 4.280 ;
        RECT 353.930 3.670 371.030 4.280 ;
        RECT 371.870 3.670 388.970 4.280 ;
        RECT 389.810 3.670 406.910 4.280 ;
        RECT 407.750 3.670 424.850 4.280 ;
        RECT 425.690 3.670 442.790 4.280 ;
        RECT 443.630 3.670 460.730 4.280 ;
        RECT 461.570 3.670 478.670 4.280 ;
        RECT 479.510 3.670 496.610 4.280 ;
        RECT 497.450 3.670 514.550 4.280 ;
        RECT 515.390 3.670 532.490 4.280 ;
        RECT 533.330 3.670 550.430 4.280 ;
        RECT 551.270 3.670 568.370 4.280 ;
        RECT 569.210 3.670 586.310 4.280 ;
        RECT 587.150 3.670 591.460 4.280 ;
      LAYER met3 ;
        RECT 3.990 569.520 560.230 587.685 ;
        RECT 4.400 568.120 560.230 569.520 ;
        RECT 3.990 554.560 560.230 568.120 ;
        RECT 4.400 553.160 560.230 554.560 ;
        RECT 3.990 539.600 560.230 553.160 ;
        RECT 4.400 538.200 560.230 539.600 ;
        RECT 3.990 524.640 560.230 538.200 ;
        RECT 4.400 523.240 560.230 524.640 ;
        RECT 3.990 509.680 560.230 523.240 ;
        RECT 4.400 508.280 560.230 509.680 ;
        RECT 3.990 494.720 560.230 508.280 ;
        RECT 4.400 493.320 560.230 494.720 ;
        RECT 3.990 479.760 560.230 493.320 ;
        RECT 4.400 478.360 560.230 479.760 ;
        RECT 3.990 464.800 560.230 478.360 ;
        RECT 4.400 463.400 560.230 464.800 ;
        RECT 3.990 449.840 560.230 463.400 ;
        RECT 4.400 448.440 560.230 449.840 ;
        RECT 3.990 434.880 560.230 448.440 ;
        RECT 4.400 433.480 560.230 434.880 ;
        RECT 3.990 419.920 560.230 433.480 ;
        RECT 4.400 418.520 560.230 419.920 ;
        RECT 3.990 404.960 560.230 418.520 ;
        RECT 4.400 403.560 560.230 404.960 ;
        RECT 3.990 390.000 560.230 403.560 ;
        RECT 4.400 388.600 560.230 390.000 ;
        RECT 3.990 375.040 560.230 388.600 ;
        RECT 4.400 373.640 560.230 375.040 ;
        RECT 3.990 360.080 560.230 373.640 ;
        RECT 4.400 358.680 560.230 360.080 ;
        RECT 3.990 345.120 560.230 358.680 ;
        RECT 4.400 343.720 560.230 345.120 ;
        RECT 3.990 330.160 560.230 343.720 ;
        RECT 4.400 328.760 560.230 330.160 ;
        RECT 3.990 315.200 560.230 328.760 ;
        RECT 4.400 313.800 560.230 315.200 ;
        RECT 3.990 300.240 560.230 313.800 ;
        RECT 4.400 298.840 560.230 300.240 ;
        RECT 3.990 285.280 560.230 298.840 ;
        RECT 4.400 283.880 560.230 285.280 ;
        RECT 3.990 270.320 560.230 283.880 ;
        RECT 4.400 268.920 560.230 270.320 ;
        RECT 3.990 255.360 560.230 268.920 ;
        RECT 4.400 253.960 560.230 255.360 ;
        RECT 3.990 240.400 560.230 253.960 ;
        RECT 4.400 239.000 560.230 240.400 ;
        RECT 3.990 225.440 560.230 239.000 ;
        RECT 4.400 224.040 560.230 225.440 ;
        RECT 3.990 210.480 560.230 224.040 ;
        RECT 4.400 209.080 560.230 210.480 ;
        RECT 3.990 195.520 560.230 209.080 ;
        RECT 4.400 194.120 560.230 195.520 ;
        RECT 3.990 180.560 560.230 194.120 ;
        RECT 4.400 179.160 560.230 180.560 ;
        RECT 3.990 165.600 560.230 179.160 ;
        RECT 4.400 164.200 560.230 165.600 ;
        RECT 3.990 150.640 560.230 164.200 ;
        RECT 4.400 149.240 560.230 150.640 ;
        RECT 3.990 135.680 560.230 149.240 ;
        RECT 4.400 134.280 560.230 135.680 ;
        RECT 3.990 120.720 560.230 134.280 ;
        RECT 4.400 119.320 560.230 120.720 ;
        RECT 3.990 105.760 560.230 119.320 ;
        RECT 4.400 104.360 560.230 105.760 ;
        RECT 3.990 90.800 560.230 104.360 ;
        RECT 4.400 89.400 560.230 90.800 ;
        RECT 3.990 75.840 560.230 89.400 ;
        RECT 4.400 74.440 560.230 75.840 ;
        RECT 3.990 60.880 560.230 74.440 ;
        RECT 4.400 59.480 560.230 60.880 ;
        RECT 3.990 45.920 560.230 59.480 ;
        RECT 4.400 44.520 560.230 45.920 ;
        RECT 3.990 30.960 560.230 44.520 ;
        RECT 4.400 29.560 560.230 30.960 ;
        RECT 3.990 10.715 560.230 29.560 ;
      LAYER met4 ;
        RECT 8.575 19.895 20.640 583.945 ;
        RECT 23.040 19.895 97.440 583.945 ;
        RECT 99.840 19.895 174.240 583.945 ;
        RECT 176.640 19.895 251.040 583.945 ;
        RECT 253.440 19.895 327.840 583.945 ;
        RECT 330.240 19.895 404.640 583.945 ;
        RECT 407.040 19.895 451.425 583.945 ;
  END
END wrapped_tholin_riscv
END LIBRARY

