// This is the unpowered netlist.
module wrapped_tholin_riscv (rst_n,
    wb_clk_i,
    custom_settings,
    io_in,
    io_oeb,
    io_out);
 input rst_n;
 input wb_clk_i;
 input [1:0] custom_settings;
 input [32:0] io_in;
 output [33:0] io_oeb;
 output [32:0] io_out;

 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net539;
 wire net535;
 wire net536;
 wire net540;
 wire net541;
 wire net537;
 wire net538;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire _16502_;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire _16552_;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire _16759_;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire _16776_;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire _16801_;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire _16808_;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire _16816_;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire _16840_;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire _16903_;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire _16912_;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire _16922_;
 wire _16923_;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire _16937_;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire _16949_;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire _17061_;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire _17130_;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire _17150_;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire _17160_;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire _17170_;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire _17175_;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire _17292_;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire _17305_;
 wire _17306_;
 wire _17307_;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire _17318_;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire _17354_;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire _17455_;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire _17532_;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire _17541_;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire _17583_;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire _17588_;
 wire _17589_;
 wire _17590_;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire _17595_;
 wire _17596_;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire _17606_;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire _17625_;
 wire _17626_;
 wire _17627_;
 wire _17628_;
 wire _17629_;
 wire _17630_;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire _17634_;
 wire _17635_;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire _17640_;
 wire _17641_;
 wire _17642_;
 wire _17643_;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire _17648_;
 wire _17649_;
 wire _17650_;
 wire _17651_;
 wire _17652_;
 wire _17653_;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire _17657_;
 wire _17658_;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire _17664_;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire _17668_;
 wire _17669_;
 wire _17670_;
 wire _17671_;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire _17675_;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire _17680_;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire _17686_;
 wire _17687_;
 wire _17688_;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire _17694_;
 wire _17695_;
 wire _17696_;
 wire _17697_;
 wire _17698_;
 wire _17699_;
 wire _17700_;
 wire _17701_;
 wire _17702_;
 wire _17703_;
 wire _17704_;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire _17708_;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire _17719_;
 wire _17720_;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire _17724_;
 wire _17725_;
 wire _17726_;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire _17736_;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire _17742_;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire _17748_;
 wire _17749_;
 wire _17750_;
 wire _17751_;
 wire _17752_;
 wire _17753_;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire _17757_;
 wire _17758_;
 wire _17759_;
 wire _17760_;
 wire _17761_;
 wire _17762_;
 wire _17763_;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire _17772_;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire _17778_;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire _17789_;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire _17794_;
 wire _17795_;
 wire _17796_;
 wire _17797_;
 wire _17798_;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire _17813_;
 wire _17814_;
 wire _17815_;
 wire _17816_;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire _17840_;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire _17846_;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire _17867_;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire _17878_;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire _17910_;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire _17922_;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire _17926_;
 wire _17927_;
 wire _17928_;
 wire _17929_;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire _17934_;
 wire _17935_;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire _17939_;
 wire _17940_;
 wire _17941_;
 wire _17942_;
 wire _17943_;
 wire _17944_;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire _17949_;
 wire _17950_;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire _17955_;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire _17961_;
 wire _17962_;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire _17968_;
 wire _17969_;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire _17978_;
 wire _17979_;
 wire _17980_;
 wire _17981_;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire _17988_;
 wire _17989_;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire _17994_;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire _17998_;
 wire _17999_;
 wire _18000_;
 wire _18001_;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire _18011_;
 wire _18012_;
 wire _18013_;
 wire _18014_;
 wire _18015_;
 wire _18016_;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire _18023_;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire _18029_;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire _18035_;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire _18041_;
 wire _18042_;
 wire _18043_;
 wire _18044_;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire _18049_;
 wire _18050_;
 wire _18051_;
 wire _18052_;
 wire _18053_;
 wire _18054_;
 wire _18055_;
 wire _18056_;
 wire _18057_;
 wire _18058_;
 wire _18059_;
 wire _18060_;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire _18066_;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire _18075_;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire _18079_;
 wire _18080_;
 wire _18081_;
 wire _18082_;
 wire _18083_;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire _18091_;
 wire _18092_;
 wire _18093_;
 wire _18094_;
 wire _18095_;
 wire _18096_;
 wire _18097_;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire _18104_;
 wire _18105_;
 wire _18106_;
 wire _18107_;
 wire _18108_;
 wire _18109_;
 wire _18110_;
 wire _18111_;
 wire _18112_;
 wire _18113_;
 wire _18114_;
 wire _18115_;
 wire _18116_;
 wire _18117_;
 wire _18118_;
 wire _18119_;
 wire _18120_;
 wire _18121_;
 wire _18122_;
 wire _18123_;
 wire _18124_;
 wire _18125_;
 wire _18126_;
 wire _18127_;
 wire _18128_;
 wire _18129_;
 wire _18130_;
 wire _18131_;
 wire _18132_;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire _18136_;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire _18140_;
 wire _18141_;
 wire _18142_;
 wire _18143_;
 wire _18144_;
 wire _18145_;
 wire _18146_;
 wire _18147_;
 wire _18148_;
 wire _18149_;
 wire _18150_;
 wire _18151_;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire _18156_;
 wire _18157_;
 wire _18158_;
 wire _18159_;
 wire _18160_;
 wire _18161_;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire _18170_;
 wire _18171_;
 wire _18172_;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire _18176_;
 wire _18177_;
 wire _18178_;
 wire _18179_;
 wire _18180_;
 wire _18181_;
 wire _18182_;
 wire _18183_;
 wire _18184_;
 wire _18185_;
 wire _18186_;
 wire _18187_;
 wire _18188_;
 wire _18189_;
 wire _18190_;
 wire _18191_;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire _18202_;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire _18208_;
 wire _18209_;
 wire _18210_;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire _18217_;
 wire _18218_;
 wire _18219_;
 wire _18220_;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire _18228_;
 wire _18229_;
 wire _18230_;
 wire _18231_;
 wire _18232_;
 wire _18233_;
 wire _18234_;
 wire _18235_;
 wire _18236_;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire _18240_;
 wire _18241_;
 wire _18242_;
 wire _18243_;
 wire _18244_;
 wire _18245_;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire _18250_;
 wire _18251_;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire _18255_;
 wire _18256_;
 wire _18257_;
 wire _18258_;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire _18267_;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire _18288_;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire _18298_;
 wire _18299_;
 wire _18300_;
 wire _18301_;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire _18308_;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire _18315_;
 wire _18316_;
 wire _18317_;
 wire _18318_;
 wire _18319_;
 wire _18320_;
 wire _18321_;
 wire _18322_;
 wire _18323_;
 wire _18324_;
 wire _18325_;
 wire _18326_;
 wire _18327_;
 wire _18328_;
 wire _18329_;
 wire _18330_;
 wire _18331_;
 wire _18332_;
 wire _18333_;
 wire _18334_;
 wire _18335_;
 wire _18336_;
 wire _18337_;
 wire _18338_;
 wire _18339_;
 wire _18340_;
 wire _18341_;
 wire _18342_;
 wire _18343_;
 wire _18344_;
 wire _18345_;
 wire _18346_;
 wire _18347_;
 wire _18348_;
 wire _18349_;
 wire _18350_;
 wire _18351_;
 wire _18352_;
 wire _18353_;
 wire _18354_;
 wire _18355_;
 wire _18356_;
 wire _18357_;
 wire _18358_;
 wire _18359_;
 wire _18360_;
 wire _18361_;
 wire _18362_;
 wire _18363_;
 wire _18364_;
 wire _18365_;
 wire _18366_;
 wire _18367_;
 wire _18368_;
 wire _18369_;
 wire _18370_;
 wire _18371_;
 wire _18372_;
 wire _18373_;
 wire _18374_;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire _18378_;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire _18382_;
 wire _18383_;
 wire _18384_;
 wire _18385_;
 wire _18386_;
 wire _18387_;
 wire _18388_;
 wire _18389_;
 wire _18390_;
 wire _18391_;
 wire _18392_;
 wire _18393_;
 wire _18394_;
 wire _18395_;
 wire _18396_;
 wire _18397_;
 wire _18398_;
 wire _18399_;
 wire _18400_;
 wire _18401_;
 wire _18402_;
 wire _18403_;
 wire _18404_;
 wire _18405_;
 wire _18406_;
 wire _18407_;
 wire _18408_;
 wire _18409_;
 wire _18410_;
 wire _18411_;
 wire _18412_;
 wire _18413_;
 wire _18414_;
 wire _18415_;
 wire _18416_;
 wire _18417_;
 wire _18418_;
 wire _18419_;
 wire _18420_;
 wire _18421_;
 wire _18422_;
 wire _18423_;
 wire _18424_;
 wire _18425_;
 wire _18426_;
 wire _18427_;
 wire _18428_;
 wire _18429_;
 wire _18430_;
 wire _18431_;
 wire _18432_;
 wire _18433_;
 wire _18434_;
 wire _18435_;
 wire _18436_;
 wire _18437_;
 wire _18438_;
 wire _18439_;
 wire _18440_;
 wire _18441_;
 wire _18442_;
 wire _18443_;
 wire _18444_;
 wire _18445_;
 wire _18446_;
 wire _18447_;
 wire _18448_;
 wire _18449_;
 wire _18450_;
 wire _18451_;
 wire _18452_;
 wire _18453_;
 wire _18454_;
 wire _18455_;
 wire _18456_;
 wire _18457_;
 wire _18458_;
 wire _18459_;
 wire _18460_;
 wire _18461_;
 wire _18462_;
 wire _18463_;
 wire _18464_;
 wire _18465_;
 wire _18466_;
 wire _18467_;
 wire _18468_;
 wire _18469_;
 wire _18470_;
 wire _18471_;
 wire _18472_;
 wire _18473_;
 wire _18474_;
 wire _18475_;
 wire _18476_;
 wire _18477_;
 wire _18478_;
 wire _18479_;
 wire _18480_;
 wire _18481_;
 wire _18482_;
 wire _18483_;
 wire _18484_;
 wire _18485_;
 wire _18486_;
 wire _18487_;
 wire _18488_;
 wire _18489_;
 wire _18490_;
 wire _18491_;
 wire _18492_;
 wire _18493_;
 wire _18494_;
 wire _18495_;
 wire _18496_;
 wire _18497_;
 wire _18498_;
 wire _18499_;
 wire _18500_;
 wire _18501_;
 wire _18502_;
 wire _18503_;
 wire _18504_;
 wire _18505_;
 wire _18506_;
 wire _18507_;
 wire _18508_;
 wire _18509_;
 wire _18510_;
 wire _18511_;
 wire _18512_;
 wire _18513_;
 wire _18514_;
 wire _18515_;
 wire _18516_;
 wire _18517_;
 wire _18518_;
 wire _18519_;
 wire _18520_;
 wire _18521_;
 wire _18522_;
 wire _18523_;
 wire _18524_;
 wire _18525_;
 wire _18526_;
 wire _18527_;
 wire _18528_;
 wire _18529_;
 wire _18530_;
 wire _18531_;
 wire _18532_;
 wire _18533_;
 wire _18534_;
 wire _18535_;
 wire _18536_;
 wire _18537_;
 wire _18538_;
 wire _18539_;
 wire _18540_;
 wire _18541_;
 wire _18542_;
 wire _18543_;
 wire _18544_;
 wire _18545_;
 wire _18546_;
 wire _18547_;
 wire _18548_;
 wire _18549_;
 wire _18550_;
 wire _18551_;
 wire _18552_;
 wire _18553_;
 wire _18554_;
 wire _18555_;
 wire _18556_;
 wire _18557_;
 wire _18558_;
 wire _18559_;
 wire _18560_;
 wire _18561_;
 wire _18562_;
 wire _18563_;
 wire _18564_;
 wire _18565_;
 wire _18566_;
 wire _18567_;
 wire _18568_;
 wire _18569_;
 wire _18570_;
 wire _18571_;
 wire _18572_;
 wire _18573_;
 wire _18574_;
 wire _18575_;
 wire _18576_;
 wire _18577_;
 wire _18578_;
 wire _18579_;
 wire _18580_;
 wire _18581_;
 wire _18582_;
 wire _18583_;
 wire _18584_;
 wire _18585_;
 wire _18586_;
 wire _18587_;
 wire _18588_;
 wire _18589_;
 wire _18590_;
 wire _18591_;
 wire _18592_;
 wire _18593_;
 wire _18594_;
 wire _18595_;
 wire _18596_;
 wire _18597_;
 wire _18598_;
 wire _18599_;
 wire _18600_;
 wire _18601_;
 wire _18602_;
 wire _18603_;
 wire _18604_;
 wire _18605_;
 wire _18606_;
 wire _18607_;
 wire _18608_;
 wire _18609_;
 wire _18610_;
 wire _18611_;
 wire _18612_;
 wire _18613_;
 wire _18614_;
 wire _18615_;
 wire _18616_;
 wire _18617_;
 wire _18618_;
 wire _18619_;
 wire _18620_;
 wire _18621_;
 wire _18622_;
 wire _18623_;
 wire _18624_;
 wire _18625_;
 wire _18626_;
 wire _18627_;
 wire _18628_;
 wire _18629_;
 wire _18630_;
 wire _18631_;
 wire _18632_;
 wire _18633_;
 wire _18634_;
 wire _18635_;
 wire _18636_;
 wire _18637_;
 wire _18638_;
 wire _18639_;
 wire _18640_;
 wire _18641_;
 wire _18642_;
 wire _18643_;
 wire _18644_;
 wire _18645_;
 wire _18646_;
 wire _18647_;
 wire _18648_;
 wire _18649_;
 wire _18650_;
 wire _18651_;
 wire _18652_;
 wire _18653_;
 wire _18654_;
 wire _18655_;
 wire _18656_;
 wire _18657_;
 wire _18658_;
 wire _18659_;
 wire _18660_;
 wire _18661_;
 wire _18662_;
 wire _18663_;
 wire _18664_;
 wire _18665_;
 wire _18666_;
 wire _18667_;
 wire _18668_;
 wire _18669_;
 wire _18670_;
 wire _18671_;
 wire _18672_;
 wire _18673_;
 wire _18674_;
 wire _18675_;
 wire _18676_;
 wire _18677_;
 wire _18678_;
 wire _18679_;
 wire _18680_;
 wire _18681_;
 wire _18682_;
 wire _18683_;
 wire _18684_;
 wire _18685_;
 wire _18686_;
 wire _18687_;
 wire _18688_;
 wire _18689_;
 wire _18690_;
 wire _18691_;
 wire _18692_;
 wire _18693_;
 wire _18694_;
 wire _18695_;
 wire _18696_;
 wire _18697_;
 wire _18698_;
 wire _18699_;
 wire _18700_;
 wire _18701_;
 wire _18702_;
 wire _18703_;
 wire _18704_;
 wire _18705_;
 wire _18706_;
 wire _18707_;
 wire _18708_;
 wire _18709_;
 wire _18710_;
 wire _18711_;
 wire _18712_;
 wire _18713_;
 wire _18714_;
 wire _18715_;
 wire _18716_;
 wire _18717_;
 wire _18718_;
 wire _18719_;
 wire _18720_;
 wire _18721_;
 wire _18722_;
 wire _18723_;
 wire _18724_;
 wire _18725_;
 wire _18726_;
 wire _18727_;
 wire _18728_;
 wire _18729_;
 wire _18730_;
 wire _18731_;
 wire _18732_;
 wire _18733_;
 wire _18734_;
 wire _18735_;
 wire _18736_;
 wire _18737_;
 wire _18738_;
 wire _18739_;
 wire _18740_;
 wire _18741_;
 wire _18742_;
 wire _18743_;
 wire _18744_;
 wire _18745_;
 wire _18746_;
 wire _18747_;
 wire _18748_;
 wire _18749_;
 wire _18750_;
 wire _18751_;
 wire _18752_;
 wire _18753_;
 wire _18754_;
 wire _18755_;
 wire _18756_;
 wire _18757_;
 wire _18758_;
 wire _18759_;
 wire _18760_;
 wire _18761_;
 wire _18762_;
 wire _18763_;
 wire _18764_;
 wire _18765_;
 wire _18766_;
 wire _18767_;
 wire _18768_;
 wire _18769_;
 wire _18770_;
 wire _18771_;
 wire _18772_;
 wire _18773_;
 wire _18774_;
 wire _18775_;
 wire _18776_;
 wire _18777_;
 wire _18778_;
 wire _18779_;
 wire _18780_;
 wire _18781_;
 wire _18782_;
 wire _18783_;
 wire _18784_;
 wire _18785_;
 wire _18786_;
 wire _18787_;
 wire _18788_;
 wire _18789_;
 wire _18790_;
 wire _18791_;
 wire _18792_;
 wire _18793_;
 wire _18794_;
 wire _18795_;
 wire _18796_;
 wire _18797_;
 wire _18798_;
 wire _18799_;
 wire _18800_;
 wire _18801_;
 wire _18802_;
 wire _18803_;
 wire _18804_;
 wire _18805_;
 wire _18806_;
 wire _18807_;
 wire _18808_;
 wire _18809_;
 wire _18810_;
 wire _18811_;
 wire _18812_;
 wire _18813_;
 wire _18814_;
 wire _18815_;
 wire _18816_;
 wire _18817_;
 wire _18818_;
 wire _18819_;
 wire _18820_;
 wire _18821_;
 wire _18822_;
 wire _18823_;
 wire _18824_;
 wire _18825_;
 wire _18826_;
 wire _18827_;
 wire _18828_;
 wire _18829_;
 wire _18830_;
 wire _18831_;
 wire _18832_;
 wire _18833_;
 wire _18834_;
 wire _18835_;
 wire _18836_;
 wire _18837_;
 wire _18838_;
 wire _18839_;
 wire _18840_;
 wire _18841_;
 wire _18842_;
 wire _18843_;
 wire _18844_;
 wire _18845_;
 wire _18846_;
 wire _18847_;
 wire _18848_;
 wire _18849_;
 wire _18850_;
 wire _18851_;
 wire _18852_;
 wire _18853_;
 wire _18854_;
 wire _18855_;
 wire _18856_;
 wire _18857_;
 wire _18858_;
 wire _18859_;
 wire _18860_;
 wire _18861_;
 wire _18862_;
 wire _18863_;
 wire _18864_;
 wire _18865_;
 wire _18866_;
 wire _18867_;
 wire _18868_;
 wire _18869_;
 wire _18870_;
 wire _18871_;
 wire _18872_;
 wire _18873_;
 wire _18874_;
 wire _18875_;
 wire _18876_;
 wire _18877_;
 wire _18878_;
 wire _18879_;
 wire _18880_;
 wire _18881_;
 wire _18882_;
 wire _18883_;
 wire _18884_;
 wire _18885_;
 wire _18886_;
 wire _18887_;
 wire _18888_;
 wire _18889_;
 wire _18890_;
 wire _18891_;
 wire _18892_;
 wire _18893_;
 wire _18894_;
 wire _18895_;
 wire _18896_;
 wire _18897_;
 wire _18898_;
 wire _18899_;
 wire _18900_;
 wire _18901_;
 wire _18902_;
 wire _18903_;
 wire _18904_;
 wire _18905_;
 wire _18906_;
 wire _18907_;
 wire _18908_;
 wire _18909_;
 wire _18910_;
 wire _18911_;
 wire _18912_;
 wire _18913_;
 wire _18914_;
 wire _18915_;
 wire _18916_;
 wire _18917_;
 wire _18918_;
 wire _18919_;
 wire _18920_;
 wire _18921_;
 wire _18922_;
 wire _18923_;
 wire _18924_;
 wire _18925_;
 wire _18926_;
 wire _18927_;
 wire _18928_;
 wire _18929_;
 wire _18930_;
 wire _18931_;
 wire _18932_;
 wire _18933_;
 wire _18934_;
 wire _18935_;
 wire _18936_;
 wire _18937_;
 wire _18938_;
 wire _18939_;
 wire _18940_;
 wire _18941_;
 wire _18942_;
 wire _18943_;
 wire _18944_;
 wire _18945_;
 wire _18946_;
 wire _18947_;
 wire _18948_;
 wire _18949_;
 wire _18950_;
 wire _18951_;
 wire _18952_;
 wire _18953_;
 wire _18954_;
 wire _18955_;
 wire _18956_;
 wire _18957_;
 wire _18958_;
 wire _18959_;
 wire _18960_;
 wire _18961_;
 wire _18962_;
 wire _18963_;
 wire _18964_;
 wire _18965_;
 wire _18966_;
 wire _18967_;
 wire _18968_;
 wire _18969_;
 wire _18970_;
 wire _18971_;
 wire _18972_;
 wire _18973_;
 wire _18974_;
 wire _18975_;
 wire _18976_;
 wire _18977_;
 wire _18978_;
 wire _18979_;
 wire _18980_;
 wire _18981_;
 wire _18982_;
 wire _18983_;
 wire _18984_;
 wire _18985_;
 wire _18986_;
 wire _18987_;
 wire _18988_;
 wire _18989_;
 wire _18990_;
 wire _18991_;
 wire _18992_;
 wire _18993_;
 wire _18994_;
 wire _18995_;
 wire _18996_;
 wire _18997_;
 wire _18998_;
 wire _18999_;
 wire _19000_;
 wire _19001_;
 wire _19002_;
 wire _19003_;
 wire _19004_;
 wire _19005_;
 wire _19006_;
 wire _19007_;
 wire _19008_;
 wire _19009_;
 wire _19010_;
 wire _19011_;
 wire _19012_;
 wire _19013_;
 wire _19014_;
 wire _19015_;
 wire _19016_;
 wire _19017_;
 wire _19018_;
 wire _19019_;
 wire _19020_;
 wire _19021_;
 wire _19022_;
 wire _19023_;
 wire _19024_;
 wire _19025_;
 wire _19026_;
 wire _19027_;
 wire _19028_;
 wire _19029_;
 wire _19030_;
 wire _19031_;
 wire _19032_;
 wire _19033_;
 wire _19034_;
 wire _19035_;
 wire _19036_;
 wire _19037_;
 wire _19038_;
 wire _19039_;
 wire _19040_;
 wire _19041_;
 wire _19042_;
 wire _19043_;
 wire _19044_;
 wire _19045_;
 wire _19046_;
 wire _19047_;
 wire _19048_;
 wire _19049_;
 wire _19050_;
 wire _19051_;
 wire _19052_;
 wire _19053_;
 wire _19054_;
 wire _19055_;
 wire _19056_;
 wire _19057_;
 wire _19058_;
 wire _19059_;
 wire _19060_;
 wire _19061_;
 wire _19062_;
 wire _19063_;
 wire _19064_;
 wire _19065_;
 wire _19066_;
 wire _19067_;
 wire _19068_;
 wire _19069_;
 wire _19070_;
 wire _19071_;
 wire _19072_;
 wire _19073_;
 wire _19074_;
 wire _19075_;
 wire _19076_;
 wire _19077_;
 wire _19078_;
 wire _19079_;
 wire _19080_;
 wire _19081_;
 wire _19082_;
 wire _19083_;
 wire _19084_;
 wire _19085_;
 wire _19086_;
 wire _19087_;
 wire _19088_;
 wire _19089_;
 wire _19090_;
 wire _19091_;
 wire _19092_;
 wire _19093_;
 wire _19094_;
 wire _19095_;
 wire _19096_;
 wire _19097_;
 wire _19098_;
 wire _19099_;
 wire _19100_;
 wire _19101_;
 wire _19102_;
 wire _19103_;
 wire _19104_;
 wire _19105_;
 wire _19106_;
 wire _19107_;
 wire _19108_;
 wire _19109_;
 wire _19110_;
 wire _19111_;
 wire _19112_;
 wire _19113_;
 wire _19114_;
 wire _19115_;
 wire _19116_;
 wire _19117_;
 wire _19118_;
 wire _19119_;
 wire _19120_;
 wire _19121_;
 wire _19122_;
 wire _19123_;
 wire _19124_;
 wire _19125_;
 wire _19126_;
 wire _19127_;
 wire _19128_;
 wire _19129_;
 wire _19130_;
 wire _19131_;
 wire _19132_;
 wire _19133_;
 wire _19134_;
 wire _19135_;
 wire _19136_;
 wire _19137_;
 wire _19138_;
 wire _19139_;
 wire _19140_;
 wire _19141_;
 wire _19142_;
 wire _19143_;
 wire _19144_;
 wire _19145_;
 wire _19146_;
 wire _19147_;
 wire _19148_;
 wire _19149_;
 wire _19150_;
 wire _19151_;
 wire _19152_;
 wire _19153_;
 wire _19154_;
 wire _19155_;
 wire _19156_;
 wire _19157_;
 wire _19158_;
 wire _19159_;
 wire _19160_;
 wire _19161_;
 wire _19162_;
 wire _19163_;
 wire _19164_;
 wire _19165_;
 wire _19166_;
 wire _19167_;
 wire _19168_;
 wire _19169_;
 wire _19170_;
 wire _19171_;
 wire _19172_;
 wire _19173_;
 wire _19174_;
 wire _19175_;
 wire _19176_;
 wire _19177_;
 wire _19178_;
 wire _19179_;
 wire _19180_;
 wire _19181_;
 wire _19182_;
 wire _19183_;
 wire _19184_;
 wire _19185_;
 wire _19186_;
 wire _19187_;
 wire _19188_;
 wire _19189_;
 wire _19190_;
 wire _19191_;
 wire _19192_;
 wire _19193_;
 wire _19194_;
 wire _19195_;
 wire _19196_;
 wire _19197_;
 wire _19198_;
 wire _19199_;
 wire _19200_;
 wire _19201_;
 wire _19202_;
 wire _19203_;
 wire _19204_;
 wire _19205_;
 wire _19206_;
 wire _19207_;
 wire _19208_;
 wire _19209_;
 wire _19210_;
 wire _19211_;
 wire _19212_;
 wire _19213_;
 wire _19214_;
 wire _19215_;
 wire _19216_;
 wire _19217_;
 wire _19218_;
 wire _19219_;
 wire _19220_;
 wire _19221_;
 wire _19222_;
 wire _19223_;
 wire _19224_;
 wire _19225_;
 wire _19226_;
 wire _19227_;
 wire _19228_;
 wire _19229_;
 wire _19230_;
 wire _19231_;
 wire _19232_;
 wire _19233_;
 wire _19234_;
 wire _19235_;
 wire _19236_;
 wire _19237_;
 wire _19238_;
 wire _19239_;
 wire _19240_;
 wire _19241_;
 wire _19242_;
 wire _19243_;
 wire _19244_;
 wire _19245_;
 wire _19246_;
 wire _19247_;
 wire _19248_;
 wire _19249_;
 wire _19250_;
 wire _19251_;
 wire _19252_;
 wire _19253_;
 wire _19254_;
 wire _19255_;
 wire _19256_;
 wire _19257_;
 wire _19258_;
 wire _19259_;
 wire _19260_;
 wire _19261_;
 wire _19262_;
 wire _19263_;
 wire _19264_;
 wire _19265_;
 wire _19266_;
 wire _19267_;
 wire _19268_;
 wire _19269_;
 wire _19270_;
 wire _19271_;
 wire _19272_;
 wire _19273_;
 wire _19274_;
 wire _19275_;
 wire _19276_;
 wire _19277_;
 wire _19278_;
 wire _19279_;
 wire _19280_;
 wire _19281_;
 wire _19282_;
 wire _19283_;
 wire _19284_;
 wire _19285_;
 wire _19286_;
 wire _19287_;
 wire _19288_;
 wire _19289_;
 wire _19290_;
 wire _19291_;
 wire _19292_;
 wire _19293_;
 wire _19294_;
 wire _19295_;
 wire _19296_;
 wire _19297_;
 wire _19298_;
 wire _19299_;
 wire _19300_;
 wire _19301_;
 wire _19302_;
 wire _19303_;
 wire _19304_;
 wire _19305_;
 wire _19306_;
 wire _19307_;
 wire _19308_;
 wire _19309_;
 wire _19310_;
 wire _19311_;
 wire _19312_;
 wire _19313_;
 wire _19314_;
 wire _19315_;
 wire _19316_;
 wire _19317_;
 wire _19318_;
 wire _19319_;
 wire _19320_;
 wire _19321_;
 wire _19322_;
 wire _19323_;
 wire _19324_;
 wire _19325_;
 wire _19326_;
 wire _19327_;
 wire _19328_;
 wire _19329_;
 wire _19330_;
 wire _19331_;
 wire _19332_;
 wire _19333_;
 wire _19334_;
 wire _19335_;
 wire _19336_;
 wire _19337_;
 wire _19338_;
 wire _19339_;
 wire _19340_;
 wire _19341_;
 wire _19342_;
 wire _19343_;
 wire _19344_;
 wire _19345_;
 wire _19346_;
 wire _19347_;
 wire _19348_;
 wire _19349_;
 wire _19350_;
 wire _19351_;
 wire _19352_;
 wire _19353_;
 wire _19354_;
 wire _19355_;
 wire _19356_;
 wire _19357_;
 wire _19358_;
 wire _19359_;
 wire _19360_;
 wire _19361_;
 wire _19362_;
 wire _19363_;
 wire _19364_;
 wire _19365_;
 wire _19366_;
 wire _19367_;
 wire _19368_;
 wire _19369_;
 wire _19370_;
 wire _19371_;
 wire _19372_;
 wire _19373_;
 wire _19374_;
 wire _19375_;
 wire _19376_;
 wire _19377_;
 wire _19378_;
 wire _19379_;
 wire _19380_;
 wire _19381_;
 wire _19382_;
 wire _19383_;
 wire _19384_;
 wire _19385_;
 wire _19386_;
 wire _19387_;
 wire _19388_;
 wire _19389_;
 wire _19390_;
 wire _19391_;
 wire _19392_;
 wire _19393_;
 wire _19394_;
 wire _19395_;
 wire _19396_;
 wire _19397_;
 wire _19398_;
 wire _19399_;
 wire _19400_;
 wire _19401_;
 wire _19402_;
 wire _19403_;
 wire _19404_;
 wire _19405_;
 wire _19406_;
 wire _19407_;
 wire _19408_;
 wire _19409_;
 wire _19410_;
 wire _19411_;
 wire _19412_;
 wire _19413_;
 wire _19414_;
 wire _19415_;
 wire _19416_;
 wire _19417_;
 wire _19418_;
 wire _19419_;
 wire _19420_;
 wire _19421_;
 wire _19422_;
 wire _19423_;
 wire _19424_;
 wire _19425_;
 wire _19426_;
 wire _19427_;
 wire _19428_;
 wire _19429_;
 wire _19430_;
 wire _19431_;
 wire _19432_;
 wire _19433_;
 wire _19434_;
 wire _19435_;
 wire _19436_;
 wire _19437_;
 wire _19438_;
 wire _19439_;
 wire _19440_;
 wire _19441_;
 wire _19442_;
 wire _19443_;
 wire _19444_;
 wire _19445_;
 wire _19446_;
 wire _19447_;
 wire _19448_;
 wire _19449_;
 wire _19450_;
 wire _19451_;
 wire _19452_;
 wire _19453_;
 wire _19454_;
 wire _19455_;
 wire _19456_;
 wire _19457_;
 wire _19458_;
 wire _19459_;
 wire _19460_;
 wire _19461_;
 wire _19462_;
 wire _19463_;
 wire _19464_;
 wire _19465_;
 wire _19466_;
 wire _19467_;
 wire _19468_;
 wire _19469_;
 wire _19470_;
 wire _19471_;
 wire _19472_;
 wire _19473_;
 wire _19474_;
 wire _19475_;
 wire _19476_;
 wire _19477_;
 wire _19478_;
 wire _19479_;
 wire _19480_;
 wire _19481_;
 wire _19482_;
 wire _19483_;
 wire _19484_;
 wire _19485_;
 wire _19486_;
 wire _19487_;
 wire _19488_;
 wire _19489_;
 wire _19490_;
 wire _19491_;
 wire _19492_;
 wire _19493_;
 wire _19494_;
 wire _19495_;
 wire _19496_;
 wire _19497_;
 wire _19498_;
 wire _19499_;
 wire _19500_;
 wire _19501_;
 wire _19502_;
 wire _19503_;
 wire _19504_;
 wire _19505_;
 wire _19506_;
 wire _19507_;
 wire _19508_;
 wire _19509_;
 wire _19510_;
 wire _19511_;
 wire _19512_;
 wire _19513_;
 wire _19514_;
 wire _19515_;
 wire _19516_;
 wire _19517_;
 wire _19518_;
 wire _19519_;
 wire _19520_;
 wire _19521_;
 wire _19522_;
 wire _19523_;
 wire _19524_;
 wire _19525_;
 wire _19526_;
 wire _19527_;
 wire _19528_;
 wire _19529_;
 wire _19530_;
 wire _19531_;
 wire _19532_;
 wire _19533_;
 wire _19534_;
 wire _19535_;
 wire _19536_;
 wire _19537_;
 wire _19538_;
 wire _19539_;
 wire _19540_;
 wire _19541_;
 wire _19542_;
 wire _19543_;
 wire _19544_;
 wire _19545_;
 wire _19546_;
 wire _19547_;
 wire _19548_;
 wire _19549_;
 wire _19550_;
 wire _19551_;
 wire _19552_;
 wire _19553_;
 wire _19554_;
 wire _19555_;
 wire _19556_;
 wire _19557_;
 wire _19558_;
 wire _19559_;
 wire _19560_;
 wire _19561_;
 wire _19562_;
 wire _19563_;
 wire _19564_;
 wire _19565_;
 wire _19566_;
 wire _19567_;
 wire _19568_;
 wire _19569_;
 wire _19570_;
 wire _19571_;
 wire _19572_;
 wire _19573_;
 wire _19574_;
 wire _19575_;
 wire _19576_;
 wire _19577_;
 wire _19578_;
 wire _19579_;
 wire _19580_;
 wire _19581_;
 wire _19582_;
 wire _19583_;
 wire _19584_;
 wire _19585_;
 wire _19586_;
 wire _19587_;
 wire _19588_;
 wire _19589_;
 wire _19590_;
 wire _19591_;
 wire _19592_;
 wire _19593_;
 wire _19594_;
 wire _19595_;
 wire _19596_;
 wire _19597_;
 wire _19598_;
 wire _19599_;
 wire _19600_;
 wire _19601_;
 wire _19602_;
 wire _19603_;
 wire _19604_;
 wire _19605_;
 wire _19606_;
 wire _19607_;
 wire _19608_;
 wire _19609_;
 wire _19610_;
 wire _19611_;
 wire _19612_;
 wire _19613_;
 wire _19614_;
 wire _19615_;
 wire _19616_;
 wire _19617_;
 wire _19618_;
 wire _19619_;
 wire _19620_;
 wire _19621_;
 wire _19622_;
 wire _19623_;
 wire _19624_;
 wire _19625_;
 wire _19626_;
 wire _19627_;
 wire _19628_;
 wire _19629_;
 wire _19630_;
 wire _19631_;
 wire _19632_;
 wire _19633_;
 wire _19634_;
 wire _19635_;
 wire _19636_;
 wire _19637_;
 wire _19638_;
 wire _19639_;
 wire _19640_;
 wire _19641_;
 wire _19642_;
 wire _19643_;
 wire _19644_;
 wire _19645_;
 wire _19646_;
 wire _19647_;
 wire _19648_;
 wire _19649_;
 wire _19650_;
 wire _19651_;
 wire _19652_;
 wire _19653_;
 wire _19654_;
 wire _19655_;
 wire _19656_;
 wire _19657_;
 wire _19658_;
 wire _19659_;
 wire _19660_;
 wire _19661_;
 wire _19662_;
 wire _19663_;
 wire _19664_;
 wire _19665_;
 wire _19666_;
 wire _19667_;
 wire _19668_;
 wire _19669_;
 wire _19670_;
 wire _19671_;
 wire _19672_;
 wire _19673_;
 wire _19674_;
 wire _19675_;
 wire _19676_;
 wire _19677_;
 wire _19678_;
 wire _19679_;
 wire _19680_;
 wire _19681_;
 wire _19682_;
 wire _19683_;
 wire _19684_;
 wire _19685_;
 wire _19686_;
 wire _19687_;
 wire _19688_;
 wire _19689_;
 wire _19690_;
 wire _19691_;
 wire _19692_;
 wire _19693_;
 wire _19694_;
 wire _19695_;
 wire _19696_;
 wire _19697_;
 wire _19698_;
 wire _19699_;
 wire _19700_;
 wire _19701_;
 wire _19702_;
 wire _19703_;
 wire _19704_;
 wire _19705_;
 wire _19706_;
 wire _19707_;
 wire _19708_;
 wire _19709_;
 wire _19710_;
 wire _19711_;
 wire _19712_;
 wire _19713_;
 wire _19714_;
 wire _19715_;
 wire _19716_;
 wire _19717_;
 wire _19718_;
 wire _19719_;
 wire _19720_;
 wire _19721_;
 wire _19722_;
 wire _19723_;
 wire _19724_;
 wire _19725_;
 wire _19726_;
 wire _19727_;
 wire _19728_;
 wire _19729_;
 wire _19730_;
 wire _19731_;
 wire _19732_;
 wire _19733_;
 wire _19734_;
 wire _19735_;
 wire _19736_;
 wire _19737_;
 wire _19738_;
 wire _19739_;
 wire _19740_;
 wire _19741_;
 wire _19742_;
 wire _19743_;
 wire _19744_;
 wire _19745_;
 wire _19746_;
 wire _19747_;
 wire _19748_;
 wire _19749_;
 wire _19750_;
 wire _19751_;
 wire _19752_;
 wire _19753_;
 wire _19754_;
 wire _19755_;
 wire _19756_;
 wire _19757_;
 wire _19758_;
 wire _19759_;
 wire _19760_;
 wire _19761_;
 wire _19762_;
 wire _19763_;
 wire _19764_;
 wire _19765_;
 wire _19766_;
 wire _19767_;
 wire _19768_;
 wire _19769_;
 wire _19770_;
 wire _19771_;
 wire _19772_;
 wire _19773_;
 wire _19774_;
 wire _19775_;
 wire _19776_;
 wire _19777_;
 wire _19778_;
 wire _19779_;
 wire _19780_;
 wire _19781_;
 wire _19782_;
 wire _19783_;
 wire _19784_;
 wire _19785_;
 wire _19786_;
 wire _19787_;
 wire _19788_;
 wire _19789_;
 wire _19790_;
 wire _19791_;
 wire _19792_;
 wire _19793_;
 wire _19794_;
 wire _19795_;
 wire _19796_;
 wire _19797_;
 wire _19798_;
 wire _19799_;
 wire _19800_;
 wire _19801_;
 wire _19802_;
 wire _19803_;
 wire _19804_;
 wire _19805_;
 wire _19806_;
 wire _19807_;
 wire _19808_;
 wire _19809_;
 wire _19810_;
 wire _19811_;
 wire _19812_;
 wire _19813_;
 wire _19814_;
 wire _19815_;
 wire _19816_;
 wire _19817_;
 wire _19818_;
 wire _19819_;
 wire _19820_;
 wire _19821_;
 wire _19822_;
 wire _19823_;
 wire _19824_;
 wire _19825_;
 wire _19826_;
 wire _19827_;
 wire _19828_;
 wire _19829_;
 wire _19830_;
 wire _19831_;
 wire _19832_;
 wire _19833_;
 wire _19834_;
 wire _19835_;
 wire _19836_;
 wire _19837_;
 wire _19838_;
 wire _19839_;
 wire _19840_;
 wire _19841_;
 wire _19842_;
 wire _19843_;
 wire _19844_;
 wire _19845_;
 wire _19846_;
 wire _19847_;
 wire _19848_;
 wire _19849_;
 wire _19850_;
 wire _19851_;
 wire _19852_;
 wire _19853_;
 wire _19854_;
 wire _19855_;
 wire _19856_;
 wire _19857_;
 wire _19858_;
 wire _19859_;
 wire _19860_;
 wire _19861_;
 wire _19862_;
 wire _19863_;
 wire _19864_;
 wire _19865_;
 wire _19866_;
 wire _19867_;
 wire _19868_;
 wire _19869_;
 wire _19870_;
 wire _19871_;
 wire _19872_;
 wire _19873_;
 wire _19874_;
 wire _19875_;
 wire _19876_;
 wire _19877_;
 wire _19878_;
 wire _19879_;
 wire _19880_;
 wire _19881_;
 wire _19882_;
 wire _19883_;
 wire _19884_;
 wire _19885_;
 wire _19886_;
 wire _19887_;
 wire _19888_;
 wire _19889_;
 wire _19890_;
 wire _19891_;
 wire _19892_;
 wire _19893_;
 wire _19894_;
 wire _19895_;
 wire _19896_;
 wire _19897_;
 wire _19898_;
 wire _19899_;
 wire _19900_;
 wire _19901_;
 wire _19902_;
 wire _19903_;
 wire _19904_;
 wire _19905_;
 wire _19906_;
 wire _19907_;
 wire _19908_;
 wire _19909_;
 wire _19910_;
 wire _19911_;
 wire _19912_;
 wire _19913_;
 wire _19914_;
 wire _19915_;
 wire _19916_;
 wire _19917_;
 wire _19918_;
 wire _19919_;
 wire _19920_;
 wire _19921_;
 wire _19922_;
 wire _19923_;
 wire _19924_;
 wire _19925_;
 wire _19926_;
 wire _19927_;
 wire _19928_;
 wire _19929_;
 wire _19930_;
 wire _19931_;
 wire _19932_;
 wire _19933_;
 wire _19934_;
 wire _19935_;
 wire _19936_;
 wire _19937_;
 wire _19938_;
 wire _19939_;
 wire _19940_;
 wire _19941_;
 wire _19942_;
 wire _19943_;
 wire _19944_;
 wire _19945_;
 wire _19946_;
 wire _19947_;
 wire _19948_;
 wire _19949_;
 wire _19950_;
 wire _19951_;
 wire _19952_;
 wire _19953_;
 wire _19954_;
 wire _19955_;
 wire _19956_;
 wire _19957_;
 wire _19958_;
 wire _19959_;
 wire _19960_;
 wire _19961_;
 wire _19962_;
 wire _19963_;
 wire _19964_;
 wire _19965_;
 wire _19966_;
 wire _19967_;
 wire _19968_;
 wire _19969_;
 wire _19970_;
 wire _19971_;
 wire _19972_;
 wire _19973_;
 wire _19974_;
 wire _19975_;
 wire _19976_;
 wire _19977_;
 wire _19978_;
 wire _19979_;
 wire _19980_;
 wire _19981_;
 wire _19982_;
 wire _19983_;
 wire _19984_;
 wire _19985_;
 wire _19986_;
 wire _19987_;
 wire _19988_;
 wire _19989_;
 wire _19990_;
 wire _19991_;
 wire _19992_;
 wire _19993_;
 wire _19994_;
 wire _19995_;
 wire _19996_;
 wire _19997_;
 wire _19998_;
 wire _19999_;
 wire _20000_;
 wire _20001_;
 wire _20002_;
 wire _20003_;
 wire _20004_;
 wire _20005_;
 wire _20006_;
 wire _20007_;
 wire _20008_;
 wire _20009_;
 wire _20010_;
 wire _20011_;
 wire _20012_;
 wire _20013_;
 wire _20014_;
 wire _20015_;
 wire _20016_;
 wire _20017_;
 wire _20018_;
 wire _20019_;
 wire _20020_;
 wire _20021_;
 wire _20022_;
 wire _20023_;
 wire _20024_;
 wire _20025_;
 wire _20026_;
 wire _20027_;
 wire _20028_;
 wire _20029_;
 wire _20030_;
 wire _20031_;
 wire _20032_;
 wire _20033_;
 wire _20034_;
 wire _20035_;
 wire _20036_;
 wire _20037_;
 wire _20038_;
 wire _20039_;
 wire _20040_;
 wire _20041_;
 wire _20042_;
 wire _20043_;
 wire _20044_;
 wire _20045_;
 wire _20046_;
 wire _20047_;
 wire _20048_;
 wire _20049_;
 wire _20050_;
 wire _20051_;
 wire _20052_;
 wire _20053_;
 wire _20054_;
 wire _20055_;
 wire _20056_;
 wire _20057_;
 wire _20058_;
 wire _20059_;
 wire _20060_;
 wire _20061_;
 wire _20062_;
 wire _20063_;
 wire _20064_;
 wire _20065_;
 wire _20066_;
 wire _20067_;
 wire _20068_;
 wire _20069_;
 wire _20070_;
 wire _20071_;
 wire _20072_;
 wire _20073_;
 wire _20074_;
 wire _20075_;
 wire _20076_;
 wire _20077_;
 wire _20078_;
 wire _20079_;
 wire _20080_;
 wire _20081_;
 wire _20082_;
 wire _20083_;
 wire _20084_;
 wire _20085_;
 wire _20086_;
 wire _20087_;
 wire _20088_;
 wire _20089_;
 wire _20090_;
 wire _20091_;
 wire _20092_;
 wire _20093_;
 wire _20094_;
 wire _20095_;
 wire _20096_;
 wire _20097_;
 wire _20098_;
 wire _20099_;
 wire _20100_;
 wire _20101_;
 wire _20102_;
 wire _20103_;
 wire _20104_;
 wire _20105_;
 wire _20106_;
 wire _20107_;
 wire _20108_;
 wire _20109_;
 wire _20110_;
 wire _20111_;
 wire _20112_;
 wire _20113_;
 wire _20114_;
 wire _20115_;
 wire _20116_;
 wire _20117_;
 wire _20118_;
 wire _20119_;
 wire _20120_;
 wire _20121_;
 wire _20122_;
 wire _20123_;
 wire _20124_;
 wire _20125_;
 wire _20126_;
 wire _20127_;
 wire _20128_;
 wire _20129_;
 wire _20130_;
 wire _20131_;
 wire _20132_;
 wire _20133_;
 wire _20134_;
 wire _20135_;
 wire _20136_;
 wire _20137_;
 wire _20138_;
 wire _20139_;
 wire _20140_;
 wire _20141_;
 wire _20142_;
 wire _20143_;
 wire _20144_;
 wire _20145_;
 wire _20146_;
 wire _20147_;
 wire _20148_;
 wire _20149_;
 wire _20150_;
 wire _20151_;
 wire _20152_;
 wire _20153_;
 wire _20154_;
 wire _20155_;
 wire _20156_;
 wire _20157_;
 wire _20158_;
 wire _20159_;
 wire _20160_;
 wire _20161_;
 wire _20162_;
 wire _20163_;
 wire _20164_;
 wire _20165_;
 wire _20166_;
 wire _20167_;
 wire _20168_;
 wire _20169_;
 wire _20170_;
 wire _20171_;
 wire _20172_;
 wire _20173_;
 wire _20174_;
 wire _20175_;
 wire _20176_;
 wire _20177_;
 wire _20178_;
 wire _20179_;
 wire _20180_;
 wire _20181_;
 wire _20182_;
 wire _20183_;
 wire _20184_;
 wire _20185_;
 wire _20186_;
 wire _20187_;
 wire _20188_;
 wire _20189_;
 wire _20190_;
 wire _20191_;
 wire _20192_;
 wire _20193_;
 wire _20194_;
 wire _20195_;
 wire _20196_;
 wire _20197_;
 wire _20198_;
 wire _20199_;
 wire _20200_;
 wire _20201_;
 wire _20202_;
 wire _20203_;
 wire _20204_;
 wire _20205_;
 wire _20206_;
 wire _20207_;
 wire _20208_;
 wire _20209_;
 wire _20210_;
 wire _20211_;
 wire _20212_;
 wire _20213_;
 wire _20214_;
 wire _20215_;
 wire _20216_;
 wire _20217_;
 wire _20218_;
 wire _20219_;
 wire _20220_;
 wire _20221_;
 wire _20222_;
 wire _20223_;
 wire _20224_;
 wire _20225_;
 wire _20226_;
 wire _20227_;
 wire _20228_;
 wire _20229_;
 wire _20230_;
 wire _20231_;
 wire _20232_;
 wire _20233_;
 wire _20234_;
 wire _20235_;
 wire _20236_;
 wire _20237_;
 wire _20238_;
 wire _20239_;
 wire _20240_;
 wire _20241_;
 wire _20242_;
 wire _20243_;
 wire _20244_;
 wire _20245_;
 wire _20246_;
 wire _20247_;
 wire _20248_;
 wire _20249_;
 wire _20250_;
 wire _20251_;
 wire _20252_;
 wire _20253_;
 wire _20254_;
 wire _20255_;
 wire _20256_;
 wire _20257_;
 wire _20258_;
 wire _20259_;
 wire _20260_;
 wire _20261_;
 wire _20262_;
 wire _20263_;
 wire _20264_;
 wire _20265_;
 wire _20266_;
 wire _20267_;
 wire _20268_;
 wire _20269_;
 wire _20270_;
 wire _20271_;
 wire _20272_;
 wire _20273_;
 wire _20274_;
 wire _20275_;
 wire _20276_;
 wire _20277_;
 wire _20278_;
 wire _20279_;
 wire _20280_;
 wire _20281_;
 wire _20282_;
 wire _20283_;
 wire _20284_;
 wire _20285_;
 wire _20286_;
 wire _20287_;
 wire _20288_;
 wire _20289_;
 wire _20290_;
 wire _20291_;
 wire _20292_;
 wire _20293_;
 wire _20294_;
 wire _20295_;
 wire _20296_;
 wire _20297_;
 wire _20298_;
 wire _20299_;
 wire _20300_;
 wire _20301_;
 wire _20302_;
 wire _20303_;
 wire _20304_;
 wire _20305_;
 wire _20306_;
 wire _20307_;
 wire _20308_;
 wire _20309_;
 wire _20310_;
 wire _20311_;
 wire _20312_;
 wire _20313_;
 wire _20314_;
 wire _20315_;
 wire _20316_;
 wire _20317_;
 wire _20318_;
 wire _20319_;
 wire _20320_;
 wire _20321_;
 wire _20322_;
 wire _20323_;
 wire _20324_;
 wire _20325_;
 wire _20326_;
 wire _20327_;
 wire _20328_;
 wire _20329_;
 wire _20330_;
 wire _20331_;
 wire _20332_;
 wire _20333_;
 wire _20334_;
 wire _20335_;
 wire _20336_;
 wire _20337_;
 wire _20338_;
 wire _20339_;
 wire _20340_;
 wire _20341_;
 wire _20342_;
 wire _20343_;
 wire _20344_;
 wire _20345_;
 wire _20346_;
 wire _20347_;
 wire _20348_;
 wire _20349_;
 wire _20350_;
 wire _20351_;
 wire _20352_;
 wire _20353_;
 wire _20354_;
 wire _20355_;
 wire _20356_;
 wire _20357_;
 wire _20358_;
 wire _20359_;
 wire _20360_;
 wire _20361_;
 wire _20362_;
 wire _20363_;
 wire _20364_;
 wire _20365_;
 wire _20366_;
 wire _20367_;
 wire _20368_;
 wire _20369_;
 wire _20370_;
 wire _20371_;
 wire _20372_;
 wire _20373_;
 wire _20374_;
 wire _20375_;
 wire _20376_;
 wire _20377_;
 wire _20378_;
 wire _20379_;
 wire _20380_;
 wire _20381_;
 wire _20382_;
 wire _20383_;
 wire _20384_;
 wire _20385_;
 wire _20386_;
 wire _20387_;
 wire _20388_;
 wire _20389_;
 wire _20390_;
 wire _20391_;
 wire _20392_;
 wire _20393_;
 wire _20394_;
 wire _20395_;
 wire _20396_;
 wire _20397_;
 wire _20398_;
 wire _20399_;
 wire _20400_;
 wire _20401_;
 wire _20402_;
 wire _20403_;
 wire _20404_;
 wire _20405_;
 wire _20406_;
 wire _20407_;
 wire _20408_;
 wire _20409_;
 wire _20410_;
 wire _20411_;
 wire _20412_;
 wire _20413_;
 wire _20414_;
 wire _20415_;
 wire _20416_;
 wire _20417_;
 wire _20418_;
 wire _20419_;
 wire _20420_;
 wire _20421_;
 wire _20422_;
 wire _20423_;
 wire _20424_;
 wire _20425_;
 wire _20426_;
 wire _20427_;
 wire _20428_;
 wire _20429_;
 wire _20430_;
 wire _20431_;
 wire _20432_;
 wire _20433_;
 wire _20434_;
 wire _20435_;
 wire _20436_;
 wire _20437_;
 wire _20438_;
 wire _20439_;
 wire _20440_;
 wire _20441_;
 wire _20442_;
 wire _20443_;
 wire _20444_;
 wire _20445_;
 wire _20446_;
 wire _20447_;
 wire _20448_;
 wire _20449_;
 wire _20450_;
 wire _20451_;
 wire _20452_;
 wire _20453_;
 wire _20454_;
 wire _20455_;
 wire _20456_;
 wire _20457_;
 wire _20458_;
 wire _20459_;
 wire _20460_;
 wire _20461_;
 wire _20462_;
 wire _20463_;
 wire _20464_;
 wire _20465_;
 wire _20466_;
 wire _20467_;
 wire _20468_;
 wire _20469_;
 wire _20470_;
 wire _20471_;
 wire _20472_;
 wire _20473_;
 wire _20474_;
 wire _20475_;
 wire _20476_;
 wire _20477_;
 wire _20478_;
 wire _20479_;
 wire _20480_;
 wire _20481_;
 wire _20482_;
 wire _20483_;
 wire _20484_;
 wire _20485_;
 wire _20486_;
 wire _20487_;
 wire _20488_;
 wire _20489_;
 wire _20490_;
 wire _20491_;
 wire _20492_;
 wire _20493_;
 wire _20494_;
 wire _20495_;
 wire _20496_;
 wire _20497_;
 wire _20498_;
 wire _20499_;
 wire _20500_;
 wire _20501_;
 wire _20502_;
 wire _20503_;
 wire _20504_;
 wire _20505_;
 wire _20506_;
 wire _20507_;
 wire _20508_;
 wire _20509_;
 wire _20510_;
 wire _20511_;
 wire _20512_;
 wire _20513_;
 wire _20514_;
 wire _20515_;
 wire _20516_;
 wire _20517_;
 wire _20518_;
 wire _20519_;
 wire _20520_;
 wire _20521_;
 wire _20522_;
 wire _20523_;
 wire _20524_;
 wire _20525_;
 wire _20526_;
 wire _20527_;
 wire _20528_;
 wire _20529_;
 wire _20530_;
 wire _20531_;
 wire _20532_;
 wire _20533_;
 wire _20534_;
 wire _20535_;
 wire _20536_;
 wire _20537_;
 wire _20538_;
 wire _20539_;
 wire _20540_;
 wire _20541_;
 wire _20542_;
 wire _20543_;
 wire _20544_;
 wire _20545_;
 wire _20546_;
 wire _20547_;
 wire _20548_;
 wire _20549_;
 wire _20550_;
 wire _20551_;
 wire _20552_;
 wire _20553_;
 wire _20554_;
 wire _20555_;
 wire _20556_;
 wire _20557_;
 wire _20558_;
 wire _20559_;
 wire _20560_;
 wire _20561_;
 wire _20562_;
 wire _20563_;
 wire _20564_;
 wire _20565_;
 wire _20566_;
 wire _20567_;
 wire _20568_;
 wire _20569_;
 wire _20570_;
 wire _20571_;
 wire _20572_;
 wire _20573_;
 wire _20574_;
 wire _20575_;
 wire _20576_;
 wire _20577_;
 wire _20578_;
 wire _20579_;
 wire _20580_;
 wire _20581_;
 wire _20582_;
 wire _20583_;
 wire _20584_;
 wire _20585_;
 wire _20586_;
 wire _20587_;
 wire _20588_;
 wire _20589_;
 wire _20590_;
 wire _20591_;
 wire _20592_;
 wire _20593_;
 wire _20594_;
 wire _20595_;
 wire _20596_;
 wire _20597_;
 wire _20598_;
 wire _20599_;
 wire _20600_;
 wire _20601_;
 wire _20602_;
 wire _20603_;
 wire _20604_;
 wire _20605_;
 wire _20606_;
 wire _20607_;
 wire _20608_;
 wire _20609_;
 wire _20610_;
 wire _20611_;
 wire _20612_;
 wire _20613_;
 wire _20614_;
 wire _20615_;
 wire _20616_;
 wire _20617_;
 wire _20618_;
 wire _20619_;
 wire _20620_;
 wire _20621_;
 wire _20622_;
 wire _20623_;
 wire _20624_;
 wire _20625_;
 wire _20626_;
 wire _20627_;
 wire _20628_;
 wire _20629_;
 wire _20630_;
 wire _20631_;
 wire _20632_;
 wire _20633_;
 wire _20634_;
 wire _20635_;
 wire _20636_;
 wire _20637_;
 wire _20638_;
 wire _20639_;
 wire _20640_;
 wire _20641_;
 wire _20642_;
 wire _20643_;
 wire _20644_;
 wire _20645_;
 wire _20646_;
 wire _20647_;
 wire _20648_;
 wire _20649_;
 wire _20650_;
 wire _20651_;
 wire _20652_;
 wire _20653_;
 wire _20654_;
 wire _20655_;
 wire _20656_;
 wire _20657_;
 wire _20658_;
 wire _20659_;
 wire _20660_;
 wire _20661_;
 wire _20662_;
 wire _20663_;
 wire _20664_;
 wire _20665_;
 wire _20666_;
 wire _20667_;
 wire _20668_;
 wire _20669_;
 wire _20670_;
 wire _20671_;
 wire _20672_;
 wire _20673_;
 wire _20674_;
 wire _20675_;
 wire _20676_;
 wire _20677_;
 wire _20678_;
 wire _20679_;
 wire _20680_;
 wire _20681_;
 wire _20682_;
 wire _20683_;
 wire _20684_;
 wire _20685_;
 wire _20686_;
 wire _20687_;
 wire _20688_;
 wire _20689_;
 wire _20690_;
 wire _20691_;
 wire _20692_;
 wire _20693_;
 wire _20694_;
 wire _20695_;
 wire _20696_;
 wire _20697_;
 wire _20698_;
 wire _20699_;
 wire _20700_;
 wire _20701_;
 wire _20702_;
 wire _20703_;
 wire _20704_;
 wire _20705_;
 wire _20706_;
 wire _20707_;
 wire _20708_;
 wire _20709_;
 wire _20710_;
 wire _20711_;
 wire _20712_;
 wire _20713_;
 wire _20714_;
 wire _20715_;
 wire _20716_;
 wire _20717_;
 wire _20718_;
 wire _20719_;
 wire _20720_;
 wire _20721_;
 wire _20722_;
 wire _20723_;
 wire _20724_;
 wire _20725_;
 wire _20726_;
 wire _20727_;
 wire _20728_;
 wire _20729_;
 wire _20730_;
 wire _20731_;
 wire _20732_;
 wire _20733_;
 wire _20734_;
 wire _20735_;
 wire _20736_;
 wire _20737_;
 wire _20738_;
 wire _20739_;
 wire _20740_;
 wire _20741_;
 wire _20742_;
 wire _20743_;
 wire _20744_;
 wire _20745_;
 wire _20746_;
 wire _20747_;
 wire _20748_;
 wire _20749_;
 wire _20750_;
 wire _20751_;
 wire _20752_;
 wire _20753_;
 wire _20754_;
 wire _20755_;
 wire _20756_;
 wire _20757_;
 wire _20758_;
 wire _20759_;
 wire _20760_;
 wire _20761_;
 wire _20762_;
 wire _20763_;
 wire _20764_;
 wire _20765_;
 wire _20766_;
 wire _20767_;
 wire _20768_;
 wire _20769_;
 wire _20770_;
 wire _20771_;
 wire _20772_;
 wire _20773_;
 wire _20774_;
 wire _20775_;
 wire _20776_;
 wire _20777_;
 wire _20778_;
 wire _20779_;
 wire _20780_;
 wire _20781_;
 wire _20782_;
 wire _20783_;
 wire _20784_;
 wire _20785_;
 wire _20786_;
 wire _20787_;
 wire _20788_;
 wire _20789_;
 wire _20790_;
 wire _20791_;
 wire _20792_;
 wire _20793_;
 wire _20794_;
 wire _20795_;
 wire _20796_;
 wire _20797_;
 wire _20798_;
 wire _20799_;
 wire _20800_;
 wire _20801_;
 wire _20802_;
 wire _20803_;
 wire _20804_;
 wire _20805_;
 wire _20806_;
 wire _20807_;
 wire _20808_;
 wire _20809_;
 wire _20810_;
 wire _20811_;
 wire _20812_;
 wire _20813_;
 wire _20814_;
 wire _20815_;
 wire _20816_;
 wire _20817_;
 wire _20818_;
 wire _20819_;
 wire _20820_;
 wire _20821_;
 wire _20822_;
 wire _20823_;
 wire _20824_;
 wire _20825_;
 wire _20826_;
 wire _20827_;
 wire _20828_;
 wire _20829_;
 wire _20830_;
 wire _20831_;
 wire _20832_;
 wire _20833_;
 wire _20834_;
 wire _20835_;
 wire _20836_;
 wire _20837_;
 wire _20838_;
 wire _20839_;
 wire _20840_;
 wire _20841_;
 wire _20842_;
 wire _20843_;
 wire _20844_;
 wire _20845_;
 wire _20846_;
 wire _20847_;
 wire _20848_;
 wire _20849_;
 wire _20850_;
 wire _20851_;
 wire _20852_;
 wire _20853_;
 wire _20854_;
 wire _20855_;
 wire _20856_;
 wire _20857_;
 wire _20858_;
 wire _20859_;
 wire _20860_;
 wire _20861_;
 wire _20862_;
 wire _20863_;
 wire _20864_;
 wire _20865_;
 wire _20866_;
 wire _20867_;
 wire _20868_;
 wire _20869_;
 wire _20870_;
 wire _20871_;
 wire _20872_;
 wire _20873_;
 wire _20874_;
 wire _20875_;
 wire _20876_;
 wire _20877_;
 wire _20878_;
 wire _20879_;
 wire _20880_;
 wire _20881_;
 wire _20882_;
 wire _20883_;
 wire _20884_;
 wire _20885_;
 wire _20886_;
 wire _20887_;
 wire _20888_;
 wire _20889_;
 wire _20890_;
 wire _20891_;
 wire _20892_;
 wire _20893_;
 wire _20894_;
 wire _20895_;
 wire _20896_;
 wire _20897_;
 wire _20898_;
 wire _20899_;
 wire _20900_;
 wire _20901_;
 wire _20902_;
 wire _20903_;
 wire _20904_;
 wire _20905_;
 wire _20906_;
 wire _20907_;
 wire _20908_;
 wire _20909_;
 wire _20910_;
 wire _20911_;
 wire _20912_;
 wire _20913_;
 wire _20914_;
 wire _20915_;
 wire _20916_;
 wire _20917_;
 wire _20918_;
 wire _20919_;
 wire _20920_;
 wire _20921_;
 wire _20922_;
 wire _20923_;
 wire _20924_;
 wire _20925_;
 wire _20926_;
 wire _20927_;
 wire _20928_;
 wire _20929_;
 wire _20930_;
 wire _20931_;
 wire _20932_;
 wire _20933_;
 wire _20934_;
 wire _20935_;
 wire _20936_;
 wire _20937_;
 wire _20938_;
 wire _20939_;
 wire _20940_;
 wire _20941_;
 wire _20942_;
 wire _20943_;
 wire _20944_;
 wire _20945_;
 wire _20946_;
 wire _20947_;
 wire _20948_;
 wire _20949_;
 wire _20950_;
 wire _20951_;
 wire _20952_;
 wire _20953_;
 wire _20954_;
 wire _20955_;
 wire _20956_;
 wire _20957_;
 wire _20958_;
 wire _20959_;
 wire _20960_;
 wire _20961_;
 wire _20962_;
 wire _20963_;
 wire _20964_;
 wire _20965_;
 wire _20966_;
 wire _20967_;
 wire _20968_;
 wire _20969_;
 wire _20970_;
 wire _20971_;
 wire _20972_;
 wire _20973_;
 wire _20974_;
 wire _20975_;
 wire _20976_;
 wire _20977_;
 wire _20978_;
 wire _20979_;
 wire _20980_;
 wire _20981_;
 wire _20982_;
 wire _20983_;
 wire _20984_;
 wire _20985_;
 wire _20986_;
 wire _20987_;
 wire _20988_;
 wire _20989_;
 wire _20990_;
 wire _20991_;
 wire _20992_;
 wire _20993_;
 wire _20994_;
 wire _20995_;
 wire _20996_;
 wire _20997_;
 wire _20998_;
 wire _20999_;
 wire _21000_;
 wire _21001_;
 wire _21002_;
 wire _21003_;
 wire _21004_;
 wire _21005_;
 wire _21006_;
 wire _21007_;
 wire _21008_;
 wire _21009_;
 wire _21010_;
 wire _21011_;
 wire _21012_;
 wire _21013_;
 wire _21014_;
 wire _21015_;
 wire _21016_;
 wire _21017_;
 wire _21018_;
 wire _21019_;
 wire _21020_;
 wire _21021_;
 wire _21022_;
 wire _21023_;
 wire _21024_;
 wire _21025_;
 wire _21026_;
 wire _21027_;
 wire _21028_;
 wire _21029_;
 wire _21030_;
 wire _21031_;
 wire _21032_;
 wire _21033_;
 wire _21034_;
 wire _21035_;
 wire _21036_;
 wire _21037_;
 wire _21038_;
 wire _21039_;
 wire _21040_;
 wire _21041_;
 wire _21042_;
 wire _21043_;
 wire _21044_;
 wire _21045_;
 wire _21046_;
 wire _21047_;
 wire _21048_;
 wire _21049_;
 wire _21050_;
 wire _21051_;
 wire _21052_;
 wire _21053_;
 wire _21054_;
 wire _21055_;
 wire _21056_;
 wire _21057_;
 wire _21058_;
 wire _21059_;
 wire _21060_;
 wire _21061_;
 wire _21062_;
 wire _21063_;
 wire _21064_;
 wire _21065_;
 wire _21066_;
 wire _21067_;
 wire _21068_;
 wire _21069_;
 wire _21070_;
 wire _21071_;
 wire _21072_;
 wire _21073_;
 wire _21074_;
 wire _21075_;
 wire _21076_;
 wire _21077_;
 wire _21078_;
 wire _21079_;
 wire _21080_;
 wire _21081_;
 wire _21082_;
 wire _21083_;
 wire _21084_;
 wire _21085_;
 wire _21086_;
 wire _21087_;
 wire _21088_;
 wire _21089_;
 wire _21090_;
 wire _21091_;
 wire _21092_;
 wire _21093_;
 wire _21094_;
 wire _21095_;
 wire _21096_;
 wire _21097_;
 wire _21098_;
 wire _21099_;
 wire _21100_;
 wire _21101_;
 wire _21102_;
 wire _21103_;
 wire _21104_;
 wire _21105_;
 wire _21106_;
 wire _21107_;
 wire _21108_;
 wire _21109_;
 wire _21110_;
 wire _21111_;
 wire _21112_;
 wire _21113_;
 wire _21114_;
 wire _21115_;
 wire _21116_;
 wire _21117_;
 wire _21118_;
 wire _21119_;
 wire _21120_;
 wire _21121_;
 wire _21122_;
 wire _21123_;
 wire _21124_;
 wire _21125_;
 wire _21126_;
 wire _21127_;
 wire _21128_;
 wire _21129_;
 wire _21130_;
 wire _21131_;
 wire _21132_;
 wire _21133_;
 wire _21134_;
 wire _21135_;
 wire _21136_;
 wire _21137_;
 wire _21138_;
 wire _21139_;
 wire _21140_;
 wire _21141_;
 wire _21142_;
 wire _21143_;
 wire _21144_;
 wire _21145_;
 wire _21146_;
 wire _21147_;
 wire _21148_;
 wire _21149_;
 wire _21150_;
 wire _21151_;
 wire _21152_;
 wire _21153_;
 wire _21154_;
 wire _21155_;
 wire _21156_;
 wire _21157_;
 wire _21158_;
 wire _21159_;
 wire _21160_;
 wire _21161_;
 wire _21162_;
 wire _21163_;
 wire _21164_;
 wire _21165_;
 wire _21166_;
 wire _21167_;
 wire _21168_;
 wire _21169_;
 wire _21170_;
 wire _21171_;
 wire _21172_;
 wire _21173_;
 wire _21174_;
 wire _21175_;
 wire _21176_;
 wire _21177_;
 wire _21178_;
 wire _21179_;
 wire _21180_;
 wire _21181_;
 wire _21182_;
 wire _21183_;
 wire _21184_;
 wire _21185_;
 wire _21186_;
 wire _21187_;
 wire _21188_;
 wire _21189_;
 wire _21190_;
 wire _21191_;
 wire _21192_;
 wire _21193_;
 wire _21194_;
 wire _21195_;
 wire _21196_;
 wire _21197_;
 wire _21198_;
 wire _21199_;
 wire _21200_;
 wire _21201_;
 wire _21202_;
 wire _21203_;
 wire _21204_;
 wire _21205_;
 wire _21206_;
 wire _21207_;
 wire _21208_;
 wire _21209_;
 wire _21210_;
 wire _21211_;
 wire _21212_;
 wire _21213_;
 wire _21214_;
 wire _21215_;
 wire _21216_;
 wire _21217_;
 wire _21218_;
 wire _21219_;
 wire _21220_;
 wire _21221_;
 wire _21222_;
 wire _21223_;
 wire _21224_;
 wire _21225_;
 wire _21226_;
 wire _21227_;
 wire _21228_;
 wire _21229_;
 wire _21230_;
 wire _21231_;
 wire _21232_;
 wire _21233_;
 wire _21234_;
 wire _21235_;
 wire _21236_;
 wire _21237_;
 wire _21238_;
 wire _21239_;
 wire _21240_;
 wire _21241_;
 wire _21242_;
 wire _21243_;
 wire _21244_;
 wire _21245_;
 wire _21246_;
 wire _21247_;
 wire _21248_;
 wire _21249_;
 wire _21250_;
 wire _21251_;
 wire _21252_;
 wire _21253_;
 wire _21254_;
 wire _21255_;
 wire _21256_;
 wire _21257_;
 wire _21258_;
 wire _21259_;
 wire _21260_;
 wire _21261_;
 wire _21262_;
 wire _21263_;
 wire _21264_;
 wire _21265_;
 wire _21266_;
 wire _21267_;
 wire _21268_;
 wire _21269_;
 wire _21270_;
 wire _21271_;
 wire _21272_;
 wire _21273_;
 wire _21274_;
 wire _21275_;
 wire _21276_;
 wire _21277_;
 wire _21278_;
 wire _21279_;
 wire _21280_;
 wire _21281_;
 wire _21282_;
 wire _21283_;
 wire _21284_;
 wire _21285_;
 wire _21286_;
 wire _21287_;
 wire _21288_;
 wire _21289_;
 wire _21290_;
 wire _21291_;
 wire _21292_;
 wire _21293_;
 wire _21294_;
 wire _21295_;
 wire _21296_;
 wire _21297_;
 wire _21298_;
 wire _21299_;
 wire _21300_;
 wire _21301_;
 wire _21302_;
 wire _21303_;
 wire _21304_;
 wire _21305_;
 wire _21306_;
 wire _21307_;
 wire _21308_;
 wire _21309_;
 wire _21310_;
 wire _21311_;
 wire _21312_;
 wire _21313_;
 wire _21314_;
 wire _21315_;
 wire _21316_;
 wire _21317_;
 wire _21318_;
 wire _21319_;
 wire _21320_;
 wire _21321_;
 wire _21322_;
 wire _21323_;
 wire _21324_;
 wire _21325_;
 wire _21326_;
 wire _21327_;
 wire _21328_;
 wire _21329_;
 wire _21330_;
 wire _21331_;
 wire _21332_;
 wire _21333_;
 wire _21334_;
 wire _21335_;
 wire _21336_;
 wire _21337_;
 wire _21338_;
 wire _21339_;
 wire _21340_;
 wire _21341_;
 wire _21342_;
 wire _21343_;
 wire _21344_;
 wire _21345_;
 wire _21346_;
 wire _21347_;
 wire _21348_;
 wire _21349_;
 wire _21350_;
 wire _21351_;
 wire _21352_;
 wire _21353_;
 wire _21354_;
 wire _21355_;
 wire _21356_;
 wire _21357_;
 wire _21358_;
 wire _21359_;
 wire _21360_;
 wire _21361_;
 wire _21362_;
 wire _21363_;
 wire _21364_;
 wire _21365_;
 wire _21366_;
 wire _21367_;
 wire _21368_;
 wire _21369_;
 wire _21370_;
 wire _21371_;
 wire _21372_;
 wire _21373_;
 wire _21374_;
 wire _21375_;
 wire _21376_;
 wire _21377_;
 wire _21378_;
 wire _21379_;
 wire _21380_;
 wire _21381_;
 wire _21382_;
 wire _21383_;
 wire _21384_;
 wire _21385_;
 wire _21386_;
 wire _21387_;
 wire _21388_;
 wire _21389_;
 wire _21390_;
 wire _21391_;
 wire _21392_;
 wire _21393_;
 wire _21394_;
 wire _21395_;
 wire _21396_;
 wire _21397_;
 wire _21398_;
 wire _21399_;
 wire _21400_;
 wire _21401_;
 wire _21402_;
 wire _21403_;
 wire _21404_;
 wire _21405_;
 wire _21406_;
 wire _21407_;
 wire _21408_;
 wire _21409_;
 wire _21410_;
 wire _21411_;
 wire _21412_;
 wire _21413_;
 wire _21414_;
 wire _21415_;
 wire _21416_;
 wire _21417_;
 wire _21418_;
 wire _21419_;
 wire _21420_;
 wire _21421_;
 wire _21422_;
 wire _21423_;
 wire _21424_;
 wire _21425_;
 wire _21426_;
 wire _21427_;
 wire _21428_;
 wire _21429_;
 wire _21430_;
 wire _21431_;
 wire _21432_;
 wire _21433_;
 wire _21434_;
 wire _21435_;
 wire _21436_;
 wire _21437_;
 wire _21438_;
 wire _21439_;
 wire _21440_;
 wire _21441_;
 wire _21442_;
 wire _21443_;
 wire _21444_;
 wire _21445_;
 wire _21446_;
 wire _21447_;
 wire _21448_;
 wire _21449_;
 wire _21450_;
 wire _21451_;
 wire _21452_;
 wire _21453_;
 wire _21454_;
 wire _21455_;
 wire _21456_;
 wire _21457_;
 wire _21458_;
 wire _21459_;
 wire _21460_;
 wire _21461_;
 wire _21462_;
 wire _21463_;
 wire _21464_;
 wire _21465_;
 wire _21466_;
 wire _21467_;
 wire _21468_;
 wire _21469_;
 wire _21470_;
 wire _21471_;
 wire _21472_;
 wire _21473_;
 wire _21474_;
 wire _21475_;
 wire _21476_;
 wire _21477_;
 wire _21478_;
 wire _21479_;
 wire _21480_;
 wire _21481_;
 wire _21482_;
 wire _21483_;
 wire _21484_;
 wire _21485_;
 wire _21486_;
 wire _21487_;
 wire _21488_;
 wire _21489_;
 wire _21490_;
 wire _21491_;
 wire _21492_;
 wire _21493_;
 wire _21494_;
 wire _21495_;
 wire _21496_;
 wire _21497_;
 wire _21498_;
 wire _21499_;
 wire _21500_;
 wire _21501_;
 wire _21502_;
 wire _21503_;
 wire _21504_;
 wire _21505_;
 wire _21506_;
 wire _21507_;
 wire _21508_;
 wire _21509_;
 wire _21510_;
 wire _21511_;
 wire _21512_;
 wire _21513_;
 wire _21514_;
 wire _21515_;
 wire _21516_;
 wire _21517_;
 wire _21518_;
 wire _21519_;
 wire _21520_;
 wire _21521_;
 wire _21522_;
 wire _21523_;
 wire _21524_;
 wire _21525_;
 wire _21526_;
 wire _21527_;
 wire _21528_;
 wire _21529_;
 wire _21530_;
 wire _21531_;
 wire _21532_;
 wire _21533_;
 wire _21534_;
 wire _21535_;
 wire _21536_;
 wire _21537_;
 wire _21538_;
 wire _21539_;
 wire _21540_;
 wire _21541_;
 wire _21542_;
 wire _21543_;
 wire _21544_;
 wire _21545_;
 wire _21546_;
 wire _21547_;
 wire _21548_;
 wire _21549_;
 wire _21550_;
 wire _21551_;
 wire _21552_;
 wire _21553_;
 wire _21554_;
 wire _21555_;
 wire _21556_;
 wire _21557_;
 wire _21558_;
 wire _21559_;
 wire _21560_;
 wire _21561_;
 wire _21562_;
 wire _21563_;
 wire _21564_;
 wire _21565_;
 wire _21566_;
 wire _21567_;
 wire _21568_;
 wire _21569_;
 wire _21570_;
 wire _21571_;
 wire _21572_;
 wire _21573_;
 wire _21574_;
 wire _21575_;
 wire _21576_;
 wire _21577_;
 wire _21578_;
 wire _21579_;
 wire _21580_;
 wire _21581_;
 wire _21582_;
 wire _21583_;
 wire _21584_;
 wire _21585_;
 wire _21586_;
 wire _21587_;
 wire _21588_;
 wire _21589_;
 wire _21590_;
 wire _21591_;
 wire _21592_;
 wire _21593_;
 wire _21594_;
 wire _21595_;
 wire _21596_;
 wire _21597_;
 wire _21598_;
 wire _21599_;
 wire _21600_;
 wire _21601_;
 wire _21602_;
 wire _21603_;
 wire _21604_;
 wire _21605_;
 wire _21606_;
 wire _21607_;
 wire _21608_;
 wire _21609_;
 wire _21610_;
 wire _21611_;
 wire _21612_;
 wire _21613_;
 wire _21614_;
 wire _21615_;
 wire _21616_;
 wire _21617_;
 wire _21618_;
 wire _21619_;
 wire _21620_;
 wire _21621_;
 wire _21622_;
 wire _21623_;
 wire _21624_;
 wire _21625_;
 wire _21626_;
 wire _21627_;
 wire _21628_;
 wire _21629_;
 wire _21630_;
 wire _21631_;
 wire _21632_;
 wire _21633_;
 wire _21634_;
 wire _21635_;
 wire _21636_;
 wire _21637_;
 wire _21638_;
 wire _21639_;
 wire _21640_;
 wire _21641_;
 wire _21642_;
 wire _21643_;
 wire _21644_;
 wire _21645_;
 wire _21646_;
 wire _21647_;
 wire _21648_;
 wire _21649_;
 wire _21650_;
 wire _21651_;
 wire _21652_;
 wire _21653_;
 wire _21654_;
 wire _21655_;
 wire _21656_;
 wire _21657_;
 wire _21658_;
 wire _21659_;
 wire _21660_;
 wire _21661_;
 wire _21662_;
 wire _21663_;
 wire _21664_;
 wire _21665_;
 wire _21666_;
 wire _21667_;
 wire _21668_;
 wire _21669_;
 wire _21670_;
 wire _21671_;
 wire _21672_;
 wire _21673_;
 wire _21674_;
 wire _21675_;
 wire _21676_;
 wire _21677_;
 wire _21678_;
 wire _21679_;
 wire _21680_;
 wire _21681_;
 wire _21682_;
 wire _21683_;
 wire _21684_;
 wire _21685_;
 wire _21686_;
 wire _21687_;
 wire _21688_;
 wire _21689_;
 wire _21690_;
 wire _21691_;
 wire _21692_;
 wire _21693_;
 wire _21694_;
 wire _21695_;
 wire _21696_;
 wire _21697_;
 wire _21698_;
 wire _21699_;
 wire _21700_;
 wire _21701_;
 wire _21702_;
 wire _21703_;
 wire _21704_;
 wire _21705_;
 wire _21706_;
 wire _21707_;
 wire _21708_;
 wire _21709_;
 wire _21710_;
 wire _21711_;
 wire _21712_;
 wire _21713_;
 wire _21714_;
 wire _21715_;
 wire _21716_;
 wire _21717_;
 wire _21718_;
 wire _21719_;
 wire _21720_;
 wire _21721_;
 wire _21722_;
 wire _21723_;
 wire _21724_;
 wire _21725_;
 wire _21726_;
 wire _21727_;
 wire _21728_;
 wire _21729_;
 wire _21730_;
 wire _21731_;
 wire _21732_;
 wire _21733_;
 wire _21734_;
 wire _21735_;
 wire _21736_;
 wire _21737_;
 wire _21738_;
 wire _21739_;
 wire _21740_;
 wire _21741_;
 wire _21742_;
 wire _21743_;
 wire _21744_;
 wire _21745_;
 wire _21746_;
 wire _21747_;
 wire _21748_;
 wire _21749_;
 wire _21750_;
 wire _21751_;
 wire _21752_;
 wire _21753_;
 wire _21754_;
 wire _21755_;
 wire _21756_;
 wire _21757_;
 wire _21758_;
 wire _21759_;
 wire _21760_;
 wire _21761_;
 wire _21762_;
 wire _21763_;
 wire _21764_;
 wire _21765_;
 wire _21766_;
 wire _21767_;
 wire _21768_;
 wire _21769_;
 wire _21770_;
 wire _21771_;
 wire _21772_;
 wire _21773_;
 wire _21774_;
 wire _21775_;
 wire _21776_;
 wire _21777_;
 wire _21778_;
 wire _21779_;
 wire _21780_;
 wire _21781_;
 wire _21782_;
 wire _21783_;
 wire _21784_;
 wire _21785_;
 wire _21786_;
 wire _21787_;
 wire _21788_;
 wire _21789_;
 wire _21790_;
 wire _21791_;
 wire _21792_;
 wire _21793_;
 wire _21794_;
 wire _21795_;
 wire _21796_;
 wire _21797_;
 wire _21798_;
 wire _21799_;
 wire _21800_;
 wire _21801_;
 wire _21802_;
 wire _21803_;
 wire _21804_;
 wire _21805_;
 wire _21806_;
 wire _21807_;
 wire _21808_;
 wire _21809_;
 wire _21810_;
 wire _21811_;
 wire _21812_;
 wire _21813_;
 wire _21814_;
 wire _21815_;
 wire _21816_;
 wire _21817_;
 wire _21818_;
 wire _21819_;
 wire _21820_;
 wire _21821_;
 wire _21822_;
 wire _21823_;
 wire _21824_;
 wire _21825_;
 wire _21826_;
 wire _21827_;
 wire _21828_;
 wire _21829_;
 wire _21830_;
 wire _21831_;
 wire _21832_;
 wire _21833_;
 wire _21834_;
 wire _21835_;
 wire _21836_;
 wire _21837_;
 wire _21838_;
 wire _21839_;
 wire _21840_;
 wire _21841_;
 wire _21842_;
 wire _21843_;
 wire _21844_;
 wire _21845_;
 wire _21846_;
 wire _21847_;
 wire _21848_;
 wire _21849_;
 wire _21850_;
 wire _21851_;
 wire _21852_;
 wire _21853_;
 wire _21854_;
 wire _21855_;
 wire _21856_;
 wire _21857_;
 wire _21858_;
 wire _21859_;
 wire _21860_;
 wire _21861_;
 wire _21862_;
 wire _21863_;
 wire _21864_;
 wire _21865_;
 wire _21866_;
 wire _21867_;
 wire _21868_;
 wire _21869_;
 wire _21870_;
 wire _21871_;
 wire _21872_;
 wire _21873_;
 wire _21874_;
 wire _21875_;
 wire _21876_;
 wire _21877_;
 wire _21878_;
 wire _21879_;
 wire _21880_;
 wire _21881_;
 wire _21882_;
 wire _21883_;
 wire _21884_;
 wire _21885_;
 wire _21886_;
 wire _21887_;
 wire _21888_;
 wire _21889_;
 wire _21890_;
 wire _21891_;
 wire _21892_;
 wire _21893_;
 wire _21894_;
 wire _21895_;
 wire _21896_;
 wire _21897_;
 wire _21898_;
 wire _21899_;
 wire _21900_;
 wire _21901_;
 wire _21902_;
 wire _21903_;
 wire _21904_;
 wire _21905_;
 wire _21906_;
 wire _21907_;
 wire _21908_;
 wire _21909_;
 wire _21910_;
 wire _21911_;
 wire _21912_;
 wire _21913_;
 wire _21914_;
 wire _21915_;
 wire _21916_;
 wire _21917_;
 wire _21918_;
 wire _21919_;
 wire _21920_;
 wire _21921_;
 wire _21922_;
 wire _21923_;
 wire _21924_;
 wire _21925_;
 wire _21926_;
 wire _21927_;
 wire _21928_;
 wire _21929_;
 wire _21930_;
 wire _21931_;
 wire _21932_;
 wire _21933_;
 wire _21934_;
 wire _21935_;
 wire _21936_;
 wire _21937_;
 wire _21938_;
 wire _21939_;
 wire _21940_;
 wire _21941_;
 wire _21942_;
 wire _21943_;
 wire _21944_;
 wire _21945_;
 wire _21946_;
 wire _21947_;
 wire _21948_;
 wire _21949_;
 wire _21950_;
 wire _21951_;
 wire _21952_;
 wire _21953_;
 wire _21954_;
 wire _21955_;
 wire _21956_;
 wire _21957_;
 wire _21958_;
 wire _21959_;
 wire _21960_;
 wire _21961_;
 wire _21962_;
 wire _21963_;
 wire _21964_;
 wire _21965_;
 wire _21966_;
 wire _21967_;
 wire _21968_;
 wire _21969_;
 wire _21970_;
 wire _21971_;
 wire _21972_;
 wire _21973_;
 wire _21974_;
 wire _21975_;
 wire _21976_;
 wire _21977_;
 wire _21978_;
 wire _21979_;
 wire _21980_;
 wire _21981_;
 wire _21982_;
 wire _21983_;
 wire _21984_;
 wire _21985_;
 wire _21986_;
 wire _21987_;
 wire _21988_;
 wire _21989_;
 wire _21990_;
 wire _21991_;
 wire _21992_;
 wire _21993_;
 wire _21994_;
 wire _21995_;
 wire _21996_;
 wire _21997_;
 wire _21998_;
 wire _21999_;
 wire _22000_;
 wire _22001_;
 wire _22002_;
 wire _22003_;
 wire _22004_;
 wire _22005_;
 wire _22006_;
 wire _22007_;
 wire _22008_;
 wire _22009_;
 wire _22010_;
 wire _22011_;
 wire _22012_;
 wire _22013_;
 wire _22014_;
 wire _22015_;
 wire _22016_;
 wire _22017_;
 wire _22018_;
 wire _22019_;
 wire _22020_;
 wire _22021_;
 wire _22022_;
 wire _22023_;
 wire _22024_;
 wire _22025_;
 wire _22026_;
 wire _22027_;
 wire _22028_;
 wire _22029_;
 wire _22030_;
 wire _22031_;
 wire _22032_;
 wire _22033_;
 wire _22034_;
 wire _22035_;
 wire _22036_;
 wire _22037_;
 wire _22038_;
 wire _22039_;
 wire _22040_;
 wire _22041_;
 wire _22042_;
 wire _22043_;
 wire _22044_;
 wire _22045_;
 wire _22046_;
 wire _22047_;
 wire _22048_;
 wire _22049_;
 wire _22050_;
 wire _22051_;
 wire _22052_;
 wire _22053_;
 wire _22054_;
 wire _22055_;
 wire _22056_;
 wire _22057_;
 wire _22058_;
 wire _22059_;
 wire _22060_;
 wire _22061_;
 wire _22062_;
 wire _22063_;
 wire _22064_;
 wire _22065_;
 wire _22066_;
 wire _22067_;
 wire _22068_;
 wire _22069_;
 wire _22070_;
 wire _22071_;
 wire _22072_;
 wire _22073_;
 wire _22074_;
 wire _22075_;
 wire _22076_;
 wire _22077_;
 wire _22078_;
 wire _22079_;
 wire _22080_;
 wire _22081_;
 wire _22082_;
 wire _22083_;
 wire _22084_;
 wire _22085_;
 wire _22086_;
 wire _22087_;
 wire _22088_;
 wire _22089_;
 wire _22090_;
 wire _22091_;
 wire _22092_;
 wire _22093_;
 wire _22094_;
 wire _22095_;
 wire _22096_;
 wire _22097_;
 wire _22098_;
 wire _22099_;
 wire _22100_;
 wire _22101_;
 wire _22102_;
 wire _22103_;
 wire _22104_;
 wire _22105_;
 wire _22106_;
 wire _22107_;
 wire _22108_;
 wire _22109_;
 wire _22110_;
 wire _22111_;
 wire _22112_;
 wire _22113_;
 wire _22114_;
 wire _22115_;
 wire _22116_;
 wire _22117_;
 wire _22118_;
 wire _22119_;
 wire _22120_;
 wire _22121_;
 wire _22122_;
 wire _22123_;
 wire _22124_;
 wire _22125_;
 wire _22126_;
 wire _22127_;
 wire _22128_;
 wire _22129_;
 wire _22130_;
 wire _22131_;
 wire _22132_;
 wire _22133_;
 wire _22134_;
 wire _22135_;
 wire _22136_;
 wire _22137_;
 wire _22138_;
 wire _22139_;
 wire _22140_;
 wire _22141_;
 wire _22142_;
 wire _22143_;
 wire _22144_;
 wire _22145_;
 wire _22146_;
 wire _22147_;
 wire _22148_;
 wire _22149_;
 wire _22150_;
 wire _22151_;
 wire _22152_;
 wire _22153_;
 wire _22154_;
 wire _22155_;
 wire _22156_;
 wire _22157_;
 wire _22158_;
 wire _22159_;
 wire _22160_;
 wire _22161_;
 wire _22162_;
 wire _22163_;
 wire _22164_;
 wire _22165_;
 wire _22166_;
 wire _22167_;
 wire _22168_;
 wire _22169_;
 wire _22170_;
 wire _22171_;
 wire _22172_;
 wire _22173_;
 wire _22174_;
 wire _22175_;
 wire _22176_;
 wire _22177_;
 wire _22178_;
 wire _22179_;
 wire _22180_;
 wire _22181_;
 wire _22182_;
 wire _22183_;
 wire _22184_;
 wire _22185_;
 wire _22186_;
 wire _22187_;
 wire _22188_;
 wire _22189_;
 wire _22190_;
 wire _22191_;
 wire _22192_;
 wire _22193_;
 wire _22194_;
 wire _22195_;
 wire _22196_;
 wire _22197_;
 wire _22198_;
 wire _22199_;
 wire _22200_;
 wire _22201_;
 wire _22202_;
 wire _22203_;
 wire _22204_;
 wire _22205_;
 wire _22206_;
 wire _22207_;
 wire _22208_;
 wire _22209_;
 wire _22210_;
 wire _22211_;
 wire _22212_;
 wire _22213_;
 wire _22214_;
 wire _22215_;
 wire _22216_;
 wire _22217_;
 wire _22218_;
 wire _22219_;
 wire _22220_;
 wire _22221_;
 wire _22222_;
 wire _22223_;
 wire _22224_;
 wire _22225_;
 wire _22226_;
 wire _22227_;
 wire _22228_;
 wire _22229_;
 wire _22230_;
 wire _22231_;
 wire _22232_;
 wire _22233_;
 wire _22234_;
 wire _22235_;
 wire _22236_;
 wire _22237_;
 wire _22238_;
 wire _22239_;
 wire _22240_;
 wire _22241_;
 wire _22242_;
 wire _22243_;
 wire _22244_;
 wire _22245_;
 wire _22246_;
 wire _22247_;
 wire _22248_;
 wire _22249_;
 wire _22250_;
 wire _22251_;
 wire _22252_;
 wire _22253_;
 wire _22254_;
 wire _22255_;
 wire _22256_;
 wire _22257_;
 wire _22258_;
 wire _22259_;
 wire _22260_;
 wire _22261_;
 wire _22262_;
 wire _22263_;
 wire _22264_;
 wire _22265_;
 wire _22266_;
 wire _22267_;
 wire _22268_;
 wire _22269_;
 wire _22270_;
 wire _22271_;
 wire _22272_;
 wire _22273_;
 wire _22274_;
 wire _22275_;
 wire _22276_;
 wire _22277_;
 wire _22278_;
 wire _22279_;
 wire _22280_;
 wire _22281_;
 wire _22282_;
 wire _22283_;
 wire _22284_;
 wire _22285_;
 wire _22286_;
 wire _22287_;
 wire _22288_;
 wire _22289_;
 wire _22290_;
 wire _22291_;
 wire _22292_;
 wire _22293_;
 wire _22294_;
 wire _22295_;
 wire _22296_;
 wire _22297_;
 wire _22298_;
 wire _22299_;
 wire _22300_;
 wire _22301_;
 wire _22302_;
 wire _22303_;
 wire _22304_;
 wire _22305_;
 wire _22306_;
 wire _22307_;
 wire _22308_;
 wire _22309_;
 wire _22310_;
 wire _22311_;
 wire _22312_;
 wire _22313_;
 wire _22314_;
 wire _22315_;
 wire _22316_;
 wire _22317_;
 wire _22318_;
 wire _22319_;
 wire _22320_;
 wire _22321_;
 wire _22322_;
 wire _22323_;
 wire _22324_;
 wire _22325_;
 wire _22326_;
 wire _22327_;
 wire _22328_;
 wire _22329_;
 wire _22330_;
 wire _22331_;
 wire _22332_;
 wire _22333_;
 wire _22334_;
 wire _22335_;
 wire _22336_;
 wire _22337_;
 wire _22338_;
 wire _22339_;
 wire _22340_;
 wire _22341_;
 wire _22342_;
 wire _22343_;
 wire _22344_;
 wire _22345_;
 wire _22346_;
 wire _22347_;
 wire _22348_;
 wire _22349_;
 wire _22350_;
 wire _22351_;
 wire _22352_;
 wire _22353_;
 wire _22354_;
 wire _22355_;
 wire _22356_;
 wire _22357_;
 wire _22358_;
 wire _22359_;
 wire _22360_;
 wire _22361_;
 wire _22362_;
 wire _22363_;
 wire _22364_;
 wire _22365_;
 wire _22366_;
 wire _22367_;
 wire _22368_;
 wire _22369_;
 wire _22370_;
 wire _22371_;
 wire _22372_;
 wire _22373_;
 wire _22374_;
 wire _22375_;
 wire _22376_;
 wire _22377_;
 wire _22378_;
 wire _22379_;
 wire _22380_;
 wire _22381_;
 wire _22382_;
 wire _22383_;
 wire _22384_;
 wire _22385_;
 wire _22386_;
 wire _22387_;
 wire _22388_;
 wire _22389_;
 wire _22390_;
 wire _22391_;
 wire _22392_;
 wire _22393_;
 wire _22394_;
 wire _22395_;
 wire _22396_;
 wire _22397_;
 wire _22398_;
 wire _22399_;
 wire _22400_;
 wire _22401_;
 wire _22402_;
 wire _22403_;
 wire _22404_;
 wire _22405_;
 wire _22406_;
 wire _22407_;
 wire _22408_;
 wire _22409_;
 wire _22410_;
 wire _22411_;
 wire _22412_;
 wire _22413_;
 wire _22414_;
 wire _22415_;
 wire _22416_;
 wire _22417_;
 wire _22418_;
 wire _22419_;
 wire _22420_;
 wire _22421_;
 wire _22422_;
 wire _22423_;
 wire _22424_;
 wire _22425_;
 wire _22426_;
 wire _22427_;
 wire _22428_;
 wire _22429_;
 wire _22430_;
 wire _22431_;
 wire _22432_;
 wire _22433_;
 wire _22434_;
 wire _22435_;
 wire _22436_;
 wire _22437_;
 wire _22438_;
 wire _22439_;
 wire _22440_;
 wire _22441_;
 wire _22442_;
 wire _22443_;
 wire _22444_;
 wire _22445_;
 wire _22446_;
 wire _22447_;
 wire _22448_;
 wire _22449_;
 wire _22450_;
 wire _22451_;
 wire _22452_;
 wire _22453_;
 wire _22454_;
 wire _22455_;
 wire _22456_;
 wire _22457_;
 wire _22458_;
 wire _22459_;
 wire _22460_;
 wire _22461_;
 wire _22462_;
 wire _22463_;
 wire _22464_;
 wire _22465_;
 wire _22466_;
 wire _22467_;
 wire _22468_;
 wire _22469_;
 wire _22470_;
 wire _22471_;
 wire _22472_;
 wire _22473_;
 wire _22474_;
 wire _22475_;
 wire _22476_;
 wire _22477_;
 wire _22478_;
 wire _22479_;
 wire _22480_;
 wire _22481_;
 wire _22482_;
 wire _22483_;
 wire _22484_;
 wire _22485_;
 wire _22486_;
 wire _22487_;
 wire _22488_;
 wire _22489_;
 wire _22490_;
 wire _22491_;
 wire _22492_;
 wire _22493_;
 wire _22494_;
 wire _22495_;
 wire _22496_;
 wire _22497_;
 wire _22498_;
 wire _22499_;
 wire _22500_;
 wire _22501_;
 wire _22502_;
 wire _22503_;
 wire _22504_;
 wire _22505_;
 wire _22506_;
 wire _22507_;
 wire _22508_;
 wire _22509_;
 wire _22510_;
 wire _22511_;
 wire _22512_;
 wire _22513_;
 wire _22514_;
 wire _22515_;
 wire _22516_;
 wire _22517_;
 wire _22518_;
 wire _22519_;
 wire _22520_;
 wire _22521_;
 wire _22522_;
 wire _22523_;
 wire _22524_;
 wire _22525_;
 wire _22526_;
 wire _22527_;
 wire _22528_;
 wire _22529_;
 wire _22530_;
 wire _22531_;
 wire _22532_;
 wire _22533_;
 wire _22534_;
 wire _22535_;
 wire _22536_;
 wire _22537_;
 wire _22538_;
 wire _22539_;
 wire _22540_;
 wire _22541_;
 wire _22542_;
 wire _22543_;
 wire _22544_;
 wire _22545_;
 wire _22546_;
 wire _22547_;
 wire _22548_;
 wire _22549_;
 wire _22550_;
 wire _22551_;
 wire _22552_;
 wire _22553_;
 wire _22554_;
 wire _22555_;
 wire _22556_;
 wire _22557_;
 wire _22558_;
 wire _22559_;
 wire _22560_;
 wire _22561_;
 wire _22562_;
 wire _22563_;
 wire _22564_;
 wire _22565_;
 wire _22566_;
 wire _22567_;
 wire _22568_;
 wire _22569_;
 wire _22570_;
 wire _22571_;
 wire _22572_;
 wire _22573_;
 wire _22574_;
 wire _22575_;
 wire _22576_;
 wire _22577_;
 wire _22578_;
 wire _22579_;
 wire _22580_;
 wire _22581_;
 wire _22582_;
 wire _22583_;
 wire _22584_;
 wire _22585_;
 wire _22586_;
 wire _22587_;
 wire _22588_;
 wire _22589_;
 wire _22590_;
 wire _22591_;
 wire _22592_;
 wire _22593_;
 wire _22594_;
 wire _22595_;
 wire _22596_;
 wire _22597_;
 wire _22598_;
 wire _22599_;
 wire _22600_;
 wire _22601_;
 wire _22602_;
 wire _22603_;
 wire _22604_;
 wire _22605_;
 wire _22606_;
 wire _22607_;
 wire _22608_;
 wire _22609_;
 wire _22610_;
 wire _22611_;
 wire _22612_;
 wire _22613_;
 wire _22614_;
 wire _22615_;
 wire _22616_;
 wire _22617_;
 wire _22618_;
 wire _22619_;
 wire _22620_;
 wire _22621_;
 wire _22622_;
 wire _22623_;
 wire _22624_;
 wire _22625_;
 wire _22626_;
 wire _22627_;
 wire _22628_;
 wire _22629_;
 wire _22630_;
 wire _22631_;
 wire _22632_;
 wire _22633_;
 wire _22634_;
 wire _22635_;
 wire _22636_;
 wire _22637_;
 wire _22638_;
 wire _22639_;
 wire _22640_;
 wire _22641_;
 wire _22642_;
 wire _22643_;
 wire _22644_;
 wire _22645_;
 wire _22646_;
 wire _22647_;
 wire _22648_;
 wire _22649_;
 wire _22650_;
 wire _22651_;
 wire _22652_;
 wire _22653_;
 wire _22654_;
 wire _22655_;
 wire _22656_;
 wire _22657_;
 wire _22658_;
 wire _22659_;
 wire _22660_;
 wire _22661_;
 wire _22662_;
 wire _22663_;
 wire _22664_;
 wire _22665_;
 wire _22666_;
 wire _22667_;
 wire _22668_;
 wire _22669_;
 wire _22670_;
 wire _22671_;
 wire _22672_;
 wire _22673_;
 wire _22674_;
 wire _22675_;
 wire _22676_;
 wire _22677_;
 wire _22678_;
 wire _22679_;
 wire _22680_;
 wire _22681_;
 wire _22682_;
 wire _22683_;
 wire _22684_;
 wire _22685_;
 wire _22686_;
 wire _22687_;
 wire _22688_;
 wire _22689_;
 wire _22690_;
 wire _22691_;
 wire _22692_;
 wire _22693_;
 wire _22694_;
 wire _22695_;
 wire _22696_;
 wire _22697_;
 wire _22698_;
 wire _22699_;
 wire _22700_;
 wire _22701_;
 wire _22702_;
 wire _22703_;
 wire _22704_;
 wire _22705_;
 wire _22706_;
 wire _22707_;
 wire _22708_;
 wire _22709_;
 wire _22710_;
 wire _22711_;
 wire _22712_;
 wire _22713_;
 wire _22714_;
 wire _22715_;
 wire _22716_;
 wire _22717_;
 wire _22718_;
 wire _22719_;
 wire _22720_;
 wire _22721_;
 wire _22722_;
 wire _22723_;
 wire _22724_;
 wire _22725_;
 wire _22726_;
 wire _22727_;
 wire _22728_;
 wire _22729_;
 wire _22730_;
 wire _22731_;
 wire _22732_;
 wire _22733_;
 wire _22734_;
 wire _22735_;
 wire _22736_;
 wire _22737_;
 wire _22738_;
 wire _22739_;
 wire _22740_;
 wire _22741_;
 wire _22742_;
 wire _22743_;
 wire _22744_;
 wire _22745_;
 wire _22746_;
 wire _22747_;
 wire _22748_;
 wire _22749_;
 wire _22750_;
 wire _22751_;
 wire _22752_;
 wire _22753_;
 wire _22754_;
 wire _22755_;
 wire _22756_;
 wire _22757_;
 wire _22758_;
 wire _22759_;
 wire _22760_;
 wire _22761_;
 wire _22762_;
 wire _22763_;
 wire _22764_;
 wire _22765_;
 wire _22766_;
 wire _22767_;
 wire _22768_;
 wire _22769_;
 wire _22770_;
 wire _22771_;
 wire _22772_;
 wire _22773_;
 wire _22774_;
 wire _22775_;
 wire _22776_;
 wire _22777_;
 wire _22778_;
 wire _22779_;
 wire _22780_;
 wire _22781_;
 wire _22782_;
 wire _22783_;
 wire _22784_;
 wire _22785_;
 wire _22786_;
 wire _22787_;
 wire _22788_;
 wire _22789_;
 wire _22790_;
 wire _22791_;
 wire _22792_;
 wire _22793_;
 wire _22794_;
 wire _22795_;
 wire _22796_;
 wire _22797_;
 wire _22798_;
 wire _22799_;
 wire _22800_;
 wire _22801_;
 wire _22802_;
 wire _22803_;
 wire _22804_;
 wire _22805_;
 wire _22806_;
 wire _22807_;
 wire _22808_;
 wire _22809_;
 wire _22810_;
 wire _22811_;
 wire _22812_;
 wire _22813_;
 wire _22814_;
 wire _22815_;
 wire _22816_;
 wire _22817_;
 wire _22818_;
 wire _22819_;
 wire _22820_;
 wire _22821_;
 wire _22822_;
 wire _22823_;
 wire _22824_;
 wire _22825_;
 wire _22826_;
 wire _22827_;
 wire _22828_;
 wire _22829_;
 wire _22830_;
 wire _22831_;
 wire _22832_;
 wire _22833_;
 wire _22834_;
 wire _22835_;
 wire _22836_;
 wire _22837_;
 wire _22838_;
 wire _22839_;
 wire _22840_;
 wire _22841_;
 wire _22842_;
 wire _22843_;
 wire _22844_;
 wire _22845_;
 wire _22846_;
 wire _22847_;
 wire _22848_;
 wire _22849_;
 wire _22850_;
 wire _22851_;
 wire _22852_;
 wire _22853_;
 wire _22854_;
 wire _22855_;
 wire _22856_;
 wire _22857_;
 wire _22858_;
 wire _22859_;
 wire _22860_;
 wire _22861_;
 wire _22862_;
 wire _22863_;
 wire _22864_;
 wire _22865_;
 wire _22866_;
 wire _22867_;
 wire _22868_;
 wire _22869_;
 wire _22870_;
 wire _22871_;
 wire _22872_;
 wire _22873_;
 wire _22874_;
 wire _22875_;
 wire _22876_;
 wire _22877_;
 wire _22878_;
 wire _22879_;
 wire _22880_;
 wire _22881_;
 wire _22882_;
 wire _22883_;
 wire _22884_;
 wire _22885_;
 wire _22886_;
 wire _22887_;
 wire _22888_;
 wire _22889_;
 wire _22890_;
 wire _22891_;
 wire _22892_;
 wire _22893_;
 wire _22894_;
 wire _22895_;
 wire _22896_;
 wire _22897_;
 wire _22898_;
 wire _22899_;
 wire _22900_;
 wire _22901_;
 wire _22902_;
 wire _22903_;
 wire _22904_;
 wire _22905_;
 wire _22906_;
 wire _22907_;
 wire _22908_;
 wire _22909_;
 wire _22910_;
 wire _22911_;
 wire _22912_;
 wire _22913_;
 wire _22914_;
 wire _22915_;
 wire _22916_;
 wire _22917_;
 wire _22918_;
 wire _22919_;
 wire _22920_;
 wire _22921_;
 wire _22922_;
 wire _22923_;
 wire _22924_;
 wire _22925_;
 wire _22926_;
 wire _22927_;
 wire _22928_;
 wire _22929_;
 wire _22930_;
 wire _22931_;
 wire _22932_;
 wire _22933_;
 wire _22934_;
 wire _22935_;
 wire _22936_;
 wire _22937_;
 wire _22938_;
 wire _22939_;
 wire _22940_;
 wire _22941_;
 wire _22942_;
 wire _22943_;
 wire _22944_;
 wire _22945_;
 wire _22946_;
 wire _22947_;
 wire _22948_;
 wire _22949_;
 wire _22950_;
 wire _22951_;
 wire _22952_;
 wire _22953_;
 wire _22954_;
 wire _22955_;
 wire _22956_;
 wire _22957_;
 wire _22958_;
 wire _22959_;
 wire _22960_;
 wire _22961_;
 wire _22962_;
 wire _22963_;
 wire _22964_;
 wire _22965_;
 wire _22966_;
 wire _22967_;
 wire _22968_;
 wire _22969_;
 wire _22970_;
 wire _22971_;
 wire _22972_;
 wire _22973_;
 wire _22974_;
 wire _22975_;
 wire _22976_;
 wire _22977_;
 wire _22978_;
 wire _22979_;
 wire _22980_;
 wire _22981_;
 wire _22982_;
 wire _22983_;
 wire _22984_;
 wire _22985_;
 wire _22986_;
 wire _22987_;
 wire _22988_;
 wire _22989_;
 wire _22990_;
 wire _22991_;
 wire _22992_;
 wire _22993_;
 wire _22994_;
 wire _22995_;
 wire _22996_;
 wire _22997_;
 wire _22998_;
 wire _22999_;
 wire _23000_;
 wire _23001_;
 wire _23002_;
 wire _23003_;
 wire _23004_;
 wire _23005_;
 wire _23006_;
 wire _23007_;
 wire _23008_;
 wire _23009_;
 wire _23010_;
 wire _23011_;
 wire _23012_;
 wire _23013_;
 wire _23014_;
 wire _23015_;
 wire _23016_;
 wire _23017_;
 wire _23018_;
 wire _23019_;
 wire _23020_;
 wire _23021_;
 wire _23022_;
 wire _23023_;
 wire _23024_;
 wire _23025_;
 wire _23026_;
 wire _23027_;
 wire _23028_;
 wire _23029_;
 wire _23030_;
 wire _23031_;
 wire _23032_;
 wire _23033_;
 wire _23034_;
 wire _23035_;
 wire _23036_;
 wire _23037_;
 wire _23038_;
 wire _23039_;
 wire _23040_;
 wire _23041_;
 wire _23042_;
 wire _23043_;
 wire _23044_;
 wire _23045_;
 wire _23046_;
 wire _23047_;
 wire _23048_;
 wire _23049_;
 wire _23050_;
 wire _23051_;
 wire _23052_;
 wire _23053_;
 wire _23054_;
 wire _23055_;
 wire _23056_;
 wire _23057_;
 wire _23058_;
 wire _23059_;
 wire _23060_;
 wire _23061_;
 wire _23062_;
 wire _23063_;
 wire _23064_;
 wire _23065_;
 wire _23066_;
 wire _23067_;
 wire _23068_;
 wire _23069_;
 wire _23070_;
 wire _23071_;
 wire _23072_;
 wire _23073_;
 wire _23074_;
 wire _23075_;
 wire _23076_;
 wire _23077_;
 wire _23078_;
 wire _23079_;
 wire _23080_;
 wire _23081_;
 wire _23082_;
 wire _23083_;
 wire _23084_;
 wire _23085_;
 wire _23086_;
 wire _23087_;
 wire _23088_;
 wire _23089_;
 wire _23090_;
 wire _23091_;
 wire _23092_;
 wire _23093_;
 wire _23094_;
 wire _23095_;
 wire _23096_;
 wire _23097_;
 wire _23098_;
 wire _23099_;
 wire _23100_;
 wire _23101_;
 wire _23102_;
 wire _23103_;
 wire _23104_;
 wire _23105_;
 wire _23106_;
 wire _23107_;
 wire _23108_;
 wire _23109_;
 wire _23110_;
 wire _23111_;
 wire _23112_;
 wire _23113_;
 wire _23114_;
 wire _23115_;
 wire _23116_;
 wire _23117_;
 wire _23118_;
 wire _23119_;
 wire _23120_;
 wire _23121_;
 wire _23122_;
 wire _23123_;
 wire _23124_;
 wire _23125_;
 wire _23126_;
 wire _23127_;
 wire _23128_;
 wire _23129_;
 wire _23130_;
 wire _23131_;
 wire _23132_;
 wire _23133_;
 wire _23134_;
 wire _23135_;
 wire _23136_;
 wire _23137_;
 wire _23138_;
 wire _23139_;
 wire _23140_;
 wire _23141_;
 wire _23142_;
 wire _23143_;
 wire _23144_;
 wire _23145_;
 wire _23146_;
 wire _23147_;
 wire _23148_;
 wire _23149_;
 wire _23150_;
 wire _23151_;
 wire _23152_;
 wire _23153_;
 wire _23154_;
 wire _23155_;
 wire _23156_;
 wire _23157_;
 wire _23158_;
 wire _23159_;
 wire _23160_;
 wire _23161_;
 wire _23162_;
 wire _23163_;
 wire _23164_;
 wire _23165_;
 wire _23166_;
 wire _23167_;
 wire _23168_;
 wire _23169_;
 wire _23170_;
 wire _23171_;
 wire _23172_;
 wire _23173_;
 wire _23174_;
 wire _23175_;
 wire _23176_;
 wire _23177_;
 wire _23178_;
 wire _23179_;
 wire _23180_;
 wire _23181_;
 wire _23182_;
 wire _23183_;
 wire _23184_;
 wire _23185_;
 wire _23186_;
 wire _23187_;
 wire _23188_;
 wire _23189_;
 wire _23190_;
 wire _23191_;
 wire _23192_;
 wire _23193_;
 wire _23194_;
 wire _23195_;
 wire _23196_;
 wire _23197_;
 wire _23198_;
 wire _23199_;
 wire _23200_;
 wire _23201_;
 wire _23202_;
 wire _23203_;
 wire _23204_;
 wire _23205_;
 wire _23206_;
 wire _23207_;
 wire _23208_;
 wire _23209_;
 wire _23210_;
 wire _23211_;
 wire _23212_;
 wire _23213_;
 wire _23214_;
 wire _23215_;
 wire _23216_;
 wire _23217_;
 wire _23218_;
 wire _23219_;
 wire _23220_;
 wire _23221_;
 wire _23222_;
 wire _23223_;
 wire _23224_;
 wire _23225_;
 wire _23226_;
 wire _23227_;
 wire _23228_;
 wire _23229_;
 wire _23230_;
 wire _23231_;
 wire _23232_;
 wire _23233_;
 wire _23234_;
 wire _23235_;
 wire _23236_;
 wire _23237_;
 wire _23238_;
 wire _23239_;
 wire _23240_;
 wire _23241_;
 wire _23242_;
 wire _23243_;
 wire _23244_;
 wire _23245_;
 wire _23246_;
 wire _23247_;
 wire _23248_;
 wire _23249_;
 wire _23250_;
 wire _23251_;
 wire _23252_;
 wire _23253_;
 wire _23254_;
 wire _23255_;
 wire _23256_;
 wire _23257_;
 wire _23258_;
 wire _23259_;
 wire _23260_;
 wire _23261_;
 wire _23262_;
 wire _23263_;
 wire _23264_;
 wire _23265_;
 wire _23266_;
 wire _23267_;
 wire _23268_;
 wire _23269_;
 wire _23270_;
 wire _23271_;
 wire _23272_;
 wire _23273_;
 wire _23274_;
 wire _23275_;
 wire _23276_;
 wire _23277_;
 wire _23278_;
 wire _23279_;
 wire _23280_;
 wire _23281_;
 wire _23282_;
 wire _23283_;
 wire _23284_;
 wire _23285_;
 wire _23286_;
 wire _23287_;
 wire _23288_;
 wire _23289_;
 wire _23290_;
 wire _23291_;
 wire _23292_;
 wire _23293_;
 wire _23294_;
 wire _23295_;
 wire _23296_;
 wire _23297_;
 wire _23298_;
 wire _23299_;
 wire _23300_;
 wire _23301_;
 wire _23302_;
 wire _23303_;
 wire _23304_;
 wire _23305_;
 wire _23306_;
 wire _23307_;
 wire _23308_;
 wire _23309_;
 wire _23310_;
 wire _23311_;
 wire _23312_;
 wire _23313_;
 wire _23314_;
 wire _23315_;
 wire _23316_;
 wire _23317_;
 wire _23318_;
 wire _23319_;
 wire _23320_;
 wire _23321_;
 wire _23322_;
 wire _23323_;
 wire _23324_;
 wire _23325_;
 wire _23326_;
 wire _23327_;
 wire _23328_;
 wire _23329_;
 wire _23330_;
 wire _23331_;
 wire _23332_;
 wire _23333_;
 wire _23334_;
 wire _23335_;
 wire _23336_;
 wire _23337_;
 wire _23338_;
 wire _23339_;
 wire _23340_;
 wire _23341_;
 wire _23342_;
 wire _23343_;
 wire _23344_;
 wire _23345_;
 wire _23346_;
 wire _23347_;
 wire _23348_;
 wire _23349_;
 wire _23350_;
 wire _23351_;
 wire _23352_;
 wire _23353_;
 wire _23354_;
 wire _23355_;
 wire _23356_;
 wire _23357_;
 wire _23358_;
 wire _23359_;
 wire _23360_;
 wire _23361_;
 wire _23362_;
 wire _23363_;
 wire _23364_;
 wire _23365_;
 wire _23366_;
 wire _23367_;
 wire _23368_;
 wire _23369_;
 wire _23370_;
 wire _23371_;
 wire _23372_;
 wire _23373_;
 wire _23374_;
 wire _23375_;
 wire _23376_;
 wire _23377_;
 wire _23378_;
 wire _23379_;
 wire _23380_;
 wire _23381_;
 wire _23382_;
 wire _23383_;
 wire _23384_;
 wire _23385_;
 wire _23386_;
 wire _23387_;
 wire _23388_;
 wire _23389_;
 wire _23390_;
 wire _23391_;
 wire _23392_;
 wire _23393_;
 wire _23394_;
 wire _23395_;
 wire _23396_;
 wire _23397_;
 wire _23398_;
 wire _23399_;
 wire _23400_;
 wire _23401_;
 wire _23402_;
 wire _23403_;
 wire _23404_;
 wire _23405_;
 wire _23406_;
 wire _23407_;
 wire _23408_;
 wire _23409_;
 wire _23410_;
 wire _23411_;
 wire _23412_;
 wire _23413_;
 wire _23414_;
 wire _23415_;
 wire _23416_;
 wire _23417_;
 wire _23418_;
 wire _23419_;
 wire _23420_;
 wire _23421_;
 wire _23422_;
 wire _23423_;
 wire _23424_;
 wire _23425_;
 wire _23426_;
 wire _23427_;
 wire _23428_;
 wire _23429_;
 wire _23430_;
 wire _23431_;
 wire _23432_;
 wire _23433_;
 wire _23434_;
 wire _23435_;
 wire _23436_;
 wire _23437_;
 wire _23438_;
 wire _23439_;
 wire _23440_;
 wire _23441_;
 wire _23442_;
 wire _23443_;
 wire _23444_;
 wire _23445_;
 wire _23446_;
 wire _23447_;
 wire _23448_;
 wire _23449_;
 wire _23450_;
 wire _23451_;
 wire _23452_;
 wire _23453_;
 wire _23454_;
 wire _23455_;
 wire _23456_;
 wire _23457_;
 wire _23458_;
 wire _23459_;
 wire _23460_;
 wire _23461_;
 wire _23462_;
 wire _23463_;
 wire _23464_;
 wire _23465_;
 wire _23466_;
 wire _23467_;
 wire _23468_;
 wire _23469_;
 wire _23470_;
 wire _23471_;
 wire _23472_;
 wire _23473_;
 wire _23474_;
 wire _23475_;
 wire _23476_;
 wire _23477_;
 wire _23478_;
 wire _23479_;
 wire _23480_;
 wire _23481_;
 wire _23482_;
 wire _23483_;
 wire _23484_;
 wire _23485_;
 wire _23486_;
 wire _23487_;
 wire _23488_;
 wire _23489_;
 wire _23490_;
 wire _23491_;
 wire _23492_;
 wire _23493_;
 wire _23494_;
 wire _23495_;
 wire _23496_;
 wire _23497_;
 wire _23498_;
 wire _23499_;
 wire _23500_;
 wire _23501_;
 wire _23502_;
 wire _23503_;
 wire _23504_;
 wire _23505_;
 wire _23506_;
 wire _23507_;
 wire _23508_;
 wire _23509_;
 wire _23510_;
 wire _23511_;
 wire _23512_;
 wire _23513_;
 wire _23514_;
 wire _23515_;
 wire _23516_;
 wire _23517_;
 wire _23518_;
 wire _23519_;
 wire _23520_;
 wire _23521_;
 wire _23522_;
 wire _23523_;
 wire _23524_;
 wire _23525_;
 wire _23526_;
 wire _23527_;
 wire _23528_;
 wire _23529_;
 wire _23530_;
 wire _23531_;
 wire _23532_;
 wire _23533_;
 wire _23534_;
 wire _23535_;
 wire _23536_;
 wire _23537_;
 wire _23538_;
 wire _23539_;
 wire _23540_;
 wire _23541_;
 wire _23542_;
 wire _23543_;
 wire _23544_;
 wire _23545_;
 wire _23546_;
 wire _23547_;
 wire _23548_;
 wire _23549_;
 wire _23550_;
 wire _23551_;
 wire _23552_;
 wire _23553_;
 wire _23554_;
 wire _23555_;
 wire _23556_;
 wire _23557_;
 wire _23558_;
 wire _23559_;
 wire _23560_;
 wire _23561_;
 wire _23562_;
 wire _23563_;
 wire _23564_;
 wire _23565_;
 wire _23566_;
 wire _23567_;
 wire _23568_;
 wire _23569_;
 wire _23570_;
 wire _23571_;
 wire _23572_;
 wire _23573_;
 wire _23574_;
 wire _23575_;
 wire _23576_;
 wire _23577_;
 wire _23578_;
 wire _23579_;
 wire _23580_;
 wire _23581_;
 wire _23582_;
 wire _23583_;
 wire _23584_;
 wire _23585_;
 wire _23586_;
 wire _23587_;
 wire _23588_;
 wire _23589_;
 wire _23590_;
 wire _23591_;
 wire _23592_;
 wire _23593_;
 wire _23594_;
 wire _23595_;
 wire _23596_;
 wire _23597_;
 wire _23598_;
 wire _23599_;
 wire _23600_;
 wire _23601_;
 wire _23602_;
 wire _23603_;
 wire _23604_;
 wire _23605_;
 wire _23606_;
 wire _23607_;
 wire _23608_;
 wire _23609_;
 wire _23610_;
 wire _23611_;
 wire _23612_;
 wire _23613_;
 wire _23614_;
 wire _23615_;
 wire _23616_;
 wire _23617_;
 wire _23618_;
 wire _23619_;
 wire _23620_;
 wire _23621_;
 wire _23622_;
 wire _23623_;
 wire _23624_;
 wire _23625_;
 wire _23626_;
 wire _23627_;
 wire _23628_;
 wire _23629_;
 wire _23630_;
 wire _23631_;
 wire _23632_;
 wire _23633_;
 wire _23634_;
 wire _23635_;
 wire _23636_;
 wire _23637_;
 wire _23638_;
 wire _23639_;
 wire _23640_;
 wire _23641_;
 wire _23642_;
 wire _23643_;
 wire _23644_;
 wire _23645_;
 wire _23646_;
 wire _23647_;
 wire _23648_;
 wire _23649_;
 wire _23650_;
 wire _23651_;
 wire _23652_;
 wire _23653_;
 wire _23654_;
 wire _23655_;
 wire _23656_;
 wire _23657_;
 wire _23658_;
 wire _23659_;
 wire _23660_;
 wire _23661_;
 wire _23662_;
 wire _23663_;
 wire _23664_;
 wire _23665_;
 wire _23666_;
 wire _23667_;
 wire _23668_;
 wire _23669_;
 wire _23670_;
 wire _23671_;
 wire _23672_;
 wire _23673_;
 wire _23674_;
 wire _23675_;
 wire _23676_;
 wire _23677_;
 wire _23678_;
 wire _23679_;
 wire _23680_;
 wire _23681_;
 wire _23682_;
 wire _23683_;
 wire _23684_;
 wire _23685_;
 wire _23686_;
 wire _23687_;
 wire _23688_;
 wire _23689_;
 wire _23690_;
 wire _23691_;
 wire _23692_;
 wire _23693_;
 wire _23694_;
 wire _23695_;
 wire _23696_;
 wire _23697_;
 wire _23698_;
 wire _23699_;
 wire _23700_;
 wire _23701_;
 wire _23702_;
 wire _23703_;
 wire _23704_;
 wire _23705_;
 wire _23706_;
 wire _23707_;
 wire _23708_;
 wire _23709_;
 wire _23710_;
 wire _23711_;
 wire _23712_;
 wire _23713_;
 wire _23714_;
 wire _23715_;
 wire _23716_;
 wire _23717_;
 wire _23718_;
 wire _23719_;
 wire _23720_;
 wire _23721_;
 wire _23722_;
 wire _23723_;
 wire _23724_;
 wire _23725_;
 wire _23726_;
 wire _23727_;
 wire _23728_;
 wire _23729_;
 wire _23730_;
 wire _23731_;
 wire _23732_;
 wire _23733_;
 wire _23734_;
 wire _23735_;
 wire _23736_;
 wire _23737_;
 wire _23738_;
 wire _23739_;
 wire _23740_;
 wire _23741_;
 wire _23742_;
 wire _23743_;
 wire _23744_;
 wire _23745_;
 wire _23746_;
 wire _23747_;
 wire _23748_;
 wire _23749_;
 wire _23750_;
 wire _23751_;
 wire _23752_;
 wire _23753_;
 wire _23754_;
 wire _23755_;
 wire _23756_;
 wire _23757_;
 wire _23758_;
 wire _23759_;
 wire _23760_;
 wire _23761_;
 wire _23762_;
 wire _23763_;
 wire _23764_;
 wire _23765_;
 wire _23766_;
 wire _23767_;
 wire _23768_;
 wire _23769_;
 wire _23770_;
 wire _23771_;
 wire _23772_;
 wire _23773_;
 wire _23774_;
 wire _23775_;
 wire _23776_;
 wire _23777_;
 wire _23778_;
 wire _23779_;
 wire _23780_;
 wire _23781_;
 wire _23782_;
 wire _23783_;
 wire _23784_;
 wire _23785_;
 wire _23786_;
 wire _23787_;
 wire _23788_;
 wire _23789_;
 wire _23790_;
 wire _23791_;
 wire _23792_;
 wire _23793_;
 wire _23794_;
 wire _23795_;
 wire _23796_;
 wire _23797_;
 wire _23798_;
 wire _23799_;
 wire _23800_;
 wire _23801_;
 wire _23802_;
 wire _23803_;
 wire _23804_;
 wire _23805_;
 wire _23806_;
 wire _23807_;
 wire _23808_;
 wire _23809_;
 wire _23810_;
 wire _23811_;
 wire _23812_;
 wire _23813_;
 wire _23814_;
 wire _23815_;
 wire _23816_;
 wire _23817_;
 wire _23818_;
 wire _23819_;
 wire _23820_;
 wire _23821_;
 wire _23822_;
 wire _23823_;
 wire _23824_;
 wire _23825_;
 wire _23826_;
 wire _23827_;
 wire _23828_;
 wire _23829_;
 wire _23830_;
 wire _23831_;
 wire _23832_;
 wire _23833_;
 wire _23834_;
 wire _23835_;
 wire _23836_;
 wire _23837_;
 wire _23838_;
 wire _23839_;
 wire _23840_;
 wire _23841_;
 wire _23842_;
 wire _23843_;
 wire _23844_;
 wire _23845_;
 wire _23846_;
 wire _23847_;
 wire _23848_;
 wire _23849_;
 wire _23850_;
 wire _23851_;
 wire _23852_;
 wire _23853_;
 wire _23854_;
 wire _23855_;
 wire _23856_;
 wire _23857_;
 wire _23858_;
 wire _23859_;
 wire _23860_;
 wire _23861_;
 wire _23862_;
 wire _23863_;
 wire _23864_;
 wire _23865_;
 wire _23866_;
 wire _23867_;
 wire _23868_;
 wire _23869_;
 wire _23870_;
 wire _23871_;
 wire _23872_;
 wire _23873_;
 wire _23874_;
 wire _23875_;
 wire _23876_;
 wire _23877_;
 wire _23878_;
 wire _23879_;
 wire _23880_;
 wire _23881_;
 wire _23882_;
 wire _23883_;
 wire _23884_;
 wire _23885_;
 wire _23886_;
 wire _23887_;
 wire _23888_;
 wire _23889_;
 wire _23890_;
 wire _23891_;
 wire _23892_;
 wire _23893_;
 wire _23894_;
 wire _23895_;
 wire _23896_;
 wire _23897_;
 wire _23898_;
 wire _23899_;
 wire _23900_;
 wire _23901_;
 wire _23902_;
 wire _23903_;
 wire _23904_;
 wire _23905_;
 wire _23906_;
 wire _23907_;
 wire _23908_;
 wire _23909_;
 wire _23910_;
 wire _23911_;
 wire _23912_;
 wire _23913_;
 wire _23914_;
 wire _23915_;
 wire _23916_;
 wire _23917_;
 wire _23918_;
 wire _23919_;
 wire _23920_;
 wire _23921_;
 wire _23922_;
 wire _23923_;
 wire _23924_;
 wire _23925_;
 wire _23926_;
 wire _23927_;
 wire _23928_;
 wire _23929_;
 wire _23930_;
 wire _23931_;
 wire _23932_;
 wire _23933_;
 wire _23934_;
 wire _23935_;
 wire _23936_;
 wire _23937_;
 wire _23938_;
 wire _23939_;
 wire _23940_;
 wire _23941_;
 wire _23942_;
 wire _23943_;
 wire _23944_;
 wire _23945_;
 wire _23946_;
 wire _23947_;
 wire _23948_;
 wire _23949_;
 wire _23950_;
 wire _23951_;
 wire _23952_;
 wire _23953_;
 wire _23954_;
 wire _23955_;
 wire _23956_;
 wire _23957_;
 wire _23958_;
 wire _23959_;
 wire _23960_;
 wire _23961_;
 wire _23962_;
 wire _23963_;
 wire _23964_;
 wire _23965_;
 wire _23966_;
 wire _23967_;
 wire _23968_;
 wire _23969_;
 wire _23970_;
 wire _23971_;
 wire _23972_;
 wire _23973_;
 wire _23974_;
 wire _23975_;
 wire _23976_;
 wire _23977_;
 wire _23978_;
 wire _23979_;
 wire _23980_;
 wire _23981_;
 wire _23982_;
 wire _23983_;
 wire _23984_;
 wire _23985_;
 wire _23986_;
 wire _23987_;
 wire _23988_;
 wire _23989_;
 wire _23990_;
 wire _23991_;
 wire _23992_;
 wire _23993_;
 wire _23994_;
 wire _23995_;
 wire _23996_;
 wire _23997_;
 wire _23998_;
 wire _23999_;
 wire _24000_;
 wire _24001_;
 wire _24002_;
 wire _24003_;
 wire _24004_;
 wire _24005_;
 wire _24006_;
 wire _24007_;
 wire _24008_;
 wire _24009_;
 wire _24010_;
 wire _24011_;
 wire _24012_;
 wire _24013_;
 wire _24014_;
 wire _24015_;
 wire _24016_;
 wire _24017_;
 wire _24018_;
 wire _24019_;
 wire _24020_;
 wire _24021_;
 wire _24022_;
 wire _24023_;
 wire _24024_;
 wire _24025_;
 wire _24026_;
 wire _24027_;
 wire _24028_;
 wire _24029_;
 wire _24030_;
 wire _24031_;
 wire _24032_;
 wire _24033_;
 wire _24034_;
 wire _24035_;
 wire _24036_;
 wire _24037_;
 wire _24038_;
 wire _24039_;
 wire _24040_;
 wire _24041_;
 wire _24042_;
 wire _24043_;
 wire _24044_;
 wire _24045_;
 wire _24046_;
 wire _24047_;
 wire _24048_;
 wire _24049_;
 wire _24050_;
 wire _24051_;
 wire _24052_;
 wire _24053_;
 wire _24054_;
 wire _24055_;
 wire _24056_;
 wire _24057_;
 wire _24058_;
 wire _24059_;
 wire _24060_;
 wire _24061_;
 wire _24062_;
 wire _24063_;
 wire _24064_;
 wire _24065_;
 wire _24066_;
 wire _24067_;
 wire _24068_;
 wire _24069_;
 wire _24070_;
 wire _24071_;
 wire _24072_;
 wire _24073_;
 wire _24074_;
 wire _24075_;
 wire _24076_;
 wire _24077_;
 wire _24078_;
 wire _24079_;
 wire _24080_;
 wire _24081_;
 wire _24082_;
 wire _24083_;
 wire _24084_;
 wire _24085_;
 wire _24086_;
 wire _24087_;
 wire _24088_;
 wire _24089_;
 wire _24090_;
 wire _24091_;
 wire _24092_;
 wire _24093_;
 wire _24094_;
 wire _24095_;
 wire _24096_;
 wire _24097_;
 wire _24098_;
 wire _24099_;
 wire _24100_;
 wire _24101_;
 wire _24102_;
 wire _24103_;
 wire _24104_;
 wire _24105_;
 wire _24106_;
 wire _24107_;
 wire _24108_;
 wire _24109_;
 wire _24110_;
 wire _24111_;
 wire _24112_;
 wire _24113_;
 wire _24114_;
 wire _24115_;
 wire _24116_;
 wire _24117_;
 wire _24118_;
 wire _24119_;
 wire _24120_;
 wire _24121_;
 wire _24122_;
 wire _24123_;
 wire _24124_;
 wire _24125_;
 wire _24126_;
 wire _24127_;
 wire _24128_;
 wire _24129_;
 wire _24130_;
 wire _24131_;
 wire _24132_;
 wire _24133_;
 wire _24134_;
 wire _24135_;
 wire _24136_;
 wire _24137_;
 wire _24138_;
 wire _24139_;
 wire _24140_;
 wire _24141_;
 wire _24142_;
 wire _24143_;
 wire _24144_;
 wire _24145_;
 wire _24146_;
 wire _24147_;
 wire _24148_;
 wire _24149_;
 wire _24150_;
 wire _24151_;
 wire _24152_;
 wire _24153_;
 wire _24154_;
 wire _24155_;
 wire _24156_;
 wire _24157_;
 wire _24158_;
 wire _24159_;
 wire _24160_;
 wire _24161_;
 wire _24162_;
 wire _24163_;
 wire _24164_;
 wire _24165_;
 wire _24166_;
 wire _24167_;
 wire _24168_;
 wire _24169_;
 wire _24170_;
 wire _24171_;
 wire _24172_;
 wire _24173_;
 wire _24174_;
 wire _24175_;
 wire _24176_;
 wire _24177_;
 wire _24178_;
 wire _24179_;
 wire _24180_;
 wire _24181_;
 wire _24182_;
 wire _24183_;
 wire _24184_;
 wire _24185_;
 wire _24186_;
 wire _24187_;
 wire _24188_;
 wire _24189_;
 wire _24190_;
 wire _24191_;
 wire _24192_;
 wire _24193_;
 wire _24194_;
 wire _24195_;
 wire _24196_;
 wire _24197_;
 wire _24198_;
 wire _24199_;
 wire _24200_;
 wire _24201_;
 wire _24202_;
 wire _24203_;
 wire _24204_;
 wire _24205_;
 wire _24206_;
 wire _24207_;
 wire _24208_;
 wire _24209_;
 wire _24210_;
 wire _24211_;
 wire _24212_;
 wire _24213_;
 wire _24214_;
 wire _24215_;
 wire _24216_;
 wire _24217_;
 wire _24218_;
 wire _24219_;
 wire _24220_;
 wire _24221_;
 wire _24222_;
 wire _24223_;
 wire _24224_;
 wire _24225_;
 wire _24226_;
 wire _24227_;
 wire _24228_;
 wire _24229_;
 wire _24230_;
 wire _24231_;
 wire _24232_;
 wire _24233_;
 wire _24234_;
 wire _24235_;
 wire _24236_;
 wire _24237_;
 wire _24238_;
 wire _24239_;
 wire _24240_;
 wire _24241_;
 wire _24242_;
 wire _24243_;
 wire _24244_;
 wire _24245_;
 wire _24246_;
 wire _24247_;
 wire _24248_;
 wire _24249_;
 wire _24250_;
 wire _24251_;
 wire _24252_;
 wire _24253_;
 wire _24254_;
 wire _24255_;
 wire _24256_;
 wire _24257_;
 wire _24258_;
 wire _24259_;
 wire _24260_;
 wire _24261_;
 wire _24262_;
 wire _24263_;
 wire _24264_;
 wire _24265_;
 wire _24266_;
 wire _24267_;
 wire _24268_;
 wire _24269_;
 wire _24270_;
 wire _24271_;
 wire _24272_;
 wire _24273_;
 wire _24274_;
 wire _24275_;
 wire _24276_;
 wire _24277_;
 wire _24278_;
 wire _24279_;
 wire _24280_;
 wire _24281_;
 wire _24282_;
 wire _24283_;
 wire _24284_;
 wire _24285_;
 wire _24286_;
 wire _24287_;
 wire _24288_;
 wire _24289_;
 wire _24290_;
 wire _24291_;
 wire _24292_;
 wire _24293_;
 wire _24294_;
 wire _24295_;
 wire _24296_;
 wire _24297_;
 wire _24298_;
 wire _24299_;
 wire _24300_;
 wire _24301_;
 wire _24302_;
 wire _24303_;
 wire _24304_;
 wire _24305_;
 wire _24306_;
 wire _24307_;
 wire _24308_;
 wire _24309_;
 wire _24310_;
 wire _24311_;
 wire _24312_;
 wire _24313_;
 wire _24314_;
 wire _24315_;
 wire _24316_;
 wire _24317_;
 wire _24318_;
 wire _24319_;
 wire _24320_;
 wire _24321_;
 wire _24322_;
 wire _24323_;
 wire _24324_;
 wire _24325_;
 wire _24326_;
 wire _24327_;
 wire _24328_;
 wire _24329_;
 wire _24330_;
 wire _24331_;
 wire _24332_;
 wire _24333_;
 wire _24334_;
 wire _24335_;
 wire _24336_;
 wire _24337_;
 wire _24338_;
 wire _24339_;
 wire _24340_;
 wire _24341_;
 wire _24342_;
 wire _24343_;
 wire _24344_;
 wire _24345_;
 wire _24346_;
 wire _24347_;
 wire _24348_;
 wire _24349_;
 wire _24350_;
 wire _24351_;
 wire _24352_;
 wire _24353_;
 wire _24354_;
 wire _24355_;
 wire _24356_;
 wire _24357_;
 wire _24358_;
 wire _24359_;
 wire _24360_;
 wire _24361_;
 wire _24362_;
 wire _24363_;
 wire _24364_;
 wire _24365_;
 wire _24366_;
 wire _24367_;
 wire _24368_;
 wire _24369_;
 wire _24370_;
 wire _24371_;
 wire _24372_;
 wire _24373_;
 wire _24374_;
 wire _24375_;
 wire _24376_;
 wire _24377_;
 wire _24378_;
 wire _24379_;
 wire _24380_;
 wire _24381_;
 wire _24382_;
 wire _24383_;
 wire _24384_;
 wire _24385_;
 wire _24386_;
 wire _24387_;
 wire _24388_;
 wire _24389_;
 wire _24390_;
 wire _24391_;
 wire _24392_;
 wire _24393_;
 wire _24394_;
 wire _24395_;
 wire _24396_;
 wire _24397_;
 wire _24398_;
 wire _24399_;
 wire _24400_;
 wire _24401_;
 wire _24402_;
 wire _24403_;
 wire _24404_;
 wire _24405_;
 wire _24406_;
 wire _24407_;
 wire _24408_;
 wire _24409_;
 wire _24410_;
 wire _24411_;
 wire _24412_;
 wire _24413_;
 wire _24414_;
 wire _24415_;
 wire _24416_;
 wire _24417_;
 wire _24418_;
 wire _24419_;
 wire _24420_;
 wire _24421_;
 wire _24422_;
 wire _24423_;
 wire _24424_;
 wire _24425_;
 wire _24426_;
 wire _24427_;
 wire _24428_;
 wire _24429_;
 wire _24430_;
 wire _24431_;
 wire _24432_;
 wire _24433_;
 wire _24434_;
 wire _24435_;
 wire _24436_;
 wire _24437_;
 wire _24438_;
 wire _24439_;
 wire _24440_;
 wire _24441_;
 wire _24442_;
 wire _24443_;
 wire _24444_;
 wire _24445_;
 wire _24446_;
 wire _24447_;
 wire _24448_;
 wire _24449_;
 wire _24450_;
 wire _24451_;
 wire _24452_;
 wire _24453_;
 wire _24454_;
 wire _24455_;
 wire _24456_;
 wire _24457_;
 wire _24458_;
 wire _24459_;
 wire _24460_;
 wire _24461_;
 wire _24462_;
 wire _24463_;
 wire _24464_;
 wire _24465_;
 wire _24466_;
 wire _24467_;
 wire _24468_;
 wire _24469_;
 wire _24470_;
 wire _24471_;
 wire _24472_;
 wire _24473_;
 wire _24474_;
 wire _24475_;
 wire _24476_;
 wire _24477_;
 wire _24478_;
 wire _24479_;
 wire _24480_;
 wire _24481_;
 wire _24482_;
 wire _24483_;
 wire _24484_;
 wire _24485_;
 wire _24486_;
 wire _24487_;
 wire _24488_;
 wire _24489_;
 wire _24490_;
 wire _24491_;
 wire _24492_;
 wire _24493_;
 wire _24494_;
 wire _24495_;
 wire _24496_;
 wire _24497_;
 wire _24498_;
 wire _24499_;
 wire _24500_;
 wire _24501_;
 wire _24502_;
 wire _24503_;
 wire _24504_;
 wire _24505_;
 wire _24506_;
 wire _24507_;
 wire _24508_;
 wire _24509_;
 wire _24510_;
 wire _24511_;
 wire _24512_;
 wire _24513_;
 wire _24514_;
 wire _24515_;
 wire _24516_;
 wire _24517_;
 wire _24518_;
 wire _24519_;
 wire _24520_;
 wire _24521_;
 wire _24522_;
 wire _24523_;
 wire _24524_;
 wire _24525_;
 wire _24526_;
 wire _24527_;
 wire _24528_;
 wire _24529_;
 wire _24530_;
 wire _24531_;
 wire _24532_;
 wire _24533_;
 wire _24534_;
 wire _24535_;
 wire _24536_;
 wire _24537_;
 wire _24538_;
 wire _24539_;
 wire _24540_;
 wire _24541_;
 wire _24542_;
 wire _24543_;
 wire _24544_;
 wire _24545_;
 wire _24546_;
 wire _24547_;
 wire _24548_;
 wire _24549_;
 wire _24550_;
 wire _24551_;
 wire _24552_;
 wire _24553_;
 wire _24554_;
 wire _24555_;
 wire _24556_;
 wire _24557_;
 wire _24558_;
 wire _24559_;
 wire _24560_;
 wire _24561_;
 wire _24562_;
 wire _24563_;
 wire _24564_;
 wire _24565_;
 wire _24566_;
 wire _24567_;
 wire _24568_;
 wire _24569_;
 wire _24570_;
 wire _24571_;
 wire _24572_;
 wire _24573_;
 wire _24574_;
 wire _24575_;
 wire _24576_;
 wire _24577_;
 wire _24578_;
 wire _24579_;
 wire _24580_;
 wire _24581_;
 wire _24582_;
 wire _24583_;
 wire _24584_;
 wire _24585_;
 wire _24586_;
 wire _24587_;
 wire _24588_;
 wire _24589_;
 wire _24590_;
 wire _24591_;
 wire _24592_;
 wire _24593_;
 wire _24594_;
 wire _24595_;
 wire _24596_;
 wire _24597_;
 wire _24598_;
 wire _24599_;
 wire _24600_;
 wire _24601_;
 wire _24602_;
 wire _24603_;
 wire _24604_;
 wire _24605_;
 wire _24606_;
 wire _24607_;
 wire _24608_;
 wire _24609_;
 wire _24610_;
 wire _24611_;
 wire _24612_;
 wire _24613_;
 wire _24614_;
 wire _24615_;
 wire _24616_;
 wire _24617_;
 wire _24618_;
 wire _24619_;
 wire _24620_;
 wire _24621_;
 wire _24622_;
 wire _24623_;
 wire _24624_;
 wire _24625_;
 wire _24626_;
 wire _24627_;
 wire _24628_;
 wire _24629_;
 wire _24630_;
 wire _24631_;
 wire _24632_;
 wire _24633_;
 wire _24634_;
 wire _24635_;
 wire _24636_;
 wire _24637_;
 wire _24638_;
 wire _24639_;
 wire _24640_;
 wire _24641_;
 wire _24642_;
 wire _24643_;
 wire _24644_;
 wire _24645_;
 wire _24646_;
 wire _24647_;
 wire _24648_;
 wire _24649_;
 wire _24650_;
 wire _24651_;
 wire _24652_;
 wire _24653_;
 wire _24654_;
 wire _24655_;
 wire _24656_;
 wire _24657_;
 wire _24658_;
 wire _24659_;
 wire _24660_;
 wire _24661_;
 wire _24662_;
 wire _24663_;
 wire _24664_;
 wire _24665_;
 wire _24666_;
 wire _24667_;
 wire _24668_;
 wire _24669_;
 wire _24670_;
 wire _24671_;
 wire _24672_;
 wire _24673_;
 wire _24674_;
 wire _24675_;
 wire _24676_;
 wire _24677_;
 wire _24678_;
 wire _24679_;
 wire _24680_;
 wire _24681_;
 wire _24682_;
 wire _24683_;
 wire _24684_;
 wire _24685_;
 wire _24686_;
 wire _24687_;
 wire _24688_;
 wire _24689_;
 wire _24690_;
 wire _24691_;
 wire _24692_;
 wire _24693_;
 wire _24694_;
 wire _24695_;
 wire _24696_;
 wire _24697_;
 wire _24698_;
 wire _24699_;
 wire _24700_;
 wire _24701_;
 wire _24702_;
 wire _24703_;
 wire _24704_;
 wire _24705_;
 wire _24706_;
 wire _24707_;
 wire _24708_;
 wire _24709_;
 wire _24710_;
 wire _24711_;
 wire _24712_;
 wire _24713_;
 wire _24714_;
 wire _24715_;
 wire _24716_;
 wire _24717_;
 wire _24718_;
 wire _24719_;
 wire _24720_;
 wire _24721_;
 wire _24722_;
 wire _24723_;
 wire _24724_;
 wire _24725_;
 wire _24726_;
 wire _24727_;
 wire _24728_;
 wire _24729_;
 wire _24730_;
 wire _24731_;
 wire _24732_;
 wire _24733_;
 wire _24734_;
 wire _24735_;
 wire _24736_;
 wire _24737_;
 wire _24738_;
 wire _24739_;
 wire _24740_;
 wire _24741_;
 wire _24742_;
 wire _24743_;
 wire _24744_;
 wire _24745_;
 wire _24746_;
 wire _24747_;
 wire _24748_;
 wire _24749_;
 wire _24750_;
 wire _24751_;
 wire _24752_;
 wire _24753_;
 wire _24754_;
 wire _24755_;
 wire _24756_;
 wire _24757_;
 wire _24758_;
 wire _24759_;
 wire _24760_;
 wire _24761_;
 wire _24762_;
 wire _24763_;
 wire _24764_;
 wire _24765_;
 wire _24766_;
 wire _24767_;
 wire _24768_;
 wire _24769_;
 wire _24770_;
 wire _24771_;
 wire _24772_;
 wire _24773_;
 wire _24774_;
 wire _24775_;
 wire _24776_;
 wire _24777_;
 wire _24778_;
 wire _24779_;
 wire _24780_;
 wire _24781_;
 wire _24782_;
 wire _24783_;
 wire _24784_;
 wire _24785_;
 wire _24786_;
 wire _24787_;
 wire _24788_;
 wire _24789_;
 wire _24790_;
 wire _24791_;
 wire _24792_;
 wire _24793_;
 wire _24794_;
 wire _24795_;
 wire _24796_;
 wire _24797_;
 wire _24798_;
 wire _24799_;
 wire _24800_;
 wire _24801_;
 wire _24802_;
 wire _24803_;
 wire _24804_;
 wire _24805_;
 wire _24806_;
 wire _24807_;
 wire _24808_;
 wire _24809_;
 wire _24810_;
 wire _24811_;
 wire _24812_;
 wire _24813_;
 wire _24814_;
 wire _24815_;
 wire _24816_;
 wire _24817_;
 wire _24818_;
 wire _24819_;
 wire _24820_;
 wire _24821_;
 wire _24822_;
 wire _24823_;
 wire _24824_;
 wire _24825_;
 wire _24826_;
 wire _24827_;
 wire _24828_;
 wire _24829_;
 wire _24830_;
 wire _24831_;
 wire _24832_;
 wire _24833_;
 wire _24834_;
 wire _24835_;
 wire _24836_;
 wire _24837_;
 wire _24838_;
 wire _24839_;
 wire _24840_;
 wire _24841_;
 wire _24842_;
 wire _24843_;
 wire _24844_;
 wire _24845_;
 wire _24846_;
 wire _24847_;
 wire _24848_;
 wire _24849_;
 wire _24850_;
 wire _24851_;
 wire _24852_;
 wire _24853_;
 wire _24854_;
 wire _24855_;
 wire _24856_;
 wire _24857_;
 wire _24858_;
 wire _24859_;
 wire _24860_;
 wire _24861_;
 wire _24862_;
 wire _24863_;
 wire _24864_;
 wire _24865_;
 wire _24866_;
 wire _24867_;
 wire _24868_;
 wire _24869_;
 wire _24870_;
 wire _24871_;
 wire _24872_;
 wire _24873_;
 wire _24874_;
 wire _24875_;
 wire _24876_;
 wire _24877_;
 wire _24878_;
 wire _24879_;
 wire _24880_;
 wire _24881_;
 wire _24882_;
 wire _24883_;
 wire _24884_;
 wire _24885_;
 wire _24886_;
 wire _24887_;
 wire _24888_;
 wire _24889_;
 wire _24890_;
 wire _24891_;
 wire _24892_;
 wire _24893_;
 wire _24894_;
 wire _24895_;
 wire _24896_;
 wire _24897_;
 wire _24898_;
 wire _24899_;
 wire _24900_;
 wire _24901_;
 wire _24902_;
 wire _24903_;
 wire _24904_;
 wire _24905_;
 wire _24906_;
 wire _24907_;
 wire _24908_;
 wire _24909_;
 wire _24910_;
 wire _24911_;
 wire _24912_;
 wire _24913_;
 wire _24914_;
 wire _24915_;
 wire _24916_;
 wire _24917_;
 wire _24918_;
 wire _24919_;
 wire _24920_;
 wire _24921_;
 wire _24922_;
 wire _24923_;
 wire _24924_;
 wire _24925_;
 wire _24926_;
 wire _24927_;
 wire _24928_;
 wire _24929_;
 wire _24930_;
 wire _24931_;
 wire _24932_;
 wire _24933_;
 wire _24934_;
 wire _24935_;
 wire _24936_;
 wire _24937_;
 wire _24938_;
 wire _24939_;
 wire _24940_;
 wire _24941_;
 wire _24942_;
 wire _24943_;
 wire _24944_;
 wire _24945_;
 wire _24946_;
 wire _24947_;
 wire _24948_;
 wire _24949_;
 wire _24950_;
 wire _24951_;
 wire _24952_;
 wire _24953_;
 wire _24954_;
 wire _24955_;
 wire _24956_;
 wire _24957_;
 wire _24958_;
 wire _24959_;
 wire _24960_;
 wire _24961_;
 wire _24962_;
 wire _24963_;
 wire _24964_;
 wire _24965_;
 wire _24966_;
 wire _24967_;
 wire _24968_;
 wire _24969_;
 wire _24970_;
 wire _24971_;
 wire _24972_;
 wire _24973_;
 wire _24974_;
 wire _24975_;
 wire _24976_;
 wire _24977_;
 wire _24978_;
 wire _24979_;
 wire _24980_;
 wire _24981_;
 wire _24982_;
 wire _24983_;
 wire _24984_;
 wire _24985_;
 wire _24986_;
 wire _24987_;
 wire _24988_;
 wire _24989_;
 wire _24990_;
 wire _24991_;
 wire _24992_;
 wire _24993_;
 wire _24994_;
 wire _24995_;
 wire _24996_;
 wire _24997_;
 wire _24998_;
 wire _24999_;
 wire _25000_;
 wire _25001_;
 wire _25002_;
 wire _25003_;
 wire _25004_;
 wire _25005_;
 wire _25006_;
 wire _25007_;
 wire _25008_;
 wire _25009_;
 wire _25010_;
 wire _25011_;
 wire _25012_;
 wire _25013_;
 wire _25014_;
 wire _25015_;
 wire _25016_;
 wire _25017_;
 wire _25018_;
 wire _25019_;
 wire _25020_;
 wire _25021_;
 wire _25022_;
 wire _25023_;
 wire _25024_;
 wire _25025_;
 wire _25026_;
 wire _25027_;
 wire _25028_;
 wire _25029_;
 wire _25030_;
 wire _25031_;
 wire _25032_;
 wire _25033_;
 wire _25034_;
 wire _25035_;
 wire _25036_;
 wire _25037_;
 wire _25038_;
 wire _25039_;
 wire _25040_;
 wire _25041_;
 wire _25042_;
 wire _25043_;
 wire _25044_;
 wire _25045_;
 wire _25046_;
 wire _25047_;
 wire _25048_;
 wire _25049_;
 wire _25050_;
 wire _25051_;
 wire _25052_;
 wire _25053_;
 wire _25054_;
 wire _25055_;
 wire _25056_;
 wire _25057_;
 wire _25058_;
 wire _25059_;
 wire _25060_;
 wire _25061_;
 wire _25062_;
 wire _25063_;
 wire _25064_;
 wire _25065_;
 wire _25066_;
 wire _25067_;
 wire _25068_;
 wire _25069_;
 wire _25070_;
 wire _25071_;
 wire _25072_;
 wire _25073_;
 wire _25074_;
 wire _25075_;
 wire _25076_;
 wire _25077_;
 wire _25078_;
 wire _25079_;
 wire _25080_;
 wire _25081_;
 wire _25082_;
 wire _25083_;
 wire _25084_;
 wire _25085_;
 wire _25086_;
 wire _25087_;
 wire _25088_;
 wire _25089_;
 wire _25090_;
 wire _25091_;
 wire _25092_;
 wire _25093_;
 wire _25094_;
 wire _25095_;
 wire _25096_;
 wire _25097_;
 wire _25098_;
 wire _25099_;
 wire _25100_;
 wire _25101_;
 wire _25102_;
 wire _25103_;
 wire _25104_;
 wire _25105_;
 wire _25106_;
 wire _25107_;
 wire _25108_;
 wire _25109_;
 wire _25110_;
 wire _25111_;
 wire _25112_;
 wire _25113_;
 wire _25114_;
 wire _25115_;
 wire _25116_;
 wire _25117_;
 wire _25118_;
 wire _25119_;
 wire _25120_;
 wire _25121_;
 wire _25122_;
 wire _25123_;
 wire _25124_;
 wire _25125_;
 wire _25126_;
 wire _25127_;
 wire _25128_;
 wire _25129_;
 wire _25130_;
 wire _25131_;
 wire _25132_;
 wire _25133_;
 wire _25134_;
 wire _25135_;
 wire _25136_;
 wire _25137_;
 wire _25138_;
 wire _25139_;
 wire _25140_;
 wire _25141_;
 wire _25142_;
 wire _25143_;
 wire _25144_;
 wire _25145_;
 wire _25146_;
 wire _25147_;
 wire _25148_;
 wire _25149_;
 wire _25150_;
 wire _25151_;
 wire _25152_;
 wire _25153_;
 wire _25154_;
 wire _25155_;
 wire _25156_;
 wire _25157_;
 wire _25158_;
 wire _25159_;
 wire _25160_;
 wire _25161_;
 wire _25162_;
 wire _25163_;
 wire _25164_;
 wire _25165_;
 wire _25166_;
 wire _25167_;
 wire _25168_;
 wire _25169_;
 wire _25170_;
 wire _25171_;
 wire _25172_;
 wire _25173_;
 wire _25174_;
 wire _25175_;
 wire _25176_;
 wire _25177_;
 wire _25178_;
 wire _25179_;
 wire _25180_;
 wire _25181_;
 wire _25182_;
 wire _25183_;
 wire _25184_;
 wire _25185_;
 wire _25186_;
 wire _25187_;
 wire _25188_;
 wire _25189_;
 wire _25190_;
 wire _25191_;
 wire _25192_;
 wire _25193_;
 wire _25194_;
 wire _25195_;
 wire _25196_;
 wire _25197_;
 wire _25198_;
 wire _25199_;
 wire _25200_;
 wire _25201_;
 wire _25202_;
 wire _25203_;
 wire _25204_;
 wire _25205_;
 wire _25206_;
 wire _25207_;
 wire _25208_;
 wire _25209_;
 wire _25210_;
 wire _25211_;
 wire _25212_;
 wire _25213_;
 wire _25214_;
 wire _25215_;
 wire _25216_;
 wire _25217_;
 wire _25218_;
 wire _25219_;
 wire _25220_;
 wire _25221_;
 wire _25222_;
 wire _25223_;
 wire _25224_;
 wire _25225_;
 wire _25226_;
 wire _25227_;
 wire _25228_;
 wire _25229_;
 wire _25230_;
 wire _25231_;
 wire _25232_;
 wire _25233_;
 wire _25234_;
 wire _25235_;
 wire _25236_;
 wire _25237_;
 wire _25238_;
 wire _25239_;
 wire _25240_;
 wire _25241_;
 wire _25242_;
 wire _25243_;
 wire _25244_;
 wire _25245_;
 wire _25246_;
 wire _25247_;
 wire _25248_;
 wire _25249_;
 wire _25250_;
 wire _25251_;
 wire _25252_;
 wire _25253_;
 wire _25254_;
 wire _25255_;
 wire _25256_;
 wire _25257_;
 wire _25258_;
 wire _25259_;
 wire _25260_;
 wire _25261_;
 wire _25262_;
 wire _25263_;
 wire _25264_;
 wire _25265_;
 wire _25266_;
 wire _25267_;
 wire _25268_;
 wire _25269_;
 wire _25270_;
 wire _25271_;
 wire _25272_;
 wire _25273_;
 wire _25274_;
 wire _25275_;
 wire _25276_;
 wire _25277_;
 wire _25278_;
 wire _25279_;
 wire _25280_;
 wire _25281_;
 wire _25282_;
 wire _25283_;
 wire _25284_;
 wire _25285_;
 wire _25286_;
 wire _25287_;
 wire _25288_;
 wire _25289_;
 wire _25290_;
 wire _25291_;
 wire _25292_;
 wire _25293_;
 wire _25294_;
 wire _25295_;
 wire _25296_;
 wire _25297_;
 wire _25298_;
 wire _25299_;
 wire _25300_;
 wire _25301_;
 wire _25302_;
 wire _25303_;
 wire _25304_;
 wire _25305_;
 wire _25306_;
 wire _25307_;
 wire _25308_;
 wire _25309_;
 wire _25310_;
 wire _25311_;
 wire _25312_;
 wire _25313_;
 wire _25314_;
 wire _25315_;
 wire _25316_;
 wire _25317_;
 wire _25318_;
 wire _25319_;
 wire _25320_;
 wire _25321_;
 wire _25322_;
 wire _25323_;
 wire _25324_;
 wire _25325_;
 wire _25326_;
 wire _25327_;
 wire _25328_;
 wire _25329_;
 wire _25330_;
 wire _25331_;
 wire _25332_;
 wire _25333_;
 wire _25334_;
 wire _25335_;
 wire _25336_;
 wire _25337_;
 wire _25338_;
 wire _25339_;
 wire _25340_;
 wire _25341_;
 wire _25342_;
 wire _25343_;
 wire _25344_;
 wire _25345_;
 wire _25346_;
 wire _25347_;
 wire _25348_;
 wire _25349_;
 wire _25350_;
 wire _25351_;
 wire _25352_;
 wire _25353_;
 wire _25354_;
 wire _25355_;
 wire _25356_;
 wire _25357_;
 wire _25358_;
 wire _25359_;
 wire _25360_;
 wire _25361_;
 wire _25362_;
 wire _25363_;
 wire _25364_;
 wire _25365_;
 wire _25366_;
 wire _25367_;
 wire _25368_;
 wire _25369_;
 wire _25370_;
 wire _25371_;
 wire _25372_;
 wire _25373_;
 wire _25374_;
 wire _25375_;
 wire _25376_;
 wire _25377_;
 wire _25378_;
 wire _25379_;
 wire _25380_;
 wire _25381_;
 wire _25382_;
 wire _25383_;
 wire _25384_;
 wire _25385_;
 wire _25386_;
 wire _25387_;
 wire _25388_;
 wire _25389_;
 wire _25390_;
 wire _25391_;
 wire _25392_;
 wire _25393_;
 wire _25394_;
 wire _25395_;
 wire _25396_;
 wire _25397_;
 wire _25398_;
 wire _25399_;
 wire _25400_;
 wire _25401_;
 wire _25402_;
 wire _25403_;
 wire _25404_;
 wire _25405_;
 wire _25406_;
 wire _25407_;
 wire _25408_;
 wire _25409_;
 wire _25410_;
 wire _25411_;
 wire _25412_;
 wire _25413_;
 wire _25414_;
 wire _25415_;
 wire _25416_;
 wire _25417_;
 wire _25418_;
 wire _25419_;
 wire _25420_;
 wire _25421_;
 wire _25422_;
 wire _25423_;
 wire _25424_;
 wire _25425_;
 wire _25426_;
 wire _25427_;
 wire _25428_;
 wire _25429_;
 wire _25430_;
 wire _25431_;
 wire _25432_;
 wire _25433_;
 wire _25434_;
 wire _25435_;
 wire _25436_;
 wire _25437_;
 wire _25438_;
 wire _25439_;
 wire _25440_;
 wire _25441_;
 wire _25442_;
 wire _25443_;
 wire _25444_;
 wire _25445_;
 wire _25446_;
 wire _25447_;
 wire _25448_;
 wire _25449_;
 wire _25450_;
 wire _25451_;
 wire _25452_;
 wire _25453_;
 wire _25454_;
 wire _25455_;
 wire _25456_;
 wire _25457_;
 wire _25458_;
 wire _25459_;
 wire _25460_;
 wire _25461_;
 wire _25462_;
 wire _25463_;
 wire _25464_;
 wire _25465_;
 wire _25466_;
 wire _25467_;
 wire _25468_;
 wire _25469_;
 wire _25470_;
 wire _25471_;
 wire _25472_;
 wire _25473_;
 wire _25474_;
 wire _25475_;
 wire _25476_;
 wire _25477_;
 wire _25478_;
 wire _25479_;
 wire _25480_;
 wire _25481_;
 wire _25482_;
 wire _25483_;
 wire _25484_;
 wire _25485_;
 wire _25486_;
 wire _25487_;
 wire _25488_;
 wire _25489_;
 wire _25490_;
 wire _25491_;
 wire _25492_;
 wire _25493_;
 wire _25494_;
 wire _25495_;
 wire _25496_;
 wire _25497_;
 wire _25498_;
 wire _25499_;
 wire _25500_;
 wire _25501_;
 wire _25502_;
 wire _25503_;
 wire _25504_;
 wire _25505_;
 wire _25506_;
 wire _25507_;
 wire _25508_;
 wire _25509_;
 wire _25510_;
 wire _25511_;
 wire _25512_;
 wire _25513_;
 wire _25514_;
 wire _25515_;
 wire _25516_;
 wire _25517_;
 wire _25518_;
 wire _25519_;
 wire _25520_;
 wire _25521_;
 wire _25522_;
 wire _25523_;
 wire _25524_;
 wire _25525_;
 wire _25526_;
 wire _25527_;
 wire _25528_;
 wire _25529_;
 wire _25530_;
 wire _25531_;
 wire _25532_;
 wire _25533_;
 wire _25534_;
 wire _25535_;
 wire _25536_;
 wire _25537_;
 wire _25538_;
 wire _25539_;
 wire _25540_;
 wire _25541_;
 wire _25542_;
 wire _25543_;
 wire _25544_;
 wire _25545_;
 wire _25546_;
 wire _25547_;
 wire _25548_;
 wire _25549_;
 wire _25550_;
 wire _25551_;
 wire _25552_;
 wire _25553_;
 wire _25554_;
 wire _25555_;
 wire _25556_;
 wire _25557_;
 wire _25558_;
 wire _25559_;
 wire _25560_;
 wire _25561_;
 wire _25562_;
 wire _25563_;
 wire _25564_;
 wire _25565_;
 wire _25566_;
 wire _25567_;
 wire _25568_;
 wire _25569_;
 wire _25570_;
 wire _25571_;
 wire _25572_;
 wire _25573_;
 wire _25574_;
 wire _25575_;
 wire _25576_;
 wire _25577_;
 wire _25578_;
 wire _25579_;
 wire _25580_;
 wire _25581_;
 wire _25582_;
 wire _25583_;
 wire _25584_;
 wire _25585_;
 wire _25586_;
 wire _25587_;
 wire _25588_;
 wire _25589_;
 wire _25590_;
 wire _25591_;
 wire _25592_;
 wire _25593_;
 wire _25594_;
 wire _25595_;
 wire _25596_;
 wire _25597_;
 wire _25598_;
 wire _25599_;
 wire _25600_;
 wire _25601_;
 wire _25602_;
 wire _25603_;
 wire _25604_;
 wire _25605_;
 wire _25606_;
 wire _25607_;
 wire _25608_;
 wire _25609_;
 wire _25610_;
 wire _25611_;
 wire _25612_;
 wire _25613_;
 wire _25614_;
 wire _25615_;
 wire _25616_;
 wire _25617_;
 wire _25618_;
 wire _25619_;
 wire _25620_;
 wire _25621_;
 wire _25622_;
 wire _25623_;
 wire _25624_;
 wire _25625_;
 wire _25626_;
 wire _25627_;
 wire _25628_;
 wire _25629_;
 wire _25630_;
 wire _25631_;
 wire _25632_;
 wire _25633_;
 wire _25634_;
 wire _25635_;
 wire _25636_;
 wire _25637_;
 wire _25638_;
 wire _25639_;
 wire _25640_;
 wire _25641_;
 wire _25642_;
 wire _25643_;
 wire _25644_;
 wire _25645_;
 wire _25646_;
 wire _25647_;
 wire _25648_;
 wire _25649_;
 wire _25650_;
 wire _25651_;
 wire _25652_;
 wire _25653_;
 wire _25654_;
 wire _25655_;
 wire _25656_;
 wire _25657_;
 wire _25658_;
 wire _25659_;
 wire _25660_;
 wire _25661_;
 wire _25662_;
 wire _25663_;
 wire _25664_;
 wire _25665_;
 wire _25666_;
 wire _25667_;
 wire _25668_;
 wire _25669_;
 wire _25670_;
 wire _25671_;
 wire _25672_;
 wire _25673_;
 wire _25674_;
 wire _25675_;
 wire _25676_;
 wire _25677_;
 wire _25678_;
 wire _25679_;
 wire _25680_;
 wire _25681_;
 wire _25682_;
 wire _25683_;
 wire _25684_;
 wire _25685_;
 wire _25686_;
 wire _25687_;
 wire _25688_;
 wire _25689_;
 wire _25690_;
 wire _25691_;
 wire _25692_;
 wire _25693_;
 wire _25694_;
 wire _25695_;
 wire _25696_;
 wire _25697_;
 wire _25698_;
 wire _25699_;
 wire _25700_;
 wire _25701_;
 wire _25702_;
 wire _25703_;
 wire _25704_;
 wire _25705_;
 wire _25706_;
 wire _25707_;
 wire _25708_;
 wire _25709_;
 wire _25710_;
 wire _25711_;
 wire _25712_;
 wire _25713_;
 wire _25714_;
 wire _25715_;
 wire _25716_;
 wire _25717_;
 wire _25718_;
 wire _25719_;
 wire _25720_;
 wire _25721_;
 wire _25722_;
 wire _25723_;
 wire _25724_;
 wire _25725_;
 wire _25726_;
 wire _25727_;
 wire _25728_;
 wire _25729_;
 wire _25730_;
 wire _25731_;
 wire _25732_;
 wire _25733_;
 wire _25734_;
 wire _25735_;
 wire _25736_;
 wire _25737_;
 wire _25738_;
 wire _25739_;
 wire _25740_;
 wire _25741_;
 wire _25742_;
 wire _25743_;
 wire _25744_;
 wire _25745_;
 wire _25746_;
 wire _25747_;
 wire _25748_;
 wire _25749_;
 wire _25750_;
 wire _25751_;
 wire _25752_;
 wire _25753_;
 wire _25754_;
 wire _25755_;
 wire _25756_;
 wire _25757_;
 wire _25758_;
 wire _25759_;
 wire _25760_;
 wire _25761_;
 wire _25762_;
 wire _25763_;
 wire _25764_;
 wire _25765_;
 wire _25766_;
 wire _25767_;
 wire _25768_;
 wire _25769_;
 wire _25770_;
 wire _25771_;
 wire _25772_;
 wire _25773_;
 wire _25774_;
 wire _25775_;
 wire _25776_;
 wire _25777_;
 wire _25778_;
 wire _25779_;
 wire _25780_;
 wire _25781_;
 wire _25782_;
 wire _25783_;
 wire _25784_;
 wire _25785_;
 wire _25786_;
 wire _25787_;
 wire _25788_;
 wire _25789_;
 wire _25790_;
 wire _25791_;
 wire _25792_;
 wire _25793_;
 wire _25794_;
 wire _25795_;
 wire _25796_;
 wire _25797_;
 wire _25798_;
 wire _25799_;
 wire _25800_;
 wire _25801_;
 wire _25802_;
 wire _25803_;
 wire _25804_;
 wire _25805_;
 wire _25806_;
 wire _25807_;
 wire _25808_;
 wire _25809_;
 wire _25810_;
 wire _25811_;
 wire _25812_;
 wire _25813_;
 wire _25814_;
 wire _25815_;
 wire _25816_;
 wire _25817_;
 wire _25818_;
 wire _25819_;
 wire _25820_;
 wire _25821_;
 wire _25822_;
 wire _25823_;
 wire _25824_;
 wire _25825_;
 wire _25826_;
 wire _25827_;
 wire _25828_;
 wire _25829_;
 wire _25830_;
 wire _25831_;
 wire _25832_;
 wire _25833_;
 wire _25834_;
 wire _25835_;
 wire _25836_;
 wire _25837_;
 wire _25838_;
 wire _25839_;
 wire _25840_;
 wire _25841_;
 wire _25842_;
 wire _25843_;
 wire _25844_;
 wire _25845_;
 wire _25846_;
 wire _25847_;
 wire _25848_;
 wire _25849_;
 wire _25850_;
 wire _25851_;
 wire _25852_;
 wire _25853_;
 wire _25854_;
 wire _25855_;
 wire _25856_;
 wire _25857_;
 wire _25858_;
 wire _25859_;
 wire _25860_;
 wire _25861_;
 wire _25862_;
 wire _25863_;
 wire _25864_;
 wire _25865_;
 wire _25866_;
 wire _25867_;
 wire _25868_;
 wire _25869_;
 wire _25870_;
 wire _25871_;
 wire _25872_;
 wire _25873_;
 wire _25874_;
 wire _25875_;
 wire _25876_;
 wire _25877_;
 wire _25878_;
 wire _25879_;
 wire _25880_;
 wire _25881_;
 wire _25882_;
 wire _25883_;
 wire _25884_;
 wire _25885_;
 wire _25886_;
 wire _25887_;
 wire _25888_;
 wire _25889_;
 wire _25890_;
 wire _25891_;
 wire _25892_;
 wire _25893_;
 wire _25894_;
 wire _25895_;
 wire _25896_;
 wire _25897_;
 wire _25898_;
 wire _25899_;
 wire _25900_;
 wire _25901_;
 wire _25902_;
 wire _25903_;
 wire _25904_;
 wire _25905_;
 wire _25906_;
 wire _25907_;
 wire _25908_;
 wire _25909_;
 wire _25910_;
 wire _25911_;
 wire _25912_;
 wire _25913_;
 wire _25914_;
 wire _25915_;
 wire _25916_;
 wire _25917_;
 wire _25918_;
 wire _25919_;
 wire _25920_;
 wire _25921_;
 wire _25922_;
 wire _25923_;
 wire _25924_;
 wire _25925_;
 wire _25926_;
 wire _25927_;
 wire _25928_;
 wire _25929_;
 wire _25930_;
 wire _25931_;
 wire _25932_;
 wire _25933_;
 wire _25934_;
 wire _25935_;
 wire _25936_;
 wire _25937_;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0_0_wb_clk_i;
 wire clknet_2_1_0_wb_clk_i;
 wire clknet_2_2_0_wb_clk_i;
 wire clknet_2_3_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_128_wb_clk_i;
 wire clknet_leaf_129_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_130_wb_clk_i;
 wire clknet_leaf_131_wb_clk_i;
 wire clknet_leaf_132_wb_clk_i;
 wire clknet_leaf_133_wb_clk_i;
 wire clknet_leaf_134_wb_clk_i;
 wire clknet_leaf_135_wb_clk_i;
 wire clknet_leaf_136_wb_clk_i;
 wire clknet_leaf_137_wb_clk_i;
 wire clknet_leaf_138_wb_clk_i;
 wire clknet_leaf_139_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_140_wb_clk_i;
 wire clknet_leaf_141_wb_clk_i;
 wire clknet_leaf_142_wb_clk_i;
 wire clknet_leaf_143_wb_clk_i;
 wire clknet_leaf_144_wb_clk_i;
 wire clknet_leaf_145_wb_clk_i;
 wire clknet_leaf_146_wb_clk_i;
 wire clknet_leaf_147_wb_clk_i;
 wire clknet_leaf_148_wb_clk_i;
 wire clknet_leaf_149_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_150_wb_clk_i;
 wire clknet_leaf_151_wb_clk_i;
 wire clknet_leaf_152_wb_clk_i;
 wire clknet_leaf_153_wb_clk_i;
 wire clknet_leaf_154_wb_clk_i;
 wire clknet_leaf_155_wb_clk_i;
 wire clknet_leaf_156_wb_clk_i;
 wire clknet_leaf_157_wb_clk_i;
 wire clknet_leaf_158_wb_clk_i;
 wire clknet_leaf_159_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_160_wb_clk_i;
 wire clknet_leaf_161_wb_clk_i;
 wire clknet_leaf_162_wb_clk_i;
 wire clknet_leaf_163_wb_clk_i;
 wire clknet_leaf_164_wb_clk_i;
 wire clknet_leaf_165_wb_clk_i;
 wire clknet_leaf_166_wb_clk_i;
 wire clknet_leaf_167_wb_clk_i;
 wire clknet_leaf_168_wb_clk_i;
 wire clknet_leaf_169_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_170_wb_clk_i;
 wire clknet_leaf_171_wb_clk_i;
 wire clknet_leaf_172_wb_clk_i;
 wire clknet_leaf_173_wb_clk_i;
 wire clknet_leaf_174_wb_clk_i;
 wire clknet_leaf_175_wb_clk_i;
 wire clknet_leaf_176_wb_clk_i;
 wire clknet_leaf_177_wb_clk_i;
 wire clknet_leaf_178_wb_clk_i;
 wire clknet_leaf_179_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_180_wb_clk_i;
 wire clknet_leaf_181_wb_clk_i;
 wire clknet_leaf_182_wb_clk_i;
 wire clknet_leaf_183_wb_clk_i;
 wire clknet_leaf_184_wb_clk_i;
 wire clknet_leaf_185_wb_clk_i;
 wire clknet_leaf_186_wb_clk_i;
 wire clknet_leaf_187_wb_clk_i;
 wire clknet_leaf_188_wb_clk_i;
 wire clknet_leaf_189_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_190_wb_clk_i;
 wire clknet_leaf_191_wb_clk_i;
 wire clknet_leaf_192_wb_clk_i;
 wire clknet_leaf_193_wb_clk_i;
 wire clknet_leaf_194_wb_clk_i;
 wire clknet_leaf_195_wb_clk_i;
 wire clknet_leaf_196_wb_clk_i;
 wire clknet_leaf_197_wb_clk_i;
 wire clknet_leaf_198_wb_clk_i;
 wire clknet_leaf_199_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_200_wb_clk_i;
 wire clknet_leaf_202_wb_clk_i;
 wire clknet_leaf_203_wb_clk_i;
 wire clknet_leaf_204_wb_clk_i;
 wire clknet_leaf_205_wb_clk_i;
 wire clknet_leaf_206_wb_clk_i;
 wire clknet_leaf_207_wb_clk_i;
 wire clknet_leaf_208_wb_clk_i;
 wire clknet_leaf_209_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_210_wb_clk_i;
 wire clknet_leaf_211_wb_clk_i;
 wire clknet_leaf_212_wb_clk_i;
 wire clknet_leaf_213_wb_clk_i;
 wire clknet_leaf_214_wb_clk_i;
 wire clknet_leaf_215_wb_clk_i;
 wire clknet_leaf_216_wb_clk_i;
 wire clknet_leaf_218_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_84_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net53;
 wire net54;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \tholin_riscv.Bimm[10] ;
 wire \tholin_riscv.Bimm[11] ;
 wire \tholin_riscv.Bimm[12] ;
 wire \tholin_riscv.Bimm[1] ;
 wire \tholin_riscv.Bimm[2] ;
 wire \tholin_riscv.Bimm[3] ;
 wire \tholin_riscv.Bimm[4] ;
 wire \tholin_riscv.Bimm[5] ;
 wire \tholin_riscv.Bimm[6] ;
 wire \tholin_riscv.Bimm[7] ;
 wire \tholin_riscv.Bimm[8] ;
 wire \tholin_riscv.Bimm[9] ;
 wire \tholin_riscv.Iimm[0] ;
 wire \tholin_riscv.Iimm[1] ;
 wire \tholin_riscv.Iimm[2] ;
 wire \tholin_riscv.Iimm[3] ;
 wire \tholin_riscv.Iimm[4] ;
 wire \tholin_riscv.Jimm[12] ;
 wire \tholin_riscv.Jimm[13] ;
 wire \tholin_riscv.Jimm[14] ;
 wire \tholin_riscv.Jimm[15] ;
 wire \tholin_riscv.Jimm[16] ;
 wire \tholin_riscv.Jimm[17] ;
 wire \tholin_riscv.Jimm[18] ;
 wire \tholin_riscv.Jimm[19] ;
 wire \tholin_riscv.PCE[0] ;
 wire \tholin_riscv.PCE[10] ;
 wire \tholin_riscv.PCE[11] ;
 wire \tholin_riscv.PCE[12] ;
 wire \tholin_riscv.PCE[13] ;
 wire \tholin_riscv.PCE[14] ;
 wire \tholin_riscv.PCE[15] ;
 wire \tholin_riscv.PCE[16] ;
 wire \tholin_riscv.PCE[17] ;
 wire \tholin_riscv.PCE[18] ;
 wire \tholin_riscv.PCE[19] ;
 wire \tholin_riscv.PCE[1] ;
 wire \tholin_riscv.PCE[20] ;
 wire \tholin_riscv.PCE[21] ;
 wire \tholin_riscv.PCE[22] ;
 wire \tholin_riscv.PCE[23] ;
 wire \tholin_riscv.PCE[24] ;
 wire \tholin_riscv.PCE[25] ;
 wire \tholin_riscv.PCE[26] ;
 wire \tholin_riscv.PCE[27] ;
 wire \tholin_riscv.PCE[28] ;
 wire \tholin_riscv.PCE[29] ;
 wire \tholin_riscv.PCE[2] ;
 wire \tholin_riscv.PCE[30] ;
 wire \tholin_riscv.PCE[31] ;
 wire \tholin_riscv.PCE[3] ;
 wire \tholin_riscv.PCE[4] ;
 wire \tholin_riscv.PCE[5] ;
 wire \tholin_riscv.PCE[6] ;
 wire \tholin_riscv.PCE[7] ;
 wire \tholin_riscv.PCE[8] ;
 wire \tholin_riscv.PCE[9] ;
 wire \tholin_riscv.PC[0] ;
 wire \tholin_riscv.PC[10] ;
 wire \tholin_riscv.PC[11] ;
 wire \tholin_riscv.PC[12] ;
 wire \tholin_riscv.PC[13] ;
 wire \tholin_riscv.PC[14] ;
 wire \tholin_riscv.PC[15] ;
 wire \tholin_riscv.PC[16] ;
 wire \tholin_riscv.PC[17] ;
 wire \tholin_riscv.PC[18] ;
 wire \tholin_riscv.PC[19] ;
 wire \tholin_riscv.PC[1] ;
 wire \tholin_riscv.PC[20] ;
 wire \tholin_riscv.PC[21] ;
 wire \tholin_riscv.PC[22] ;
 wire \tholin_riscv.PC[23] ;
 wire \tholin_riscv.PC[24] ;
 wire \tholin_riscv.PC[25] ;
 wire \tholin_riscv.PC[26] ;
 wire \tholin_riscv.PC[27] ;
 wire \tholin_riscv.PC[28] ;
 wire \tholin_riscv.PC[29] ;
 wire \tholin_riscv.PC[2] ;
 wire \tholin_riscv.PC[30] ;
 wire \tholin_riscv.PC[31] ;
 wire \tholin_riscv.PC[3] ;
 wire \tholin_riscv.PC[4] ;
 wire \tholin_riscv.PC[5] ;
 wire \tholin_riscv.PC[6] ;
 wire \tholin_riscv.PC[7] ;
 wire \tholin_riscv.PC[8] ;
 wire \tholin_riscv.PC[9] ;
 wire \tholin_riscv.PORT_dir[0] ;
 wire \tholin_riscv.PORT_dir[1] ;
 wire \tholin_riscv.PORT_dir[2] ;
 wire \tholin_riscv.PORT_dir[3] ;
 wire \tholin_riscv.PORT_dir[4] ;
 wire \tholin_riscv.PORT_dir[5] ;
 wire \tholin_riscv.current_irq[0] ;
 wire \tholin_riscv.current_irq[1] ;
 wire \tholin_riscv.cycle[0] ;
 wire \tholin_riscv.cycle[1] ;
 wire \tholin_riscv.cycle[2] ;
 wire \tholin_riscv.cycle[3] ;
 wire \tholin_riscv.div_counter[0] ;
 wire \tholin_riscv.div_counter[1] ;
 wire \tholin_riscv.div_counter[2] ;
 wire \tholin_riscv.div_counter[3] ;
 wire \tholin_riscv.div_counter[4] ;
 wire \tholin_riscv.div_res[0] ;
 wire \tholin_riscv.div_res[10] ;
 wire \tholin_riscv.div_res[11] ;
 wire \tholin_riscv.div_res[12] ;
 wire \tholin_riscv.div_res[13] ;
 wire \tholin_riscv.div_res[14] ;
 wire \tholin_riscv.div_res[15] ;
 wire \tholin_riscv.div_res[16] ;
 wire \tholin_riscv.div_res[17] ;
 wire \tholin_riscv.div_res[18] ;
 wire \tholin_riscv.div_res[19] ;
 wire \tholin_riscv.div_res[1] ;
 wire \tholin_riscv.div_res[20] ;
 wire \tholin_riscv.div_res[21] ;
 wire \tholin_riscv.div_res[22] ;
 wire \tholin_riscv.div_res[23] ;
 wire \tholin_riscv.div_res[24] ;
 wire \tholin_riscv.div_res[25] ;
 wire \tholin_riscv.div_res[26] ;
 wire \tholin_riscv.div_res[27] ;
 wire \tholin_riscv.div_res[28] ;
 wire \tholin_riscv.div_res[29] ;
 wire \tholin_riscv.div_res[2] ;
 wire \tholin_riscv.div_res[30] ;
 wire \tholin_riscv.div_res[31] ;
 wire \tholin_riscv.div_res[3] ;
 wire \tholin_riscv.div_res[4] ;
 wire \tholin_riscv.div_res[5] ;
 wire \tholin_riscv.div_res[6] ;
 wire \tholin_riscv.div_res[7] ;
 wire \tholin_riscv.div_res[8] ;
 wire \tholin_riscv.div_res[9] ;
 wire \tholin_riscv.div_shifter[0] ;
 wire \tholin_riscv.div_shifter[10] ;
 wire \tholin_riscv.div_shifter[11] ;
 wire \tholin_riscv.div_shifter[12] ;
 wire \tholin_riscv.div_shifter[13] ;
 wire \tholin_riscv.div_shifter[14] ;
 wire \tholin_riscv.div_shifter[15] ;
 wire \tholin_riscv.div_shifter[16] ;
 wire \tholin_riscv.div_shifter[17] ;
 wire \tholin_riscv.div_shifter[18] ;
 wire \tholin_riscv.div_shifter[19] ;
 wire \tholin_riscv.div_shifter[1] ;
 wire \tholin_riscv.div_shifter[20] ;
 wire \tholin_riscv.div_shifter[21] ;
 wire \tholin_riscv.div_shifter[22] ;
 wire \tholin_riscv.div_shifter[23] ;
 wire \tholin_riscv.div_shifter[24] ;
 wire \tholin_riscv.div_shifter[25] ;
 wire \tholin_riscv.div_shifter[26] ;
 wire \tholin_riscv.div_shifter[27] ;
 wire \tholin_riscv.div_shifter[28] ;
 wire \tholin_riscv.div_shifter[29] ;
 wire \tholin_riscv.div_shifter[2] ;
 wire \tholin_riscv.div_shifter[30] ;
 wire \tholin_riscv.div_shifter[31] ;
 wire \tholin_riscv.div_shifter[32] ;
 wire \tholin_riscv.div_shifter[33] ;
 wire \tholin_riscv.div_shifter[34] ;
 wire \tholin_riscv.div_shifter[35] ;
 wire \tholin_riscv.div_shifter[36] ;
 wire \tholin_riscv.div_shifter[37] ;
 wire \tholin_riscv.div_shifter[38] ;
 wire \tholin_riscv.div_shifter[39] ;
 wire \tholin_riscv.div_shifter[3] ;
 wire \tholin_riscv.div_shifter[40] ;
 wire \tholin_riscv.div_shifter[41] ;
 wire \tholin_riscv.div_shifter[42] ;
 wire \tholin_riscv.div_shifter[43] ;
 wire \tholin_riscv.div_shifter[44] ;
 wire \tholin_riscv.div_shifter[45] ;
 wire \tholin_riscv.div_shifter[46] ;
 wire \tholin_riscv.div_shifter[47] ;
 wire \tholin_riscv.div_shifter[48] ;
 wire \tholin_riscv.div_shifter[49] ;
 wire \tholin_riscv.div_shifter[4] ;
 wire \tholin_riscv.div_shifter[50] ;
 wire \tholin_riscv.div_shifter[51] ;
 wire \tholin_riscv.div_shifter[52] ;
 wire \tholin_riscv.div_shifter[53] ;
 wire \tholin_riscv.div_shifter[54] ;
 wire \tholin_riscv.div_shifter[55] ;
 wire \tholin_riscv.div_shifter[56] ;
 wire \tholin_riscv.div_shifter[57] ;
 wire \tholin_riscv.div_shifter[58] ;
 wire \tholin_riscv.div_shifter[59] ;
 wire \tholin_riscv.div_shifter[5] ;
 wire \tholin_riscv.div_shifter[60] ;
 wire \tholin_riscv.div_shifter[61] ;
 wire \tholin_riscv.div_shifter[62] ;
 wire \tholin_riscv.div_shifter[63] ;
 wire \tholin_riscv.div_shifter[6] ;
 wire \tholin_riscv.div_shifter[7] ;
 wire \tholin_riscv.div_shifter[8] ;
 wire \tholin_riscv.div_shifter[9] ;
 wire \tholin_riscv.instr[0] ;
 wire \tholin_riscv.instr[1] ;
 wire \tholin_riscv.instr[2] ;
 wire \tholin_riscv.instr[3] ;
 wire \tholin_riscv.instr[4] ;
 wire \tholin_riscv.instr[5] ;
 wire \tholin_riscv.instr[6] ;
 wire \tholin_riscv.int_enabled ;
 wire \tholin_riscv.intr_vec[0] ;
 wire \tholin_riscv.intr_vec[10] ;
 wire \tholin_riscv.intr_vec[11] ;
 wire \tholin_riscv.intr_vec[12] ;
 wire \tholin_riscv.intr_vec[13] ;
 wire \tholin_riscv.intr_vec[14] ;
 wire \tholin_riscv.intr_vec[15] ;
 wire \tholin_riscv.intr_vec[16] ;
 wire \tholin_riscv.intr_vec[17] ;
 wire \tholin_riscv.intr_vec[18] ;
 wire \tholin_riscv.intr_vec[19] ;
 wire \tholin_riscv.intr_vec[1] ;
 wire \tholin_riscv.intr_vec[20] ;
 wire \tholin_riscv.intr_vec[21] ;
 wire \tholin_riscv.intr_vec[22] ;
 wire \tholin_riscv.intr_vec[23] ;
 wire \tholin_riscv.intr_vec[24] ;
 wire \tholin_riscv.intr_vec[25] ;
 wire \tholin_riscv.intr_vec[26] ;
 wire \tholin_riscv.intr_vec[27] ;
 wire \tholin_riscv.intr_vec[28] ;
 wire \tholin_riscv.intr_vec[29] ;
 wire \tholin_riscv.intr_vec[2] ;
 wire \tholin_riscv.intr_vec[3] ;
 wire \tholin_riscv.intr_vec[4] ;
 wire \tholin_riscv.intr_vec[5] ;
 wire \tholin_riscv.intr_vec[6] ;
 wire \tholin_riscv.intr_vec[7] ;
 wire \tholin_riscv.intr_vec[8] ;
 wire \tholin_riscv.intr_vec[9] ;
 wire \tholin_riscv.io_int_enable ;
 wire \tholin_riscv.io_size[0] ;
 wire \tholin_riscv.io_size[1] ;
 wire \tholin_riscv.irqs[0] ;
 wire \tholin_riscv.irqs[1] ;
 wire \tholin_riscv.irqs[2] ;
 wire \tholin_riscv.is_write ;
 wire \tholin_riscv.last_io_state ;
 wire \tholin_riscv.load_dest[0] ;
 wire \tholin_riscv.load_dest[1] ;
 wire \tholin_riscv.load_dest[2] ;
 wire \tholin_riscv.load_dest[3] ;
 wire \tholin_riscv.load_dest[4] ;
 wire \tholin_riscv.load_funct ;
 wire \tholin_riscv.mul_delay ;
 wire \tholin_riscv.regs[0][0] ;
 wire \tholin_riscv.regs[0][10] ;
 wire \tholin_riscv.regs[0][11] ;
 wire \tholin_riscv.regs[0][12] ;
 wire \tholin_riscv.regs[0][13] ;
 wire \tholin_riscv.regs[0][14] ;
 wire \tholin_riscv.regs[0][15] ;
 wire \tholin_riscv.regs[0][16] ;
 wire \tholin_riscv.regs[0][17] ;
 wire \tholin_riscv.regs[0][18] ;
 wire \tholin_riscv.regs[0][19] ;
 wire \tholin_riscv.regs[0][1] ;
 wire \tholin_riscv.regs[0][20] ;
 wire \tholin_riscv.regs[0][21] ;
 wire \tholin_riscv.regs[0][22] ;
 wire \tholin_riscv.regs[0][23] ;
 wire \tholin_riscv.regs[0][24] ;
 wire \tholin_riscv.regs[0][25] ;
 wire \tholin_riscv.regs[0][26] ;
 wire \tholin_riscv.regs[0][27] ;
 wire \tholin_riscv.regs[0][28] ;
 wire \tholin_riscv.regs[0][29] ;
 wire \tholin_riscv.regs[0][2] ;
 wire \tholin_riscv.regs[0][30] ;
 wire \tholin_riscv.regs[0][31] ;
 wire \tholin_riscv.regs[0][3] ;
 wire \tholin_riscv.regs[0][4] ;
 wire \tholin_riscv.regs[0][5] ;
 wire \tholin_riscv.regs[0][6] ;
 wire \tholin_riscv.regs[0][7] ;
 wire \tholin_riscv.regs[0][8] ;
 wire \tholin_riscv.regs[0][9] ;
 wire \tholin_riscv.regs[10][0] ;
 wire \tholin_riscv.regs[10][10] ;
 wire \tholin_riscv.regs[10][11] ;
 wire \tholin_riscv.regs[10][12] ;
 wire \tholin_riscv.regs[10][13] ;
 wire \tholin_riscv.regs[10][14] ;
 wire \tholin_riscv.regs[10][15] ;
 wire \tholin_riscv.regs[10][16] ;
 wire \tholin_riscv.regs[10][17] ;
 wire \tholin_riscv.regs[10][18] ;
 wire \tholin_riscv.regs[10][19] ;
 wire \tholin_riscv.regs[10][1] ;
 wire \tholin_riscv.regs[10][20] ;
 wire \tholin_riscv.regs[10][21] ;
 wire \tholin_riscv.regs[10][22] ;
 wire \tholin_riscv.regs[10][23] ;
 wire \tholin_riscv.regs[10][24] ;
 wire \tholin_riscv.regs[10][25] ;
 wire \tholin_riscv.regs[10][26] ;
 wire \tholin_riscv.regs[10][27] ;
 wire \tholin_riscv.regs[10][28] ;
 wire \tholin_riscv.regs[10][29] ;
 wire \tholin_riscv.regs[10][2] ;
 wire \tholin_riscv.regs[10][30] ;
 wire \tholin_riscv.regs[10][31] ;
 wire \tholin_riscv.regs[10][3] ;
 wire \tholin_riscv.regs[10][4] ;
 wire \tholin_riscv.regs[10][5] ;
 wire \tholin_riscv.regs[10][6] ;
 wire \tholin_riscv.regs[10][7] ;
 wire \tholin_riscv.regs[10][8] ;
 wire \tholin_riscv.regs[10][9] ;
 wire \tholin_riscv.regs[11][0] ;
 wire \tholin_riscv.regs[11][10] ;
 wire \tholin_riscv.regs[11][11] ;
 wire \tholin_riscv.regs[11][12] ;
 wire \tholin_riscv.regs[11][13] ;
 wire \tholin_riscv.regs[11][14] ;
 wire \tholin_riscv.regs[11][15] ;
 wire \tholin_riscv.regs[11][16] ;
 wire \tholin_riscv.regs[11][17] ;
 wire \tholin_riscv.regs[11][18] ;
 wire \tholin_riscv.regs[11][19] ;
 wire \tholin_riscv.regs[11][1] ;
 wire \tholin_riscv.regs[11][20] ;
 wire \tholin_riscv.regs[11][21] ;
 wire \tholin_riscv.regs[11][22] ;
 wire \tholin_riscv.regs[11][23] ;
 wire \tholin_riscv.regs[11][24] ;
 wire \tholin_riscv.regs[11][25] ;
 wire \tholin_riscv.regs[11][26] ;
 wire \tholin_riscv.regs[11][27] ;
 wire \tholin_riscv.regs[11][28] ;
 wire \tholin_riscv.regs[11][29] ;
 wire \tholin_riscv.regs[11][2] ;
 wire \tholin_riscv.regs[11][30] ;
 wire \tholin_riscv.regs[11][31] ;
 wire \tholin_riscv.regs[11][3] ;
 wire \tholin_riscv.regs[11][4] ;
 wire \tholin_riscv.regs[11][5] ;
 wire \tholin_riscv.regs[11][6] ;
 wire \tholin_riscv.regs[11][7] ;
 wire \tholin_riscv.regs[11][8] ;
 wire \tholin_riscv.regs[11][9] ;
 wire \tholin_riscv.regs[12][0] ;
 wire \tholin_riscv.regs[12][10] ;
 wire \tholin_riscv.regs[12][11] ;
 wire \tholin_riscv.regs[12][12] ;
 wire \tholin_riscv.regs[12][13] ;
 wire \tholin_riscv.regs[12][14] ;
 wire \tholin_riscv.regs[12][15] ;
 wire \tholin_riscv.regs[12][16] ;
 wire \tholin_riscv.regs[12][17] ;
 wire \tholin_riscv.regs[12][18] ;
 wire \tholin_riscv.regs[12][19] ;
 wire \tholin_riscv.regs[12][1] ;
 wire \tholin_riscv.regs[12][20] ;
 wire \tholin_riscv.regs[12][21] ;
 wire \tholin_riscv.regs[12][22] ;
 wire \tholin_riscv.regs[12][23] ;
 wire \tholin_riscv.regs[12][24] ;
 wire \tholin_riscv.regs[12][25] ;
 wire \tholin_riscv.regs[12][26] ;
 wire \tholin_riscv.regs[12][27] ;
 wire \tholin_riscv.regs[12][28] ;
 wire \tholin_riscv.regs[12][29] ;
 wire \tholin_riscv.regs[12][2] ;
 wire \tholin_riscv.regs[12][30] ;
 wire \tholin_riscv.regs[12][31] ;
 wire \tholin_riscv.regs[12][3] ;
 wire \tholin_riscv.regs[12][4] ;
 wire \tholin_riscv.regs[12][5] ;
 wire \tholin_riscv.regs[12][6] ;
 wire \tholin_riscv.regs[12][7] ;
 wire \tholin_riscv.regs[12][8] ;
 wire \tholin_riscv.regs[12][9] ;
 wire \tholin_riscv.regs[13][0] ;
 wire \tholin_riscv.regs[13][10] ;
 wire \tholin_riscv.regs[13][11] ;
 wire \tholin_riscv.regs[13][12] ;
 wire \tholin_riscv.regs[13][13] ;
 wire \tholin_riscv.regs[13][14] ;
 wire \tholin_riscv.regs[13][15] ;
 wire \tholin_riscv.regs[13][16] ;
 wire \tholin_riscv.regs[13][17] ;
 wire \tholin_riscv.regs[13][18] ;
 wire \tholin_riscv.regs[13][19] ;
 wire \tholin_riscv.regs[13][1] ;
 wire \tholin_riscv.regs[13][20] ;
 wire \tholin_riscv.regs[13][21] ;
 wire \tholin_riscv.regs[13][22] ;
 wire \tholin_riscv.regs[13][23] ;
 wire \tholin_riscv.regs[13][24] ;
 wire \tholin_riscv.regs[13][25] ;
 wire \tholin_riscv.regs[13][26] ;
 wire \tholin_riscv.regs[13][27] ;
 wire \tholin_riscv.regs[13][28] ;
 wire \tholin_riscv.regs[13][29] ;
 wire \tholin_riscv.regs[13][2] ;
 wire \tholin_riscv.regs[13][30] ;
 wire \tholin_riscv.regs[13][31] ;
 wire \tholin_riscv.regs[13][3] ;
 wire \tholin_riscv.regs[13][4] ;
 wire \tholin_riscv.regs[13][5] ;
 wire \tholin_riscv.regs[13][6] ;
 wire \tholin_riscv.regs[13][7] ;
 wire \tholin_riscv.regs[13][8] ;
 wire \tholin_riscv.regs[13][9] ;
 wire \tholin_riscv.regs[14][0] ;
 wire \tholin_riscv.regs[14][10] ;
 wire \tholin_riscv.regs[14][11] ;
 wire \tholin_riscv.regs[14][12] ;
 wire \tholin_riscv.regs[14][13] ;
 wire \tholin_riscv.regs[14][14] ;
 wire \tholin_riscv.regs[14][15] ;
 wire \tholin_riscv.regs[14][16] ;
 wire \tholin_riscv.regs[14][17] ;
 wire \tholin_riscv.regs[14][18] ;
 wire \tholin_riscv.regs[14][19] ;
 wire \tholin_riscv.regs[14][1] ;
 wire \tholin_riscv.regs[14][20] ;
 wire \tholin_riscv.regs[14][21] ;
 wire \tholin_riscv.regs[14][22] ;
 wire \tholin_riscv.regs[14][23] ;
 wire \tholin_riscv.regs[14][24] ;
 wire \tholin_riscv.regs[14][25] ;
 wire \tholin_riscv.regs[14][26] ;
 wire \tholin_riscv.regs[14][27] ;
 wire \tholin_riscv.regs[14][28] ;
 wire \tholin_riscv.regs[14][29] ;
 wire \tholin_riscv.regs[14][2] ;
 wire \tholin_riscv.regs[14][30] ;
 wire \tholin_riscv.regs[14][31] ;
 wire \tholin_riscv.regs[14][3] ;
 wire \tholin_riscv.regs[14][4] ;
 wire \tholin_riscv.regs[14][5] ;
 wire \tholin_riscv.regs[14][6] ;
 wire \tholin_riscv.regs[14][7] ;
 wire \tholin_riscv.regs[14][8] ;
 wire \tholin_riscv.regs[14][9] ;
 wire \tholin_riscv.regs[15][0] ;
 wire \tholin_riscv.regs[15][10] ;
 wire \tholin_riscv.regs[15][11] ;
 wire \tholin_riscv.regs[15][12] ;
 wire \tholin_riscv.regs[15][13] ;
 wire \tholin_riscv.regs[15][14] ;
 wire \tholin_riscv.regs[15][15] ;
 wire \tholin_riscv.regs[15][16] ;
 wire \tholin_riscv.regs[15][17] ;
 wire \tholin_riscv.regs[15][18] ;
 wire \tholin_riscv.regs[15][19] ;
 wire \tholin_riscv.regs[15][1] ;
 wire \tholin_riscv.regs[15][20] ;
 wire \tholin_riscv.regs[15][21] ;
 wire \tholin_riscv.regs[15][22] ;
 wire \tholin_riscv.regs[15][23] ;
 wire \tholin_riscv.regs[15][24] ;
 wire \tholin_riscv.regs[15][25] ;
 wire \tholin_riscv.regs[15][26] ;
 wire \tholin_riscv.regs[15][27] ;
 wire \tholin_riscv.regs[15][28] ;
 wire \tholin_riscv.regs[15][29] ;
 wire \tholin_riscv.regs[15][2] ;
 wire \tholin_riscv.regs[15][30] ;
 wire \tholin_riscv.regs[15][31] ;
 wire \tholin_riscv.regs[15][3] ;
 wire \tholin_riscv.regs[15][4] ;
 wire \tholin_riscv.regs[15][5] ;
 wire \tholin_riscv.regs[15][6] ;
 wire \tholin_riscv.regs[15][7] ;
 wire \tholin_riscv.regs[15][8] ;
 wire \tholin_riscv.regs[15][9] ;
 wire \tholin_riscv.regs[16][0] ;
 wire \tholin_riscv.regs[16][10] ;
 wire \tholin_riscv.regs[16][11] ;
 wire \tholin_riscv.regs[16][12] ;
 wire \tholin_riscv.regs[16][13] ;
 wire \tholin_riscv.regs[16][14] ;
 wire \tholin_riscv.regs[16][15] ;
 wire \tholin_riscv.regs[16][16] ;
 wire \tholin_riscv.regs[16][17] ;
 wire \tholin_riscv.regs[16][18] ;
 wire \tholin_riscv.regs[16][19] ;
 wire \tholin_riscv.regs[16][1] ;
 wire \tholin_riscv.regs[16][20] ;
 wire \tholin_riscv.regs[16][21] ;
 wire \tholin_riscv.regs[16][22] ;
 wire \tholin_riscv.regs[16][23] ;
 wire \tholin_riscv.regs[16][24] ;
 wire \tholin_riscv.regs[16][25] ;
 wire \tholin_riscv.regs[16][26] ;
 wire \tholin_riscv.regs[16][27] ;
 wire \tholin_riscv.regs[16][28] ;
 wire \tholin_riscv.regs[16][29] ;
 wire \tholin_riscv.regs[16][2] ;
 wire \tholin_riscv.regs[16][30] ;
 wire \tholin_riscv.regs[16][31] ;
 wire \tholin_riscv.regs[16][3] ;
 wire \tholin_riscv.regs[16][4] ;
 wire \tholin_riscv.regs[16][5] ;
 wire \tholin_riscv.regs[16][6] ;
 wire \tholin_riscv.regs[16][7] ;
 wire \tholin_riscv.regs[16][8] ;
 wire \tholin_riscv.regs[16][9] ;
 wire \tholin_riscv.regs[17][0] ;
 wire \tholin_riscv.regs[17][10] ;
 wire \tholin_riscv.regs[17][11] ;
 wire \tholin_riscv.regs[17][12] ;
 wire \tholin_riscv.regs[17][13] ;
 wire \tholin_riscv.regs[17][14] ;
 wire \tholin_riscv.regs[17][15] ;
 wire \tholin_riscv.regs[17][16] ;
 wire \tholin_riscv.regs[17][17] ;
 wire \tholin_riscv.regs[17][18] ;
 wire \tholin_riscv.regs[17][19] ;
 wire \tholin_riscv.regs[17][1] ;
 wire \tholin_riscv.regs[17][20] ;
 wire \tholin_riscv.regs[17][21] ;
 wire \tholin_riscv.regs[17][22] ;
 wire \tholin_riscv.regs[17][23] ;
 wire \tholin_riscv.regs[17][24] ;
 wire \tholin_riscv.regs[17][25] ;
 wire \tholin_riscv.regs[17][26] ;
 wire \tholin_riscv.regs[17][27] ;
 wire \tholin_riscv.regs[17][28] ;
 wire \tholin_riscv.regs[17][29] ;
 wire \tholin_riscv.regs[17][2] ;
 wire \tholin_riscv.regs[17][30] ;
 wire \tholin_riscv.regs[17][31] ;
 wire \tholin_riscv.regs[17][3] ;
 wire \tholin_riscv.regs[17][4] ;
 wire \tholin_riscv.regs[17][5] ;
 wire \tholin_riscv.regs[17][6] ;
 wire \tholin_riscv.regs[17][7] ;
 wire \tholin_riscv.regs[17][8] ;
 wire \tholin_riscv.regs[17][9] ;
 wire \tholin_riscv.regs[18][0] ;
 wire \tholin_riscv.regs[18][10] ;
 wire \tholin_riscv.regs[18][11] ;
 wire \tholin_riscv.regs[18][12] ;
 wire \tholin_riscv.regs[18][13] ;
 wire \tholin_riscv.regs[18][14] ;
 wire \tholin_riscv.regs[18][15] ;
 wire \tholin_riscv.regs[18][16] ;
 wire \tholin_riscv.regs[18][17] ;
 wire \tholin_riscv.regs[18][18] ;
 wire \tholin_riscv.regs[18][19] ;
 wire \tholin_riscv.regs[18][1] ;
 wire \tholin_riscv.regs[18][20] ;
 wire \tholin_riscv.regs[18][21] ;
 wire \tholin_riscv.regs[18][22] ;
 wire \tholin_riscv.regs[18][23] ;
 wire \tholin_riscv.regs[18][24] ;
 wire \tholin_riscv.regs[18][25] ;
 wire \tholin_riscv.regs[18][26] ;
 wire \tholin_riscv.regs[18][27] ;
 wire \tholin_riscv.regs[18][28] ;
 wire \tholin_riscv.regs[18][29] ;
 wire \tholin_riscv.regs[18][2] ;
 wire \tholin_riscv.regs[18][30] ;
 wire \tholin_riscv.regs[18][31] ;
 wire \tholin_riscv.regs[18][3] ;
 wire \tholin_riscv.regs[18][4] ;
 wire \tholin_riscv.regs[18][5] ;
 wire \tholin_riscv.regs[18][6] ;
 wire \tholin_riscv.regs[18][7] ;
 wire \tholin_riscv.regs[18][8] ;
 wire \tholin_riscv.regs[18][9] ;
 wire \tholin_riscv.regs[19][0] ;
 wire \tholin_riscv.regs[19][10] ;
 wire \tholin_riscv.regs[19][11] ;
 wire \tholin_riscv.regs[19][12] ;
 wire \tholin_riscv.regs[19][13] ;
 wire \tholin_riscv.regs[19][14] ;
 wire \tholin_riscv.regs[19][15] ;
 wire \tholin_riscv.regs[19][16] ;
 wire \tholin_riscv.regs[19][17] ;
 wire \tholin_riscv.regs[19][18] ;
 wire \tholin_riscv.regs[19][19] ;
 wire \tholin_riscv.regs[19][1] ;
 wire \tholin_riscv.regs[19][20] ;
 wire \tholin_riscv.regs[19][21] ;
 wire \tholin_riscv.regs[19][22] ;
 wire \tholin_riscv.regs[19][23] ;
 wire \tholin_riscv.regs[19][24] ;
 wire \tholin_riscv.regs[19][25] ;
 wire \tholin_riscv.regs[19][26] ;
 wire \tholin_riscv.regs[19][27] ;
 wire \tholin_riscv.regs[19][28] ;
 wire \tholin_riscv.regs[19][29] ;
 wire \tholin_riscv.regs[19][2] ;
 wire \tholin_riscv.regs[19][30] ;
 wire \tholin_riscv.regs[19][31] ;
 wire \tholin_riscv.regs[19][3] ;
 wire \tholin_riscv.regs[19][4] ;
 wire \tholin_riscv.regs[19][5] ;
 wire \tholin_riscv.regs[19][6] ;
 wire \tholin_riscv.regs[19][7] ;
 wire \tholin_riscv.regs[19][8] ;
 wire \tholin_riscv.regs[19][9] ;
 wire \tholin_riscv.regs[1][0] ;
 wire \tholin_riscv.regs[1][10] ;
 wire \tholin_riscv.regs[1][11] ;
 wire \tholin_riscv.regs[1][12] ;
 wire \tholin_riscv.regs[1][13] ;
 wire \tholin_riscv.regs[1][14] ;
 wire \tholin_riscv.regs[1][15] ;
 wire \tholin_riscv.regs[1][16] ;
 wire \tholin_riscv.regs[1][17] ;
 wire \tholin_riscv.regs[1][18] ;
 wire \tholin_riscv.regs[1][19] ;
 wire \tholin_riscv.regs[1][1] ;
 wire \tholin_riscv.regs[1][20] ;
 wire \tholin_riscv.regs[1][21] ;
 wire \tholin_riscv.regs[1][22] ;
 wire \tholin_riscv.regs[1][23] ;
 wire \tholin_riscv.regs[1][24] ;
 wire \tholin_riscv.regs[1][25] ;
 wire \tholin_riscv.regs[1][26] ;
 wire \tholin_riscv.regs[1][27] ;
 wire \tholin_riscv.regs[1][28] ;
 wire \tholin_riscv.regs[1][29] ;
 wire \tholin_riscv.regs[1][2] ;
 wire \tholin_riscv.regs[1][30] ;
 wire \tholin_riscv.regs[1][31] ;
 wire \tholin_riscv.regs[1][3] ;
 wire \tholin_riscv.regs[1][4] ;
 wire \tholin_riscv.regs[1][5] ;
 wire \tholin_riscv.regs[1][6] ;
 wire \tholin_riscv.regs[1][7] ;
 wire \tholin_riscv.regs[1][8] ;
 wire \tholin_riscv.regs[1][9] ;
 wire \tholin_riscv.regs[20][0] ;
 wire \tholin_riscv.regs[20][10] ;
 wire \tholin_riscv.regs[20][11] ;
 wire \tholin_riscv.regs[20][12] ;
 wire \tholin_riscv.regs[20][13] ;
 wire \tholin_riscv.regs[20][14] ;
 wire \tholin_riscv.regs[20][15] ;
 wire \tholin_riscv.regs[20][16] ;
 wire \tholin_riscv.regs[20][17] ;
 wire \tholin_riscv.regs[20][18] ;
 wire \tholin_riscv.regs[20][19] ;
 wire \tholin_riscv.regs[20][1] ;
 wire \tholin_riscv.regs[20][20] ;
 wire \tholin_riscv.regs[20][21] ;
 wire \tholin_riscv.regs[20][22] ;
 wire \tholin_riscv.regs[20][23] ;
 wire \tholin_riscv.regs[20][24] ;
 wire \tholin_riscv.regs[20][25] ;
 wire \tholin_riscv.regs[20][26] ;
 wire \tholin_riscv.regs[20][27] ;
 wire \tholin_riscv.regs[20][28] ;
 wire \tholin_riscv.regs[20][29] ;
 wire \tholin_riscv.regs[20][2] ;
 wire \tholin_riscv.regs[20][30] ;
 wire \tholin_riscv.regs[20][31] ;
 wire \tholin_riscv.regs[20][3] ;
 wire \tholin_riscv.regs[20][4] ;
 wire \tholin_riscv.regs[20][5] ;
 wire \tholin_riscv.regs[20][6] ;
 wire \tholin_riscv.regs[20][7] ;
 wire \tholin_riscv.regs[20][8] ;
 wire \tholin_riscv.regs[20][9] ;
 wire \tholin_riscv.regs[21][0] ;
 wire \tholin_riscv.regs[21][10] ;
 wire \tholin_riscv.regs[21][11] ;
 wire \tholin_riscv.regs[21][12] ;
 wire \tholin_riscv.regs[21][13] ;
 wire \tholin_riscv.regs[21][14] ;
 wire \tholin_riscv.regs[21][15] ;
 wire \tholin_riscv.regs[21][16] ;
 wire \tholin_riscv.regs[21][17] ;
 wire \tholin_riscv.regs[21][18] ;
 wire \tholin_riscv.regs[21][19] ;
 wire \tholin_riscv.regs[21][1] ;
 wire \tholin_riscv.regs[21][20] ;
 wire \tholin_riscv.regs[21][21] ;
 wire \tholin_riscv.regs[21][22] ;
 wire \tholin_riscv.regs[21][23] ;
 wire \tholin_riscv.regs[21][24] ;
 wire \tholin_riscv.regs[21][25] ;
 wire \tholin_riscv.regs[21][26] ;
 wire \tholin_riscv.regs[21][27] ;
 wire \tholin_riscv.regs[21][28] ;
 wire \tholin_riscv.regs[21][29] ;
 wire \tholin_riscv.regs[21][2] ;
 wire \tholin_riscv.regs[21][30] ;
 wire \tholin_riscv.regs[21][31] ;
 wire \tholin_riscv.regs[21][3] ;
 wire \tholin_riscv.regs[21][4] ;
 wire \tholin_riscv.regs[21][5] ;
 wire \tholin_riscv.regs[21][6] ;
 wire \tholin_riscv.regs[21][7] ;
 wire \tholin_riscv.regs[21][8] ;
 wire \tholin_riscv.regs[21][9] ;
 wire \tholin_riscv.regs[22][0] ;
 wire \tholin_riscv.regs[22][10] ;
 wire \tholin_riscv.regs[22][11] ;
 wire \tholin_riscv.regs[22][12] ;
 wire \tholin_riscv.regs[22][13] ;
 wire \tholin_riscv.regs[22][14] ;
 wire \tholin_riscv.regs[22][15] ;
 wire \tholin_riscv.regs[22][16] ;
 wire \tholin_riscv.regs[22][17] ;
 wire \tholin_riscv.regs[22][18] ;
 wire \tholin_riscv.regs[22][19] ;
 wire \tholin_riscv.regs[22][1] ;
 wire \tholin_riscv.regs[22][20] ;
 wire \tholin_riscv.regs[22][21] ;
 wire \tholin_riscv.regs[22][22] ;
 wire \tholin_riscv.regs[22][23] ;
 wire \tholin_riscv.regs[22][24] ;
 wire \tholin_riscv.regs[22][25] ;
 wire \tholin_riscv.regs[22][26] ;
 wire \tholin_riscv.regs[22][27] ;
 wire \tholin_riscv.regs[22][28] ;
 wire \tholin_riscv.regs[22][29] ;
 wire \tholin_riscv.regs[22][2] ;
 wire \tholin_riscv.regs[22][30] ;
 wire \tholin_riscv.regs[22][31] ;
 wire \tholin_riscv.regs[22][3] ;
 wire \tholin_riscv.regs[22][4] ;
 wire \tholin_riscv.regs[22][5] ;
 wire \tholin_riscv.regs[22][6] ;
 wire \tholin_riscv.regs[22][7] ;
 wire \tholin_riscv.regs[22][8] ;
 wire \tholin_riscv.regs[22][9] ;
 wire \tholin_riscv.regs[23][0] ;
 wire \tholin_riscv.regs[23][10] ;
 wire \tholin_riscv.regs[23][11] ;
 wire \tholin_riscv.regs[23][12] ;
 wire \tholin_riscv.regs[23][13] ;
 wire \tholin_riscv.regs[23][14] ;
 wire \tholin_riscv.regs[23][15] ;
 wire \tholin_riscv.regs[23][16] ;
 wire \tholin_riscv.regs[23][17] ;
 wire \tholin_riscv.regs[23][18] ;
 wire \tholin_riscv.regs[23][19] ;
 wire \tholin_riscv.regs[23][1] ;
 wire \tholin_riscv.regs[23][20] ;
 wire \tholin_riscv.regs[23][21] ;
 wire \tholin_riscv.regs[23][22] ;
 wire \tholin_riscv.regs[23][23] ;
 wire \tholin_riscv.regs[23][24] ;
 wire \tholin_riscv.regs[23][25] ;
 wire \tholin_riscv.regs[23][26] ;
 wire \tholin_riscv.regs[23][27] ;
 wire \tholin_riscv.regs[23][28] ;
 wire \tholin_riscv.regs[23][29] ;
 wire \tholin_riscv.regs[23][2] ;
 wire \tholin_riscv.regs[23][30] ;
 wire \tholin_riscv.regs[23][31] ;
 wire \tholin_riscv.regs[23][3] ;
 wire \tholin_riscv.regs[23][4] ;
 wire \tholin_riscv.regs[23][5] ;
 wire \tholin_riscv.regs[23][6] ;
 wire \tholin_riscv.regs[23][7] ;
 wire \tholin_riscv.regs[23][8] ;
 wire \tholin_riscv.regs[23][9] ;
 wire \tholin_riscv.regs[24][0] ;
 wire \tholin_riscv.regs[24][10] ;
 wire \tholin_riscv.regs[24][11] ;
 wire \tholin_riscv.regs[24][12] ;
 wire \tholin_riscv.regs[24][13] ;
 wire \tholin_riscv.regs[24][14] ;
 wire \tholin_riscv.regs[24][15] ;
 wire \tholin_riscv.regs[24][16] ;
 wire \tholin_riscv.regs[24][17] ;
 wire \tholin_riscv.regs[24][18] ;
 wire \tholin_riscv.regs[24][19] ;
 wire \tholin_riscv.regs[24][1] ;
 wire \tholin_riscv.regs[24][20] ;
 wire \tholin_riscv.regs[24][21] ;
 wire \tholin_riscv.regs[24][22] ;
 wire \tholin_riscv.regs[24][23] ;
 wire \tholin_riscv.regs[24][24] ;
 wire \tholin_riscv.regs[24][25] ;
 wire \tholin_riscv.regs[24][26] ;
 wire \tholin_riscv.regs[24][27] ;
 wire \tholin_riscv.regs[24][28] ;
 wire \tholin_riscv.regs[24][29] ;
 wire \tholin_riscv.regs[24][2] ;
 wire \tholin_riscv.regs[24][30] ;
 wire \tholin_riscv.regs[24][31] ;
 wire \tholin_riscv.regs[24][3] ;
 wire \tholin_riscv.regs[24][4] ;
 wire \tholin_riscv.regs[24][5] ;
 wire \tholin_riscv.regs[24][6] ;
 wire \tholin_riscv.regs[24][7] ;
 wire \tholin_riscv.regs[24][8] ;
 wire \tholin_riscv.regs[24][9] ;
 wire \tholin_riscv.regs[25][0] ;
 wire \tholin_riscv.regs[25][10] ;
 wire \tholin_riscv.regs[25][11] ;
 wire \tholin_riscv.regs[25][12] ;
 wire \tholin_riscv.regs[25][13] ;
 wire \tholin_riscv.regs[25][14] ;
 wire \tholin_riscv.regs[25][15] ;
 wire \tholin_riscv.regs[25][16] ;
 wire \tholin_riscv.regs[25][17] ;
 wire \tholin_riscv.regs[25][18] ;
 wire \tholin_riscv.regs[25][19] ;
 wire \tholin_riscv.regs[25][1] ;
 wire \tholin_riscv.regs[25][20] ;
 wire \tholin_riscv.regs[25][21] ;
 wire \tholin_riscv.regs[25][22] ;
 wire \tholin_riscv.regs[25][23] ;
 wire \tholin_riscv.regs[25][24] ;
 wire \tholin_riscv.regs[25][25] ;
 wire \tholin_riscv.regs[25][26] ;
 wire \tholin_riscv.regs[25][27] ;
 wire \tholin_riscv.regs[25][28] ;
 wire \tholin_riscv.regs[25][29] ;
 wire \tholin_riscv.regs[25][2] ;
 wire \tholin_riscv.regs[25][30] ;
 wire \tholin_riscv.regs[25][31] ;
 wire \tholin_riscv.regs[25][3] ;
 wire \tholin_riscv.regs[25][4] ;
 wire \tholin_riscv.regs[25][5] ;
 wire \tholin_riscv.regs[25][6] ;
 wire \tholin_riscv.regs[25][7] ;
 wire \tholin_riscv.regs[25][8] ;
 wire \tholin_riscv.regs[25][9] ;
 wire \tholin_riscv.regs[26][0] ;
 wire \tholin_riscv.regs[26][10] ;
 wire \tholin_riscv.regs[26][11] ;
 wire \tholin_riscv.regs[26][12] ;
 wire \tholin_riscv.regs[26][13] ;
 wire \tholin_riscv.regs[26][14] ;
 wire \tholin_riscv.regs[26][15] ;
 wire \tholin_riscv.regs[26][16] ;
 wire \tholin_riscv.regs[26][17] ;
 wire \tholin_riscv.regs[26][18] ;
 wire \tholin_riscv.regs[26][19] ;
 wire \tholin_riscv.regs[26][1] ;
 wire \tholin_riscv.regs[26][20] ;
 wire \tholin_riscv.regs[26][21] ;
 wire \tholin_riscv.regs[26][22] ;
 wire \tholin_riscv.regs[26][23] ;
 wire \tholin_riscv.regs[26][24] ;
 wire \tholin_riscv.regs[26][25] ;
 wire \tholin_riscv.regs[26][26] ;
 wire \tholin_riscv.regs[26][27] ;
 wire \tholin_riscv.regs[26][28] ;
 wire \tholin_riscv.regs[26][29] ;
 wire \tholin_riscv.regs[26][2] ;
 wire \tholin_riscv.regs[26][30] ;
 wire \tholin_riscv.regs[26][31] ;
 wire \tholin_riscv.regs[26][3] ;
 wire \tholin_riscv.regs[26][4] ;
 wire \tholin_riscv.regs[26][5] ;
 wire \tholin_riscv.regs[26][6] ;
 wire \tholin_riscv.regs[26][7] ;
 wire \tholin_riscv.regs[26][8] ;
 wire \tholin_riscv.regs[26][9] ;
 wire \tholin_riscv.regs[27][0] ;
 wire \tholin_riscv.regs[27][10] ;
 wire \tholin_riscv.regs[27][11] ;
 wire \tholin_riscv.regs[27][12] ;
 wire \tholin_riscv.regs[27][13] ;
 wire \tholin_riscv.regs[27][14] ;
 wire \tholin_riscv.regs[27][15] ;
 wire \tholin_riscv.regs[27][16] ;
 wire \tholin_riscv.regs[27][17] ;
 wire \tholin_riscv.regs[27][18] ;
 wire \tholin_riscv.regs[27][19] ;
 wire \tholin_riscv.regs[27][1] ;
 wire \tholin_riscv.regs[27][20] ;
 wire \tholin_riscv.regs[27][21] ;
 wire \tholin_riscv.regs[27][22] ;
 wire \tholin_riscv.regs[27][23] ;
 wire \tholin_riscv.regs[27][24] ;
 wire \tholin_riscv.regs[27][25] ;
 wire \tholin_riscv.regs[27][26] ;
 wire \tholin_riscv.regs[27][27] ;
 wire \tholin_riscv.regs[27][28] ;
 wire \tholin_riscv.regs[27][29] ;
 wire \tholin_riscv.regs[27][2] ;
 wire \tholin_riscv.regs[27][30] ;
 wire \tholin_riscv.regs[27][31] ;
 wire \tholin_riscv.regs[27][3] ;
 wire \tholin_riscv.regs[27][4] ;
 wire \tholin_riscv.regs[27][5] ;
 wire \tholin_riscv.regs[27][6] ;
 wire \tholin_riscv.regs[27][7] ;
 wire \tholin_riscv.regs[27][8] ;
 wire \tholin_riscv.regs[27][9] ;
 wire \tholin_riscv.regs[28][0] ;
 wire \tholin_riscv.regs[28][10] ;
 wire \tholin_riscv.regs[28][11] ;
 wire \tholin_riscv.regs[28][12] ;
 wire \tholin_riscv.regs[28][13] ;
 wire \tholin_riscv.regs[28][14] ;
 wire \tholin_riscv.regs[28][15] ;
 wire \tholin_riscv.regs[28][16] ;
 wire \tholin_riscv.regs[28][17] ;
 wire \tholin_riscv.regs[28][18] ;
 wire \tholin_riscv.regs[28][19] ;
 wire \tholin_riscv.regs[28][1] ;
 wire \tholin_riscv.regs[28][20] ;
 wire \tholin_riscv.regs[28][21] ;
 wire \tholin_riscv.regs[28][22] ;
 wire \tholin_riscv.regs[28][23] ;
 wire \tholin_riscv.regs[28][24] ;
 wire \tholin_riscv.regs[28][25] ;
 wire \tholin_riscv.regs[28][26] ;
 wire \tholin_riscv.regs[28][27] ;
 wire \tholin_riscv.regs[28][28] ;
 wire \tholin_riscv.regs[28][29] ;
 wire \tholin_riscv.regs[28][2] ;
 wire \tholin_riscv.regs[28][30] ;
 wire \tholin_riscv.regs[28][31] ;
 wire \tholin_riscv.regs[28][3] ;
 wire \tholin_riscv.regs[28][4] ;
 wire \tholin_riscv.regs[28][5] ;
 wire \tholin_riscv.regs[28][6] ;
 wire \tholin_riscv.regs[28][7] ;
 wire \tholin_riscv.regs[28][8] ;
 wire \tholin_riscv.regs[28][9] ;
 wire \tholin_riscv.regs[29][0] ;
 wire \tholin_riscv.regs[29][10] ;
 wire \tholin_riscv.regs[29][11] ;
 wire \tholin_riscv.regs[29][12] ;
 wire \tholin_riscv.regs[29][13] ;
 wire \tholin_riscv.regs[29][14] ;
 wire \tholin_riscv.regs[29][15] ;
 wire \tholin_riscv.regs[29][16] ;
 wire \tholin_riscv.regs[29][17] ;
 wire \tholin_riscv.regs[29][18] ;
 wire \tholin_riscv.regs[29][19] ;
 wire \tholin_riscv.regs[29][1] ;
 wire \tholin_riscv.regs[29][20] ;
 wire \tholin_riscv.regs[29][21] ;
 wire \tholin_riscv.regs[29][22] ;
 wire \tholin_riscv.regs[29][23] ;
 wire \tholin_riscv.regs[29][24] ;
 wire \tholin_riscv.regs[29][25] ;
 wire \tholin_riscv.regs[29][26] ;
 wire \tholin_riscv.regs[29][27] ;
 wire \tholin_riscv.regs[29][28] ;
 wire \tholin_riscv.regs[29][29] ;
 wire \tholin_riscv.regs[29][2] ;
 wire \tholin_riscv.regs[29][30] ;
 wire \tholin_riscv.regs[29][31] ;
 wire \tholin_riscv.regs[29][3] ;
 wire \tholin_riscv.regs[29][4] ;
 wire \tholin_riscv.regs[29][5] ;
 wire \tholin_riscv.regs[29][6] ;
 wire \tholin_riscv.regs[29][7] ;
 wire \tholin_riscv.regs[29][8] ;
 wire \tholin_riscv.regs[29][9] ;
 wire \tholin_riscv.regs[2][0] ;
 wire \tholin_riscv.regs[2][10] ;
 wire \tholin_riscv.regs[2][11] ;
 wire \tholin_riscv.regs[2][12] ;
 wire \tholin_riscv.regs[2][13] ;
 wire \tholin_riscv.regs[2][14] ;
 wire \tholin_riscv.regs[2][15] ;
 wire \tholin_riscv.regs[2][16] ;
 wire \tholin_riscv.regs[2][17] ;
 wire \tholin_riscv.regs[2][18] ;
 wire \tholin_riscv.regs[2][19] ;
 wire \tholin_riscv.regs[2][1] ;
 wire \tholin_riscv.regs[2][20] ;
 wire \tholin_riscv.regs[2][21] ;
 wire \tholin_riscv.regs[2][22] ;
 wire \tholin_riscv.regs[2][23] ;
 wire \tholin_riscv.regs[2][24] ;
 wire \tholin_riscv.regs[2][25] ;
 wire \tholin_riscv.regs[2][26] ;
 wire \tholin_riscv.regs[2][27] ;
 wire \tholin_riscv.regs[2][28] ;
 wire \tholin_riscv.regs[2][29] ;
 wire \tholin_riscv.regs[2][2] ;
 wire \tholin_riscv.regs[2][30] ;
 wire \tholin_riscv.regs[2][31] ;
 wire \tholin_riscv.regs[2][3] ;
 wire \tholin_riscv.regs[2][4] ;
 wire \tholin_riscv.regs[2][5] ;
 wire \tholin_riscv.regs[2][6] ;
 wire \tholin_riscv.regs[2][7] ;
 wire \tholin_riscv.regs[2][8] ;
 wire \tholin_riscv.regs[2][9] ;
 wire \tholin_riscv.regs[30][0] ;
 wire \tholin_riscv.regs[30][10] ;
 wire \tholin_riscv.regs[30][11] ;
 wire \tholin_riscv.regs[30][12] ;
 wire \tholin_riscv.regs[30][13] ;
 wire \tholin_riscv.regs[30][14] ;
 wire \tholin_riscv.regs[30][15] ;
 wire \tholin_riscv.regs[30][16] ;
 wire \tholin_riscv.regs[30][17] ;
 wire \tholin_riscv.regs[30][18] ;
 wire \tholin_riscv.regs[30][19] ;
 wire \tholin_riscv.regs[30][1] ;
 wire \tholin_riscv.regs[30][20] ;
 wire \tholin_riscv.regs[30][21] ;
 wire \tholin_riscv.regs[30][22] ;
 wire \tholin_riscv.regs[30][23] ;
 wire \tholin_riscv.regs[30][24] ;
 wire \tholin_riscv.regs[30][25] ;
 wire \tholin_riscv.regs[30][26] ;
 wire \tholin_riscv.regs[30][27] ;
 wire \tholin_riscv.regs[30][28] ;
 wire \tholin_riscv.regs[30][29] ;
 wire \tholin_riscv.regs[30][2] ;
 wire \tholin_riscv.regs[30][30] ;
 wire \tholin_riscv.regs[30][31] ;
 wire \tholin_riscv.regs[30][3] ;
 wire \tholin_riscv.regs[30][4] ;
 wire \tholin_riscv.regs[30][5] ;
 wire \tholin_riscv.regs[30][6] ;
 wire \tholin_riscv.regs[30][7] ;
 wire \tholin_riscv.regs[30][8] ;
 wire \tholin_riscv.regs[30][9] ;
 wire \tholin_riscv.regs[31][0] ;
 wire \tholin_riscv.regs[31][10] ;
 wire \tholin_riscv.regs[31][11] ;
 wire \tholin_riscv.regs[31][12] ;
 wire \tholin_riscv.regs[31][13] ;
 wire \tholin_riscv.regs[31][14] ;
 wire \tholin_riscv.regs[31][15] ;
 wire \tholin_riscv.regs[31][16] ;
 wire \tholin_riscv.regs[31][17] ;
 wire \tholin_riscv.regs[31][18] ;
 wire \tholin_riscv.regs[31][19] ;
 wire \tholin_riscv.regs[31][1] ;
 wire \tholin_riscv.regs[31][20] ;
 wire \tholin_riscv.regs[31][21] ;
 wire \tholin_riscv.regs[31][22] ;
 wire \tholin_riscv.regs[31][23] ;
 wire \tholin_riscv.regs[31][24] ;
 wire \tholin_riscv.regs[31][25] ;
 wire \tholin_riscv.regs[31][26] ;
 wire \tholin_riscv.regs[31][27] ;
 wire \tholin_riscv.regs[31][28] ;
 wire \tholin_riscv.regs[31][29] ;
 wire \tholin_riscv.regs[31][2] ;
 wire \tholin_riscv.regs[31][30] ;
 wire \tholin_riscv.regs[31][31] ;
 wire \tholin_riscv.regs[31][3] ;
 wire \tholin_riscv.regs[31][4] ;
 wire \tholin_riscv.regs[31][5] ;
 wire \tholin_riscv.regs[31][6] ;
 wire \tholin_riscv.regs[31][7] ;
 wire \tholin_riscv.regs[31][8] ;
 wire \tholin_riscv.regs[31][9] ;
 wire \tholin_riscv.regs[3][0] ;
 wire \tholin_riscv.regs[3][10] ;
 wire \tholin_riscv.regs[3][11] ;
 wire \tholin_riscv.regs[3][12] ;
 wire \tholin_riscv.regs[3][13] ;
 wire \tholin_riscv.regs[3][14] ;
 wire \tholin_riscv.regs[3][15] ;
 wire \tholin_riscv.regs[3][16] ;
 wire \tholin_riscv.regs[3][17] ;
 wire \tholin_riscv.regs[3][18] ;
 wire \tholin_riscv.regs[3][19] ;
 wire \tholin_riscv.regs[3][1] ;
 wire \tholin_riscv.regs[3][20] ;
 wire \tholin_riscv.regs[3][21] ;
 wire \tholin_riscv.regs[3][22] ;
 wire \tholin_riscv.regs[3][23] ;
 wire \tholin_riscv.regs[3][24] ;
 wire \tholin_riscv.regs[3][25] ;
 wire \tholin_riscv.regs[3][26] ;
 wire \tholin_riscv.regs[3][27] ;
 wire \tholin_riscv.regs[3][28] ;
 wire \tholin_riscv.regs[3][29] ;
 wire \tholin_riscv.regs[3][2] ;
 wire \tholin_riscv.regs[3][30] ;
 wire \tholin_riscv.regs[3][31] ;
 wire \tholin_riscv.regs[3][3] ;
 wire \tholin_riscv.regs[3][4] ;
 wire \tholin_riscv.regs[3][5] ;
 wire \tholin_riscv.regs[3][6] ;
 wire \tholin_riscv.regs[3][7] ;
 wire \tholin_riscv.regs[3][8] ;
 wire \tholin_riscv.regs[3][9] ;
 wire \tholin_riscv.regs[4][0] ;
 wire \tholin_riscv.regs[4][10] ;
 wire \tholin_riscv.regs[4][11] ;
 wire \tholin_riscv.regs[4][12] ;
 wire \tholin_riscv.regs[4][13] ;
 wire \tholin_riscv.regs[4][14] ;
 wire \tholin_riscv.regs[4][15] ;
 wire \tholin_riscv.regs[4][16] ;
 wire \tholin_riscv.regs[4][17] ;
 wire \tholin_riscv.regs[4][18] ;
 wire \tholin_riscv.regs[4][19] ;
 wire \tholin_riscv.regs[4][1] ;
 wire \tholin_riscv.regs[4][20] ;
 wire \tholin_riscv.regs[4][21] ;
 wire \tholin_riscv.regs[4][22] ;
 wire \tholin_riscv.regs[4][23] ;
 wire \tholin_riscv.regs[4][24] ;
 wire \tholin_riscv.regs[4][25] ;
 wire \tholin_riscv.regs[4][26] ;
 wire \tholin_riscv.regs[4][27] ;
 wire \tholin_riscv.regs[4][28] ;
 wire \tholin_riscv.regs[4][29] ;
 wire \tholin_riscv.regs[4][2] ;
 wire \tholin_riscv.regs[4][30] ;
 wire \tholin_riscv.regs[4][31] ;
 wire \tholin_riscv.regs[4][3] ;
 wire \tholin_riscv.regs[4][4] ;
 wire \tholin_riscv.regs[4][5] ;
 wire \tholin_riscv.regs[4][6] ;
 wire \tholin_riscv.regs[4][7] ;
 wire \tholin_riscv.regs[4][8] ;
 wire \tholin_riscv.regs[4][9] ;
 wire \tholin_riscv.regs[5][0] ;
 wire \tholin_riscv.regs[5][10] ;
 wire \tholin_riscv.regs[5][11] ;
 wire \tholin_riscv.regs[5][12] ;
 wire \tholin_riscv.regs[5][13] ;
 wire \tholin_riscv.regs[5][14] ;
 wire \tholin_riscv.regs[5][15] ;
 wire \tholin_riscv.regs[5][16] ;
 wire \tholin_riscv.regs[5][17] ;
 wire \tholin_riscv.regs[5][18] ;
 wire \tholin_riscv.regs[5][19] ;
 wire \tholin_riscv.regs[5][1] ;
 wire \tholin_riscv.regs[5][20] ;
 wire \tholin_riscv.regs[5][21] ;
 wire \tholin_riscv.regs[5][22] ;
 wire \tholin_riscv.regs[5][23] ;
 wire \tholin_riscv.regs[5][24] ;
 wire \tholin_riscv.regs[5][25] ;
 wire \tholin_riscv.regs[5][26] ;
 wire \tholin_riscv.regs[5][27] ;
 wire \tholin_riscv.regs[5][28] ;
 wire \tholin_riscv.regs[5][29] ;
 wire \tholin_riscv.regs[5][2] ;
 wire \tholin_riscv.regs[5][30] ;
 wire \tholin_riscv.regs[5][31] ;
 wire \tholin_riscv.regs[5][3] ;
 wire \tholin_riscv.regs[5][4] ;
 wire \tholin_riscv.regs[5][5] ;
 wire \tholin_riscv.regs[5][6] ;
 wire \tholin_riscv.regs[5][7] ;
 wire \tholin_riscv.regs[5][8] ;
 wire \tholin_riscv.regs[5][9] ;
 wire \tholin_riscv.regs[6][0] ;
 wire \tholin_riscv.regs[6][10] ;
 wire \tholin_riscv.regs[6][11] ;
 wire \tholin_riscv.regs[6][12] ;
 wire \tholin_riscv.regs[6][13] ;
 wire \tholin_riscv.regs[6][14] ;
 wire \tholin_riscv.regs[6][15] ;
 wire \tholin_riscv.regs[6][16] ;
 wire \tholin_riscv.regs[6][17] ;
 wire \tholin_riscv.regs[6][18] ;
 wire \tholin_riscv.regs[6][19] ;
 wire \tholin_riscv.regs[6][1] ;
 wire \tholin_riscv.regs[6][20] ;
 wire \tholin_riscv.regs[6][21] ;
 wire \tholin_riscv.regs[6][22] ;
 wire \tholin_riscv.regs[6][23] ;
 wire \tholin_riscv.regs[6][24] ;
 wire \tholin_riscv.regs[6][25] ;
 wire \tholin_riscv.regs[6][26] ;
 wire \tholin_riscv.regs[6][27] ;
 wire \tholin_riscv.regs[6][28] ;
 wire \tholin_riscv.regs[6][29] ;
 wire \tholin_riscv.regs[6][2] ;
 wire \tholin_riscv.regs[6][30] ;
 wire \tholin_riscv.regs[6][31] ;
 wire \tholin_riscv.regs[6][3] ;
 wire \tholin_riscv.regs[6][4] ;
 wire \tholin_riscv.regs[6][5] ;
 wire \tholin_riscv.regs[6][6] ;
 wire \tholin_riscv.regs[6][7] ;
 wire \tholin_riscv.regs[6][8] ;
 wire \tholin_riscv.regs[6][9] ;
 wire \tholin_riscv.regs[7][0] ;
 wire \tholin_riscv.regs[7][10] ;
 wire \tholin_riscv.regs[7][11] ;
 wire \tholin_riscv.regs[7][12] ;
 wire \tholin_riscv.regs[7][13] ;
 wire \tholin_riscv.regs[7][14] ;
 wire \tholin_riscv.regs[7][15] ;
 wire \tholin_riscv.regs[7][16] ;
 wire \tholin_riscv.regs[7][17] ;
 wire \tholin_riscv.regs[7][18] ;
 wire \tholin_riscv.regs[7][19] ;
 wire \tholin_riscv.regs[7][1] ;
 wire \tholin_riscv.regs[7][20] ;
 wire \tholin_riscv.regs[7][21] ;
 wire \tholin_riscv.regs[7][22] ;
 wire \tholin_riscv.regs[7][23] ;
 wire \tholin_riscv.regs[7][24] ;
 wire \tholin_riscv.regs[7][25] ;
 wire \tholin_riscv.regs[7][26] ;
 wire \tholin_riscv.regs[7][27] ;
 wire \tholin_riscv.regs[7][28] ;
 wire \tholin_riscv.regs[7][29] ;
 wire \tholin_riscv.regs[7][2] ;
 wire \tholin_riscv.regs[7][30] ;
 wire \tholin_riscv.regs[7][31] ;
 wire \tholin_riscv.regs[7][3] ;
 wire \tholin_riscv.regs[7][4] ;
 wire \tholin_riscv.regs[7][5] ;
 wire \tholin_riscv.regs[7][6] ;
 wire \tholin_riscv.regs[7][7] ;
 wire \tholin_riscv.regs[7][8] ;
 wire \tholin_riscv.regs[7][9] ;
 wire \tholin_riscv.regs[8][0] ;
 wire \tholin_riscv.regs[8][10] ;
 wire \tholin_riscv.regs[8][11] ;
 wire \tholin_riscv.regs[8][12] ;
 wire \tholin_riscv.regs[8][13] ;
 wire \tholin_riscv.regs[8][14] ;
 wire \tholin_riscv.regs[8][15] ;
 wire \tholin_riscv.regs[8][16] ;
 wire \tholin_riscv.regs[8][17] ;
 wire \tholin_riscv.regs[8][18] ;
 wire \tholin_riscv.regs[8][19] ;
 wire \tholin_riscv.regs[8][1] ;
 wire \tholin_riscv.regs[8][20] ;
 wire \tholin_riscv.regs[8][21] ;
 wire \tholin_riscv.regs[8][22] ;
 wire \tholin_riscv.regs[8][23] ;
 wire \tholin_riscv.regs[8][24] ;
 wire \tholin_riscv.regs[8][25] ;
 wire \tholin_riscv.regs[8][26] ;
 wire \tholin_riscv.regs[8][27] ;
 wire \tholin_riscv.regs[8][28] ;
 wire \tholin_riscv.regs[8][29] ;
 wire \tholin_riscv.regs[8][2] ;
 wire \tholin_riscv.regs[8][30] ;
 wire \tholin_riscv.regs[8][31] ;
 wire \tholin_riscv.regs[8][3] ;
 wire \tholin_riscv.regs[8][4] ;
 wire \tholin_riscv.regs[8][5] ;
 wire \tholin_riscv.regs[8][6] ;
 wire \tholin_riscv.regs[8][7] ;
 wire \tholin_riscv.regs[8][8] ;
 wire \tholin_riscv.regs[8][9] ;
 wire \tholin_riscv.regs[9][0] ;
 wire \tholin_riscv.regs[9][10] ;
 wire \tholin_riscv.regs[9][11] ;
 wire \tholin_riscv.regs[9][12] ;
 wire \tholin_riscv.regs[9][13] ;
 wire \tholin_riscv.regs[9][14] ;
 wire \tholin_riscv.regs[9][15] ;
 wire \tholin_riscv.regs[9][16] ;
 wire \tholin_riscv.regs[9][17] ;
 wire \tholin_riscv.regs[9][18] ;
 wire \tholin_riscv.regs[9][19] ;
 wire \tholin_riscv.regs[9][1] ;
 wire \tholin_riscv.regs[9][20] ;
 wire \tholin_riscv.regs[9][21] ;
 wire \tholin_riscv.regs[9][22] ;
 wire \tholin_riscv.regs[9][23] ;
 wire \tholin_riscv.regs[9][24] ;
 wire \tholin_riscv.regs[9][25] ;
 wire \tholin_riscv.regs[9][26] ;
 wire \tholin_riscv.regs[9][27] ;
 wire \tholin_riscv.regs[9][28] ;
 wire \tholin_riscv.regs[9][29] ;
 wire \tholin_riscv.regs[9][2] ;
 wire \tholin_riscv.regs[9][30] ;
 wire \tholin_riscv.regs[9][31] ;
 wire \tholin_riscv.regs[9][3] ;
 wire \tholin_riscv.regs[9][4] ;
 wire \tholin_riscv.regs[9][5] ;
 wire \tholin_riscv.regs[9][6] ;
 wire \tholin_riscv.regs[9][7] ;
 wire \tholin_riscv.regs[9][8] ;
 wire \tholin_riscv.regs[9][9] ;
 wire \tholin_riscv.requested_addr[0] ;
 wire \tholin_riscv.requested_addr[10] ;
 wire \tholin_riscv.requested_addr[11] ;
 wire \tholin_riscv.requested_addr[12] ;
 wire \tholin_riscv.requested_addr[13] ;
 wire \tholin_riscv.requested_addr[14] ;
 wire \tholin_riscv.requested_addr[15] ;
 wire \tholin_riscv.requested_addr[16] ;
 wire \tholin_riscv.requested_addr[17] ;
 wire \tholin_riscv.requested_addr[18] ;
 wire \tholin_riscv.requested_addr[19] ;
 wire \tholin_riscv.requested_addr[1] ;
 wire \tholin_riscv.requested_addr[20] ;
 wire \tholin_riscv.requested_addr[21] ;
 wire \tholin_riscv.requested_addr[22] ;
 wire \tholin_riscv.requested_addr[23] ;
 wire \tholin_riscv.requested_addr[24] ;
 wire \tholin_riscv.requested_addr[25] ;
 wire \tholin_riscv.requested_addr[26] ;
 wire \tholin_riscv.requested_addr[27] ;
 wire \tholin_riscv.requested_addr[28] ;
 wire \tholin_riscv.requested_addr[29] ;
 wire \tholin_riscv.requested_addr[2] ;
 wire \tholin_riscv.requested_addr[30] ;
 wire \tholin_riscv.requested_addr[31] ;
 wire \tholin_riscv.requested_addr[3] ;
 wire \tholin_riscv.requested_addr[4] ;
 wire \tholin_riscv.requested_addr[5] ;
 wire \tholin_riscv.requested_addr[6] ;
 wire \tholin_riscv.requested_addr[7] ;
 wire \tholin_riscv.requested_addr[8] ;
 wire \tholin_riscv.requested_addr[9] ;
 wire \tholin_riscv.ret_cycle[0] ;
 wire \tholin_riscv.ret_cycle[1] ;
 wire \tholin_riscv.spi.busy ;
 wire \tholin_riscv.spi.counter[0] ;
 wire \tholin_riscv.spi.counter[1] ;
 wire \tholin_riscv.spi.counter[2] ;
 wire \tholin_riscv.spi.counter[3] ;
 wire \tholin_riscv.spi.counter[4] ;
 wire \tholin_riscv.spi.data_in_buff[0] ;
 wire \tholin_riscv.spi.data_in_buff[1] ;
 wire \tholin_riscv.spi.data_in_buff[2] ;
 wire \tholin_riscv.spi.data_in_buff[3] ;
 wire \tholin_riscv.spi.data_in_buff[4] ;
 wire \tholin_riscv.spi.data_in_buff[5] ;
 wire \tholin_riscv.spi.data_in_buff[6] ;
 wire \tholin_riscv.spi.data_in_buff[7] ;
 wire \tholin_riscv.spi.data_out_buff[0] ;
 wire \tholin_riscv.spi.data_out_buff[1] ;
 wire \tholin_riscv.spi.data_out_buff[2] ;
 wire \tholin_riscv.spi.data_out_buff[3] ;
 wire \tholin_riscv.spi.data_out_buff[4] ;
 wire \tholin_riscv.spi.data_out_buff[5] ;
 wire \tholin_riscv.spi.data_out_buff[6] ;
 wire \tholin_riscv.spi.data_out_buff[7] ;
 wire \tholin_riscv.spi.div_counter[0] ;
 wire \tholin_riscv.spi.div_counter[1] ;
 wire \tholin_riscv.spi.div_counter[2] ;
 wire \tholin_riscv.spi.div_counter[3] ;
 wire \tholin_riscv.spi.div_counter[4] ;
 wire \tholin_riscv.spi.div_counter[5] ;
 wire \tholin_riscv.spi.div_counter[6] ;
 wire \tholin_riscv.spi.div_counter[7] ;
 wire \tholin_riscv.spi.divisor[0] ;
 wire \tholin_riscv.spi.divisor[1] ;
 wire \tholin_riscv.spi.divisor[2] ;
 wire \tholin_riscv.spi.divisor[3] ;
 wire \tholin_riscv.spi.divisor[4] ;
 wire \tholin_riscv.spi.divisor[5] ;
 wire \tholin_riscv.spi.divisor[6] ;
 wire \tholin_riscv.spi.divisor[7] ;
 wire \tholin_riscv.spi.dout[0] ;
 wire \tholin_riscv.spi.dout[1] ;
 wire \tholin_riscv.spi.dout[2] ;
 wire \tholin_riscv.spi.dout[3] ;
 wire \tholin_riscv.spi.dout[4] ;
 wire \tholin_riscv.spi.dout[5] ;
 wire \tholin_riscv.spi.dout[6] ;
 wire \tholin_riscv.spi.dout[7] ;
 wire \tholin_riscv.timer_int_enable ;
 wire \tholin_riscv.tmr0[0] ;
 wire \tholin_riscv.tmr0[10] ;
 wire \tholin_riscv.tmr0[11] ;
 wire \tholin_riscv.tmr0[12] ;
 wire \tholin_riscv.tmr0[13] ;
 wire \tholin_riscv.tmr0[14] ;
 wire \tholin_riscv.tmr0[15] ;
 wire \tholin_riscv.tmr0[16] ;
 wire \tholin_riscv.tmr0[17] ;
 wire \tholin_riscv.tmr0[18] ;
 wire \tholin_riscv.tmr0[19] ;
 wire \tholin_riscv.tmr0[1] ;
 wire \tholin_riscv.tmr0[20] ;
 wire \tholin_riscv.tmr0[21] ;
 wire \tholin_riscv.tmr0[22] ;
 wire \tholin_riscv.tmr0[23] ;
 wire \tholin_riscv.tmr0[24] ;
 wire \tholin_riscv.tmr0[25] ;
 wire \tholin_riscv.tmr0[26] ;
 wire \tholin_riscv.tmr0[27] ;
 wire \tholin_riscv.tmr0[28] ;
 wire \tholin_riscv.tmr0[29] ;
 wire \tholin_riscv.tmr0[2] ;
 wire \tholin_riscv.tmr0[30] ;
 wire \tholin_riscv.tmr0[31] ;
 wire \tholin_riscv.tmr0[3] ;
 wire \tholin_riscv.tmr0[4] ;
 wire \tholin_riscv.tmr0[5] ;
 wire \tholin_riscv.tmr0[6] ;
 wire \tholin_riscv.tmr0[7] ;
 wire \tholin_riscv.tmr0[8] ;
 wire \tholin_riscv.tmr0[9] ;
 wire \tholin_riscv.tmr0_pre[0] ;
 wire \tholin_riscv.tmr0_pre[10] ;
 wire \tholin_riscv.tmr0_pre[11] ;
 wire \tholin_riscv.tmr0_pre[12] ;
 wire \tholin_riscv.tmr0_pre[13] ;
 wire \tholin_riscv.tmr0_pre[14] ;
 wire \tholin_riscv.tmr0_pre[15] ;
 wire \tholin_riscv.tmr0_pre[16] ;
 wire \tholin_riscv.tmr0_pre[17] ;
 wire \tholin_riscv.tmr0_pre[18] ;
 wire \tholin_riscv.tmr0_pre[19] ;
 wire \tholin_riscv.tmr0_pre[1] ;
 wire \tholin_riscv.tmr0_pre[20] ;
 wire \tholin_riscv.tmr0_pre[21] ;
 wire \tholin_riscv.tmr0_pre[22] ;
 wire \tholin_riscv.tmr0_pre[23] ;
 wire \tholin_riscv.tmr0_pre[24] ;
 wire \tholin_riscv.tmr0_pre[25] ;
 wire \tholin_riscv.tmr0_pre[26] ;
 wire \tholin_riscv.tmr0_pre[27] ;
 wire \tholin_riscv.tmr0_pre[28] ;
 wire \tholin_riscv.tmr0_pre[29] ;
 wire \tholin_riscv.tmr0_pre[2] ;
 wire \tholin_riscv.tmr0_pre[30] ;
 wire \tholin_riscv.tmr0_pre[31] ;
 wire \tholin_riscv.tmr0_pre[3] ;
 wire \tholin_riscv.tmr0_pre[4] ;
 wire \tholin_riscv.tmr0_pre[5] ;
 wire \tholin_riscv.tmr0_pre[6] ;
 wire \tholin_riscv.tmr0_pre[7] ;
 wire \tholin_riscv.tmr0_pre[8] ;
 wire \tholin_riscv.tmr0_pre[9] ;
 wire \tholin_riscv.tmr0_pre_ctr[0] ;
 wire \tholin_riscv.tmr0_pre_ctr[10] ;
 wire \tholin_riscv.tmr0_pre_ctr[11] ;
 wire \tholin_riscv.tmr0_pre_ctr[12] ;
 wire \tholin_riscv.tmr0_pre_ctr[13] ;
 wire \tholin_riscv.tmr0_pre_ctr[14] ;
 wire \tholin_riscv.tmr0_pre_ctr[15] ;
 wire \tholin_riscv.tmr0_pre_ctr[16] ;
 wire \tholin_riscv.tmr0_pre_ctr[17] ;
 wire \tholin_riscv.tmr0_pre_ctr[18] ;
 wire \tholin_riscv.tmr0_pre_ctr[19] ;
 wire \tholin_riscv.tmr0_pre_ctr[1] ;
 wire \tholin_riscv.tmr0_pre_ctr[20] ;
 wire \tholin_riscv.tmr0_pre_ctr[21] ;
 wire \tholin_riscv.tmr0_pre_ctr[22] ;
 wire \tholin_riscv.tmr0_pre_ctr[23] ;
 wire \tholin_riscv.tmr0_pre_ctr[24] ;
 wire \tholin_riscv.tmr0_pre_ctr[25] ;
 wire \tholin_riscv.tmr0_pre_ctr[26] ;
 wire \tholin_riscv.tmr0_pre_ctr[27] ;
 wire \tholin_riscv.tmr0_pre_ctr[28] ;
 wire \tholin_riscv.tmr0_pre_ctr[29] ;
 wire \tholin_riscv.tmr0_pre_ctr[2] ;
 wire \tholin_riscv.tmr0_pre_ctr[30] ;
 wire \tholin_riscv.tmr0_pre_ctr[31] ;
 wire \tholin_riscv.tmr0_pre_ctr[3] ;
 wire \tholin_riscv.tmr0_pre_ctr[4] ;
 wire \tholin_riscv.tmr0_pre_ctr[5] ;
 wire \tholin_riscv.tmr0_pre_ctr[6] ;
 wire \tholin_riscv.tmr0_pre_ctr[7] ;
 wire \tholin_riscv.tmr0_pre_ctr[8] ;
 wire \tholin_riscv.tmr0_pre_ctr[9] ;
 wire \tholin_riscv.tmr0_top[0] ;
 wire \tholin_riscv.tmr0_top[10] ;
 wire \tholin_riscv.tmr0_top[11] ;
 wire \tholin_riscv.tmr0_top[12] ;
 wire \tholin_riscv.tmr0_top[13] ;
 wire \tholin_riscv.tmr0_top[14] ;
 wire \tholin_riscv.tmr0_top[15] ;
 wire \tholin_riscv.tmr0_top[16] ;
 wire \tholin_riscv.tmr0_top[17] ;
 wire \tholin_riscv.tmr0_top[18] ;
 wire \tholin_riscv.tmr0_top[19] ;
 wire \tholin_riscv.tmr0_top[1] ;
 wire \tholin_riscv.tmr0_top[20] ;
 wire \tholin_riscv.tmr0_top[21] ;
 wire \tholin_riscv.tmr0_top[22] ;
 wire \tholin_riscv.tmr0_top[23] ;
 wire \tholin_riscv.tmr0_top[24] ;
 wire \tholin_riscv.tmr0_top[25] ;
 wire \tholin_riscv.tmr0_top[26] ;
 wire \tholin_riscv.tmr0_top[27] ;
 wire \tholin_riscv.tmr0_top[28] ;
 wire \tholin_riscv.tmr0_top[29] ;
 wire \tholin_riscv.tmr0_top[2] ;
 wire \tholin_riscv.tmr0_top[30] ;
 wire \tholin_riscv.tmr0_top[31] ;
 wire \tholin_riscv.tmr0_top[3] ;
 wire \tholin_riscv.tmr0_top[4] ;
 wire \tholin_riscv.tmr0_top[5] ;
 wire \tholin_riscv.tmr0_top[6] ;
 wire \tholin_riscv.tmr0_top[7] ;
 wire \tholin_riscv.tmr0_top[8] ;
 wire \tholin_riscv.tmr0_top[9] ;
 wire \tholin_riscv.tmr1[0] ;
 wire \tholin_riscv.tmr1[10] ;
 wire \tholin_riscv.tmr1[11] ;
 wire \tholin_riscv.tmr1[12] ;
 wire \tholin_riscv.tmr1[13] ;
 wire \tholin_riscv.tmr1[14] ;
 wire \tholin_riscv.tmr1[15] ;
 wire \tholin_riscv.tmr1[16] ;
 wire \tholin_riscv.tmr1[17] ;
 wire \tholin_riscv.tmr1[18] ;
 wire \tholin_riscv.tmr1[19] ;
 wire \tholin_riscv.tmr1[1] ;
 wire \tholin_riscv.tmr1[20] ;
 wire \tholin_riscv.tmr1[21] ;
 wire \tholin_riscv.tmr1[22] ;
 wire \tholin_riscv.tmr1[23] ;
 wire \tholin_riscv.tmr1[24] ;
 wire \tholin_riscv.tmr1[25] ;
 wire \tholin_riscv.tmr1[26] ;
 wire \tholin_riscv.tmr1[27] ;
 wire \tholin_riscv.tmr1[28] ;
 wire \tholin_riscv.tmr1[29] ;
 wire \tholin_riscv.tmr1[2] ;
 wire \tholin_riscv.tmr1[30] ;
 wire \tholin_riscv.tmr1[31] ;
 wire \tholin_riscv.tmr1[3] ;
 wire \tholin_riscv.tmr1[4] ;
 wire \tholin_riscv.tmr1[5] ;
 wire \tholin_riscv.tmr1[6] ;
 wire \tholin_riscv.tmr1[7] ;
 wire \tholin_riscv.tmr1[8] ;
 wire \tholin_riscv.tmr1[9] ;
 wire \tholin_riscv.tmr1_pre[0] ;
 wire \tholin_riscv.tmr1_pre[10] ;
 wire \tholin_riscv.tmr1_pre[11] ;
 wire \tholin_riscv.tmr1_pre[12] ;
 wire \tholin_riscv.tmr1_pre[13] ;
 wire \tholin_riscv.tmr1_pre[14] ;
 wire \tholin_riscv.tmr1_pre[15] ;
 wire \tholin_riscv.tmr1_pre[16] ;
 wire \tholin_riscv.tmr1_pre[17] ;
 wire \tholin_riscv.tmr1_pre[18] ;
 wire \tholin_riscv.tmr1_pre[19] ;
 wire \tholin_riscv.tmr1_pre[1] ;
 wire \tholin_riscv.tmr1_pre[20] ;
 wire \tholin_riscv.tmr1_pre[21] ;
 wire \tholin_riscv.tmr1_pre[22] ;
 wire \tholin_riscv.tmr1_pre[23] ;
 wire \tholin_riscv.tmr1_pre[24] ;
 wire \tholin_riscv.tmr1_pre[25] ;
 wire \tholin_riscv.tmr1_pre[26] ;
 wire \tholin_riscv.tmr1_pre[27] ;
 wire \tholin_riscv.tmr1_pre[28] ;
 wire \tholin_riscv.tmr1_pre[29] ;
 wire \tholin_riscv.tmr1_pre[2] ;
 wire \tholin_riscv.tmr1_pre[30] ;
 wire \tholin_riscv.tmr1_pre[31] ;
 wire \tholin_riscv.tmr1_pre[3] ;
 wire \tholin_riscv.tmr1_pre[4] ;
 wire \tholin_riscv.tmr1_pre[5] ;
 wire \tholin_riscv.tmr1_pre[6] ;
 wire \tholin_riscv.tmr1_pre[7] ;
 wire \tholin_riscv.tmr1_pre[8] ;
 wire \tholin_riscv.tmr1_pre[9] ;
 wire \tholin_riscv.tmr1_pre_ctr[0] ;
 wire \tholin_riscv.tmr1_pre_ctr[10] ;
 wire \tholin_riscv.tmr1_pre_ctr[11] ;
 wire \tholin_riscv.tmr1_pre_ctr[12] ;
 wire \tholin_riscv.tmr1_pre_ctr[13] ;
 wire \tholin_riscv.tmr1_pre_ctr[14] ;
 wire \tholin_riscv.tmr1_pre_ctr[15] ;
 wire \tholin_riscv.tmr1_pre_ctr[16] ;
 wire \tholin_riscv.tmr1_pre_ctr[17] ;
 wire \tholin_riscv.tmr1_pre_ctr[18] ;
 wire \tholin_riscv.tmr1_pre_ctr[19] ;
 wire \tholin_riscv.tmr1_pre_ctr[1] ;
 wire \tholin_riscv.tmr1_pre_ctr[20] ;
 wire \tholin_riscv.tmr1_pre_ctr[21] ;
 wire \tholin_riscv.tmr1_pre_ctr[22] ;
 wire \tholin_riscv.tmr1_pre_ctr[23] ;
 wire \tholin_riscv.tmr1_pre_ctr[24] ;
 wire \tholin_riscv.tmr1_pre_ctr[25] ;
 wire \tholin_riscv.tmr1_pre_ctr[26] ;
 wire \tholin_riscv.tmr1_pre_ctr[27] ;
 wire \tholin_riscv.tmr1_pre_ctr[28] ;
 wire \tholin_riscv.tmr1_pre_ctr[29] ;
 wire \tholin_riscv.tmr1_pre_ctr[2] ;
 wire \tholin_riscv.tmr1_pre_ctr[30] ;
 wire \tholin_riscv.tmr1_pre_ctr[31] ;
 wire \tholin_riscv.tmr1_pre_ctr[3] ;
 wire \tholin_riscv.tmr1_pre_ctr[4] ;
 wire \tholin_riscv.tmr1_pre_ctr[5] ;
 wire \tholin_riscv.tmr1_pre_ctr[6] ;
 wire \tholin_riscv.tmr1_pre_ctr[7] ;
 wire \tholin_riscv.tmr1_pre_ctr[8] ;
 wire \tholin_riscv.tmr1_pre_ctr[9] ;
 wire \tholin_riscv.tmr1_top[0] ;
 wire \tholin_riscv.tmr1_top[10] ;
 wire \tholin_riscv.tmr1_top[11] ;
 wire \tholin_riscv.tmr1_top[12] ;
 wire \tholin_riscv.tmr1_top[13] ;
 wire \tholin_riscv.tmr1_top[14] ;
 wire \tholin_riscv.tmr1_top[15] ;
 wire \tholin_riscv.tmr1_top[16] ;
 wire \tholin_riscv.tmr1_top[17] ;
 wire \tholin_riscv.tmr1_top[18] ;
 wire \tholin_riscv.tmr1_top[19] ;
 wire \tholin_riscv.tmr1_top[1] ;
 wire \tholin_riscv.tmr1_top[20] ;
 wire \tholin_riscv.tmr1_top[21] ;
 wire \tholin_riscv.tmr1_top[22] ;
 wire \tholin_riscv.tmr1_top[23] ;
 wire \tholin_riscv.tmr1_top[24] ;
 wire \tholin_riscv.tmr1_top[25] ;
 wire \tholin_riscv.tmr1_top[26] ;
 wire \tholin_riscv.tmr1_top[27] ;
 wire \tholin_riscv.tmr1_top[28] ;
 wire \tholin_riscv.tmr1_top[29] ;
 wire \tholin_riscv.tmr1_top[2] ;
 wire \tholin_riscv.tmr1_top[30] ;
 wire \tholin_riscv.tmr1_top[31] ;
 wire \tholin_riscv.tmr1_top[3] ;
 wire \tholin_riscv.tmr1_top[4] ;
 wire \tholin_riscv.tmr1_top[5] ;
 wire \tholin_riscv.tmr1_top[6] ;
 wire \tholin_riscv.tmr1_top[7] ;
 wire \tholin_riscv.tmr1_top[8] ;
 wire \tholin_riscv.tmr1_top[9] ;
 wire \tholin_riscv.uart.busy ;
 wire \tholin_riscv.uart.counter[0] ;
 wire \tholin_riscv.uart.counter[1] ;
 wire \tholin_riscv.uart.counter[2] ;
 wire \tholin_riscv.uart.counter[3] ;
 wire \tholin_riscv.uart.data_buff[0] ;
 wire \tholin_riscv.uart.data_buff[1] ;
 wire \tholin_riscv.uart.data_buff[2] ;
 wire \tholin_riscv.uart.data_buff[3] ;
 wire \tholin_riscv.uart.data_buff[4] ;
 wire \tholin_riscv.uart.data_buff[5] ;
 wire \tholin_riscv.uart.data_buff[6] ;
 wire \tholin_riscv.uart.data_buff[7] ;
 wire \tholin_riscv.uart.data_buff[8] ;
 wire \tholin_riscv.uart.data_buff[9] ;
 wire \tholin_riscv.uart.div_counter[0] ;
 wire \tholin_riscv.uart.div_counter[10] ;
 wire \tholin_riscv.uart.div_counter[11] ;
 wire \tholin_riscv.uart.div_counter[12] ;
 wire \tholin_riscv.uart.div_counter[13] ;
 wire \tholin_riscv.uart.div_counter[14] ;
 wire \tholin_riscv.uart.div_counter[15] ;
 wire \tholin_riscv.uart.div_counter[1] ;
 wire \tholin_riscv.uart.div_counter[2] ;
 wire \tholin_riscv.uart.div_counter[3] ;
 wire \tholin_riscv.uart.div_counter[4] ;
 wire \tholin_riscv.uart.div_counter[5] ;
 wire \tholin_riscv.uart.div_counter[6] ;
 wire \tholin_riscv.uart.div_counter[7] ;
 wire \tholin_riscv.uart.div_counter[8] ;
 wire \tholin_riscv.uart.div_counter[9] ;
 wire \tholin_riscv.uart.divisor[0] ;
 wire \tholin_riscv.uart.divisor[10] ;
 wire \tholin_riscv.uart.divisor[11] ;
 wire \tholin_riscv.uart.divisor[12] ;
 wire \tholin_riscv.uart.divisor[13] ;
 wire \tholin_riscv.uart.divisor[14] ;
 wire \tholin_riscv.uart.divisor[15] ;
 wire \tholin_riscv.uart.divisor[1] ;
 wire \tholin_riscv.uart.divisor[2] ;
 wire \tholin_riscv.uart.divisor[3] ;
 wire \tholin_riscv.uart.divisor[4] ;
 wire \tholin_riscv.uart.divisor[5] ;
 wire \tholin_riscv.uart.divisor[6] ;
 wire \tholin_riscv.uart.divisor[7] ;
 wire \tholin_riscv.uart.divisor[8] ;
 wire \tholin_riscv.uart.divisor[9] ;
 wire \tholin_riscv.uart.dout[0] ;
 wire \tholin_riscv.uart.dout[1] ;
 wire \tholin_riscv.uart.dout[2] ;
 wire \tholin_riscv.uart.dout[3] ;
 wire \tholin_riscv.uart.dout[4] ;
 wire \tholin_riscv.uart.dout[5] ;
 wire \tholin_riscv.uart.dout[6] ;
 wire \tholin_riscv.uart.dout[7] ;
 wire \tholin_riscv.uart.has_byte ;
 wire \tholin_riscv.uart.receive_buff[0] ;
 wire \tholin_riscv.uart.receive_buff[1] ;
 wire \tholin_riscv.uart.receive_buff[2] ;
 wire \tholin_riscv.uart.receive_buff[3] ;
 wire \tholin_riscv.uart.receive_buff[4] ;
 wire \tholin_riscv.uart.receive_buff[5] ;
 wire \tholin_riscv.uart.receive_buff[6] ;
 wire \tholin_riscv.uart.receive_buff[7] ;
 wire \tholin_riscv.uart.receive_counter[0] ;
 wire \tholin_riscv.uart.receive_counter[1] ;
 wire \tholin_riscv.uart.receive_counter[2] ;
 wire \tholin_riscv.uart.receive_counter[3] ;
 wire \tholin_riscv.uart.receive_div_counter[0] ;
 wire \tholin_riscv.uart.receive_div_counter[10] ;
 wire \tholin_riscv.uart.receive_div_counter[11] ;
 wire \tholin_riscv.uart.receive_div_counter[12] ;
 wire \tholin_riscv.uart.receive_div_counter[13] ;
 wire \tholin_riscv.uart.receive_div_counter[14] ;
 wire \tholin_riscv.uart.receive_div_counter[15] ;
 wire \tholin_riscv.uart.receive_div_counter[1] ;
 wire \tholin_riscv.uart.receive_div_counter[2] ;
 wire \tholin_riscv.uart.receive_div_counter[3] ;
 wire \tholin_riscv.uart.receive_div_counter[4] ;
 wire \tholin_riscv.uart.receive_div_counter[5] ;
 wire \tholin_riscv.uart.receive_div_counter[6] ;
 wire \tholin_riscv.uart.receive_div_counter[7] ;
 wire \tholin_riscv.uart.receive_div_counter[8] ;
 wire \tholin_riscv.uart.receive_div_counter[9] ;
 wire \tholin_riscv.uart.receiving ;
 wire \tholin_riscv.uart_int_enable ;

 sky130_as_sc_hs__diode_2 ANTENNA_1 (.DIODE(wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA__26229__A (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__26229__B (.DIODE(_19755_));
 sky130_as_sc_hs__diode_2 ANTENNA__26239__B (.DIODE(_19764_));
 sky130_as_sc_hs__diode_2 ANTENNA__26241__B (.DIODE(_19764_));
 sky130_as_sc_hs__diode_2 ANTENNA__26243__A (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__26244__A (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__26249__A (.DIODE(clknet_4_0__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA__26256__A (.DIODE(_19754_));
 sky130_as_sc_hs__diode_2 ANTENNA__26259__A (.DIODE(_19761_));
 sky130_as_sc_hs__diode_2 ANTENNA__26264__A (.DIODE(\tholin_riscv.requested_addr[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26269__A (.DIODE(_19784_));
 sky130_as_sc_hs__diode_2 ANTENNA__26271__A (.DIODE(\tholin_riscv.requested_addr[3] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26275__A (.DIODE(_19790_));
 sky130_as_sc_hs__diode_2 ANTENNA__26277__A (.DIODE(\tholin_riscv.requested_addr[4] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26281__A (.DIODE(_19795_));
 sky130_as_sc_hs__diode_2 ANTENNA__26283__A (.DIODE(\tholin_riscv.requested_addr[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26287__A (.DIODE(_19800_));
 sky130_as_sc_hs__diode_2 ANTENNA__26289__A (.DIODE(\tholin_riscv.requested_addr[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26293__A (.DIODE(_19805_));
 sky130_as_sc_hs__diode_2 ANTENNA__26295__A (.DIODE(\tholin_riscv.requested_addr[7] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26299__A (.DIODE(_19810_));
 sky130_as_sc_hs__diode_2 ANTENNA__26305__A (.DIODE(_19815_));
 sky130_as_sc_hs__diode_2 ANTENNA__26306__A (.DIODE(\tholin_riscv.Bimm[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26307__A (.DIODE(\tholin_riscv.instr[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26315__A (.DIODE(\tholin_riscv.Bimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26316__A (.DIODE(\tholin_riscv.instr[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26324__A (.DIODE(\tholin_riscv.Bimm[3] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26333__A (.DIODE(\tholin_riscv.Bimm[4] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26342__A (.DIODE(\tholin_riscv.Jimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26351__A (.DIODE(\tholin_riscv.Jimm[13] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26360__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__26369__A (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA__26370__A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26397__A (.DIODE(\tholin_riscv.requested_addr[7] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26397__B (.DIODE(\tholin_riscv.requested_addr[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26398__A (.DIODE(\tholin_riscv.requested_addr[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26398__B (.DIODE(\tholin_riscv.requested_addr[4] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26401__A (.DIODE(\tholin_riscv.requested_addr[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26403__B (.DIODE(\tholin_riscv.requested_addr[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26405__B (.DIODE(\tholin_riscv.requested_addr[4] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26407__A (.DIODE(\tholin_riscv.requested_addr[3] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26411__A (.DIODE(\tholin_riscv.requested_addr[3] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26411__B (.DIODE(\tholin_riscv.requested_addr[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26413__B (.DIODE(\tholin_riscv.requested_addr[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26414__A (.DIODE(\tholin_riscv.requested_addr[3] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26414__B (.DIODE(\tholin_riscv.requested_addr[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26418__B (.DIODE(_19920_));
 sky130_as_sc_hs__diode_2 ANTENNA__26438__B (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__26441__A (.DIODE(\tholin_riscv.instr[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26441__B (.DIODE(\tholin_riscv.instr[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26446__A (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__26446__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__26447__A (.DIODE(\tholin_riscv.requested_addr[4] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26458__C (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__26476__A (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__26476__B (.DIODE(\tholin_riscv.Bimm[10] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26477__A (.DIODE(\tholin_riscv.Bimm[9] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26479__B (.DIODE(\tholin_riscv.Bimm[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26480__A (.DIODE(\tholin_riscv.Bimm[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__26490__B (.DIODE(_19764_));
 sky130_as_sc_hs__diode_2 ANTENNA__26492__A (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__26493__A (.DIODE(_19920_));
 sky130_as_sc_hs__diode_2 ANTENNA__26493__B (.DIODE(_19993_));
 sky130_as_sc_hs__diode_2 ANTENNA__26502__C (.DIODE(_19993_));
 sky130_as_sc_hs__diode_2 ANTENNA__26503__A (.DIODE(_20005_));
 sky130_as_sc_hs__diode_2 ANTENNA__26505__A (.DIODE(net145));
 sky130_as_sc_hs__diode_2 ANTENNA__26509__A (.DIODE(_19761_));
 sky130_as_sc_hs__diode_2 ANTENNA__26531__A (.DIODE(_19920_));
 sky130_as_sc_hs__diode_2 ANTENNA__26538__A (.DIODE(_19534_));
 sky130_as_sc_hs__diode_2 ANTENNA__26540__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__26541__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26544__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__26545__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26548__A (.DIODE(_19534_));
 sky130_as_sc_hs__diode_2 ANTENNA__26550__A (.DIODE(net281));
 sky130_as_sc_hs__diode_2 ANTENNA__26551__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__26552__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26555__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__26557__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__26558__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__26559__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__26561__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__26562__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__26564__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__26565__A (.DIODE(net262));
 sky130_as_sc_hs__diode_2 ANTENNA__26566__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__26567__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__26568__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__26569__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26570__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__26571__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__26572__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26573__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__26574__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__26575__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__26576__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26578__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__26579__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26581__A (.DIODE(net281));
 sky130_as_sc_hs__diode_2 ANTENNA__26582__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__26583__A (.DIODE(net198));
 sky130_as_sc_hs__diode_2 ANTENNA__26584__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__26585__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__26586__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26587__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__26588__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__26589__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__26590__A (.DIODE(net198));
 sky130_as_sc_hs__diode_2 ANTENNA__26592__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__26593__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__26595__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__26596__A (.DIODE(net262));
 sky130_as_sc_hs__diode_2 ANTENNA__26597__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__26598__A (.DIODE(net253));
 sky130_as_sc_hs__diode_2 ANTENNA__26599__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__26603__A (.DIODE(net20));
 sky130_as_sc_hs__diode_2 ANTENNA__26603__B (.DIODE(_19755_));
 sky130_as_sc_hs__diode_2 ANTENNA__26604__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__26605__A (.DIODE(net1710));
 sky130_as_sc_hs__diode_2 ANTENNA__26605__B (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__26606__A (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__26625__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__26628__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__26629__A (.DIODE(net333));
 sky130_as_sc_hs__diode_2 ANTENNA__26630__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__26631__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__26632__A (.DIODE(net198));
 sky130_as_sc_hs__diode_2 ANTENNA__26634__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__26635__A (.DIODE(net198));
 sky130_as_sc_hs__diode_2 ANTENNA__26637__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__26638__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__26639__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__26642__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__26643__A (.DIODE(net320));
 sky130_as_sc_hs__diode_2 ANTENNA__26645__A (.DIODE(net160));
 sky130_as_sc_hs__diode_2 ANTENNA__26646__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__26647__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__26648__A (.DIODE(net274));
 sky130_as_sc_hs__diode_2 ANTENNA__26649__A (.DIODE(net198));
 sky130_as_sc_hs__diode_2 ANTENNA__26651__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__26652__A (.DIODE(net259));
 sky130_as_sc_hs__diode_2 ANTENNA__26653__A (.DIODE(net153));
 sky130_as_sc_hs__diode_2 ANTENNA__26654__A (.DIODE(net250));
 sky130_as_sc_hs__diode_2 ANTENNA__26655__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__26656__A (.DIODE(net198));
 sky130_as_sc_hs__diode_2 ANTENNA__26657__A (.DIODE(net333));
 sky130_as_sc_hs__diode_2 ANTENNA__26658__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__26659__A (.DIODE(net198));
 sky130_as_sc_hs__diode_2 ANTENNA__26661__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__26662__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__26663__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26664__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__26665__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__26666__A (.DIODE(net198));
 sky130_as_sc_hs__diode_2 ANTENNA__26667__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__26668__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__26669__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__26670__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26671__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__26672__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__26673__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26674__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__26675__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__26676__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__26677__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26678__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__26679__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__26680__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26681__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__26682__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__26683__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__26684__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__26685__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__26686__A (.DIODE(_19538_));
 sky130_as_sc_hs__diode_2 ANTENNA__26690__A (.DIODE(net21));
 sky130_as_sc_hs__diode_2 ANTENNA__26690__B (.DIODE(_19755_));
 sky130_as_sc_hs__diode_2 ANTENNA__26691__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__26692__A (.DIODE(net1780));
 sky130_as_sc_hs__diode_2 ANTENNA__26692__B (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__26693__A (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__26712__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__26715__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__26716__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__26717__A (.DIODE(net274));
 sky130_as_sc_hs__diode_2 ANTENNA__26718__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__26719__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__26722__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__26723__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__26724__A (.DIODE(net274));
 sky130_as_sc_hs__diode_2 ANTENNA__26725__A (.DIODE(net259));
 sky130_as_sc_hs__diode_2 ANTENNA__26726__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__26729__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__26731__A (.DIODE(net274));
 sky130_as_sc_hs__diode_2 ANTENNA__26732__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__26733__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__26734__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__26735__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__26736__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__26737__A (.DIODE(net333));
 sky130_as_sc_hs__diode_2 ANTENNA__26738__A (.DIODE(net175));
 sky130_as_sc_hs__diode_2 ANTENNA__26739__A (.DIODE(net259));
 sky130_as_sc_hs__diode_2 ANTENNA__26740__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__26741__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__26742__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__26744__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__26745__A (.DIODE(net175));
 sky130_as_sc_hs__diode_2 ANTENNA__26747__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__26748__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__26749__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__26751__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__26752__A (.DIODE(net175));
 sky130_as_sc_hs__diode_2 ANTENNA__26753__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__26754__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__26755__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__26756__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__26757__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__26759__A (.DIODE(net175));
 sky130_as_sc_hs__diode_2 ANTENNA__26760__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__26761__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__26762__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__26763__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__26765__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__26766__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__26767__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__26768__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__26769__A (.DIODE(net175));
 sky130_as_sc_hs__diode_2 ANTENNA__26770__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__26771__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__26772__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__26773__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__26776__A (.DIODE(net4));
 sky130_as_sc_hs__diode_2 ANTENNA__26776__B (.DIODE(_19755_));
 sky130_as_sc_hs__diode_2 ANTENNA__26777__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__26778__A (.DIODE(net1791));
 sky130_as_sc_hs__diode_2 ANTENNA__26778__B (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__26779__A (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__26793__A (.DIODE(_19993_));
 sky130_as_sc_hs__diode_2 ANTENNA__26798__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__26799__A (.DIODE(net190));
 sky130_as_sc_hs__diode_2 ANTENNA__26801__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__26802__A (.DIODE(net190));
 sky130_as_sc_hs__diode_2 ANTENNA__26804__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__26805__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__26806__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__26808__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__26809__A (.DIODE(net195));
 sky130_as_sc_hs__diode_2 ANTENNA__26811__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__26812__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__26813__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__26814__A (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__26815__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__26816__A (.DIODE(net190));
 sky130_as_sc_hs__diode_2 ANTENNA__26818__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__26819__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__26820__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__26821__A (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__26822__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__26823__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__26825__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__26826__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__26827__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__26828__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__26829__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__26831__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__26832__A (.DIODE(net175));
 sky130_as_sc_hs__diode_2 ANTENNA__26833__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__26834__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__26835__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__26836__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__26837__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__26838__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__26839__A (.DIODE(net175));
 sky130_as_sc_hs__diode_2 ANTENNA__26841__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__26842__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__26843__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__26846__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__26847__A (.DIODE(net190));
 sky130_as_sc_hs__diode_2 ANTENNA__26849__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__26850__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__26851__A (.DIODE(net190));
 sky130_as_sc_hs__diode_2 ANTENNA__26853__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__26854__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__26856__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__26857__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__26858__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__26859__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__26860__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__26864__A (.DIODE(net5));
 sky130_as_sc_hs__diode_2 ANTENNA__26864__B (.DIODE(_19755_));
 sky130_as_sc_hs__diode_2 ANTENNA__26865__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__26866__A (.DIODE(net1792));
 sky130_as_sc_hs__diode_2 ANTENNA__26866__B (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__26867__A (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__26868__A (.DIODE(net502));
 sky130_as_sc_hs__diode_2 ANTENNA__26888__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__26891__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__26892__A (.DIODE(net160));
 sky130_as_sc_hs__diode_2 ANTENNA__26895__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__26898__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__26899__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__26902__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__26905__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__26906__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__26909__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__26912__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__26913__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__26914__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__26915__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__26916__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__26922__A (.DIODE(net274));
 sky130_as_sc_hs__diode_2 ANTENNA__26923__A (.DIODE(net160));
 sky130_as_sc_hs__diode_2 ANTENNA__26926__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__26929__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__26930__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__26931__B (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__26932__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__26934__B (.DIODE(net320));
 sky130_as_sc_hs__diode_2 ANTENNA__26937__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__26940__A (.DIODE(net274));
 sky130_as_sc_hs__diode_2 ANTENNA__26944__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__26945__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__26946__A (.DIODE(net250));
 sky130_as_sc_hs__diode_2 ANTENNA__26947__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__26950__A (.DIODE(net6));
 sky130_as_sc_hs__diode_2 ANTENNA__26950__B (.DIODE(_19755_));
 sky130_as_sc_hs__diode_2 ANTENNA__26951__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__26952__B (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__26953__A (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__26967__A (.DIODE(_19920_));
 sky130_as_sc_hs__diode_2 ANTENNA__26975__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__26978__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__26979__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__26982__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__26985__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__26986__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__26987__B (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__26988__A (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__26989__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__26990__B (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__26991__A (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__26992__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__26993__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__26994__B (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__26995__A (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__26996__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__26997__B (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__26998__A (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__26999__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__27000__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__27001__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__27002__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__27003__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__27006__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__27009__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__27010__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__27013__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__27016__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__27017__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__27020__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__27023__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__27024__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__27027__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__27030__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__27031__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__27032__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__27033__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__27034__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__27038__A (.DIODE(net7));
 sky130_as_sc_hs__diode_2 ANTENNA__27038__B (.DIODE(_19755_));
 sky130_as_sc_hs__diode_2 ANTENNA__27039__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__27040__B (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__27041__A (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__27055__A (.DIODE(_19993_));
 sky130_as_sc_hs__diode_2 ANTENNA__27063__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27066__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27067__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__27070__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27073__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27074__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__27077__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27080__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27081__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__27084__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27087__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27088__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__27089__A (.DIODE(net153));
 sky130_as_sc_hs__diode_2 ANTENNA__27090__A (.DIODE(net250));
 sky130_as_sc_hs__diode_2 ANTENNA__27091__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__27094__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27097__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27098__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__27101__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27104__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27105__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__27108__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27109__B (.DIODE(net292));
 sky130_as_sc_hs__diode_2 ANTENNA__27110__A (.DIODE(net292));
 sky130_as_sc_hs__diode_2 ANTENNA__27111__A (.DIODE(net282));
 sky130_as_sc_hs__diode_2 ANTENNA__27112__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__27115__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27116__B (.DIODE(net292));
 sky130_as_sc_hs__diode_2 ANTENNA__27117__A (.DIODE(net292));
 sky130_as_sc_hs__diode_2 ANTENNA__27118__A (.DIODE(net173));
 sky130_as_sc_hs__diode_2 ANTENNA__27119__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__27120__A (.DIODE(net153));
 sky130_as_sc_hs__diode_2 ANTENNA__27121__A (.DIODE(net250));
 sky130_as_sc_hs__diode_2 ANTENNA__27122__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__27124__A (.DIODE(_19754_));
 sky130_as_sc_hs__diode_2 ANTENNA__27124__B (.DIODE(_20622_));
 sky130_as_sc_hs__diode_2 ANTENNA__27125__A (.DIODE(net8));
 sky130_as_sc_hs__diode_2 ANTENNA__27125__B (.DIODE(_19755_));
 sky130_as_sc_hs__diode_2 ANTENNA__27126__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__27127__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__27127__B (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__27128__A (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__27149__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27152__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27153__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__27156__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27159__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27160__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__27163__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27166__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27167__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__27170__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27173__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27174__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__27175__A (.DIODE(net153));
 sky130_as_sc_hs__diode_2 ANTENNA__27176__A (.DIODE(net250));
 sky130_as_sc_hs__diode_2 ANTENNA__27177__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__27178__B (.DIODE(net291));
 sky130_as_sc_hs__diode_2 ANTENNA__27180__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27183__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27184__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__27187__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27190__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__27191__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__27194__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__27197__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27198__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__27201__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__27204__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27205__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__27206__A (.DIODE(net153));
 sky130_as_sc_hs__diode_2 ANTENNA__27207__A (.DIODE(net250));
 sky130_as_sc_hs__diode_2 ANTENNA__27208__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__27210__A (.DIODE(_19754_));
 sky130_as_sc_hs__diode_2 ANTENNA__27210__B (.DIODE(_20707_));
 sky130_as_sc_hs__diode_2 ANTENNA__27211__A (.DIODE(net9));
 sky130_as_sc_hs__diode_2 ANTENNA__27211__B (.DIODE(_19755_));
 sky130_as_sc_hs__diode_2 ANTENNA__27212__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__27213__A (.DIODE(net373));
 sky130_as_sc_hs__diode_2 ANTENNA__27213__B (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__27214__A (.DIODE(_20021_));
 sky130_as_sc_hs__diode_2 ANTENNA__27257__A (.DIODE(_19993_));
 sky130_as_sc_hs__diode_2 ANTENNA__27265__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__27268__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__27271__A (.DIODE(net266));
 sky130_as_sc_hs__diode_2 ANTENNA__27272__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__27275__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__27278__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__27279__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__27282__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__27285__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__27286__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__27289__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__27292__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__27293__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__27294__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__27295__A (.DIODE(net253));
 sky130_as_sc_hs__diode_2 ANTENNA__27296__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__27299__A (.DIODE(net169));
 sky130_as_sc_hs__diode_2 ANTENNA__27302__A (.DIODE(net266));
 sky130_as_sc_hs__diode_2 ANTENNA__27303__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__27306__A (.DIODE(net169));
 sky130_as_sc_hs__diode_2 ANTENNA__27309__A (.DIODE(net266));
 sky130_as_sc_hs__diode_2 ANTENNA__27310__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__27313__A (.DIODE(net169));
 sky130_as_sc_hs__diode_2 ANTENNA__27315__A (.DIODE(net307));
 sky130_as_sc_hs__diode_2 ANTENNA__27316__A (.DIODE(net266));
 sky130_as_sc_hs__diode_2 ANTENNA__27317__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__27319__A (.DIODE(net307));
 sky130_as_sc_hs__diode_2 ANTENNA__27320__A (.DIODE(net266));
 sky130_as_sc_hs__diode_2 ANTENNA__27322__A (.DIODE(net307));
 sky130_as_sc_hs__diode_2 ANTENNA__27323__A (.DIODE(net169));
 sky130_as_sc_hs__diode_2 ANTENNA__27324__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__27325__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__27326__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__27327__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__27333__A (.DIODE(_19754_));
 sky130_as_sc_hs__diode_2 ANTENNA__27334__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__27336__A (.DIODE(\tholin_riscv.instr[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__27337__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__27364__A (.DIODE(_19993_));
 sky130_as_sc_hs__diode_2 ANTENNA__27375__A (.DIODE(net169));
 sky130_as_sc_hs__diode_2 ANTENNA__27378__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__27379__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__27382__A (.DIODE(net169));
 sky130_as_sc_hs__diode_2 ANTENNA__27385__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__27386__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__27389__A (.DIODE(net169));
 sky130_as_sc_hs__diode_2 ANTENNA__27392__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__27393__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__27396__A (.DIODE(net266));
 sky130_as_sc_hs__diode_2 ANTENNA__27399__A (.DIODE(net169));
 sky130_as_sc_hs__diode_2 ANTENNA__27400__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__27401__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__27402__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__27403__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__27406__A (.DIODE(net169));
 sky130_as_sc_hs__diode_2 ANTENNA__27409__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__27410__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__27413__A (.DIODE(net169));
 sky130_as_sc_hs__diode_2 ANTENNA__27416__A (.DIODE(net266));
 sky130_as_sc_hs__diode_2 ANTENNA__27417__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__27420__A (.DIODE(net169));
 sky130_as_sc_hs__diode_2 ANTENNA__27423__A (.DIODE(net266));
 sky130_as_sc_hs__diode_2 ANTENNA__27424__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__27427__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__27430__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__27431__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__27432__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__27433__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__27434__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__27440__A (.DIODE(_19754_));
 sky130_as_sc_hs__diode_2 ANTENNA__27441__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__27443__A (.DIODE(net1684));
 sky130_as_sc_hs__diode_2 ANTENNA__27444__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__27479__B (.DIODE(net292));
 sky130_as_sc_hs__diode_2 ANTENNA__27480__A (.DIODE(net292));
 sky130_as_sc_hs__diode_2 ANTENNA__27481__A (.DIODE(net173));
 sky130_as_sc_hs__diode_2 ANTENNA__27484__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__27485__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__27488__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__27491__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__27492__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__27493__B (.DIODE(net292));
 sky130_as_sc_hs__diode_2 ANTENNA__27494__A (.DIODE(net292));
 sky130_as_sc_hs__diode_2 ANTENNA__27495__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__27498__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__27499__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__27502__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__27505__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__27506__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__27507__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__27508__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__27509__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__27512__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__27515__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__27516__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__27519__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__27522__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__27523__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__27526__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__27529__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__27530__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__27533__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__27536__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__27537__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__27538__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__27539__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__27540__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__27546__A (.DIODE(_19754_));
 sky130_as_sc_hs__diode_2 ANTENNA__27547__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__27550__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__27581__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__27584__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27587__A (.DIODE(net264));
 sky130_as_sc_hs__diode_2 ANTENNA__27588__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__27591__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27594__A (.DIODE(net264));
 sky130_as_sc_hs__diode_2 ANTENNA__27595__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__27598__A (.DIODE(net173));
 sky130_as_sc_hs__diode_2 ANTENNA__27601__A (.DIODE(net264));
 sky130_as_sc_hs__diode_2 ANTENNA__27602__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__27603__B (.DIODE(net292));
 sky130_as_sc_hs__diode_2 ANTENNA__27604__A (.DIODE(net292));
 sky130_as_sc_hs__diode_2 ANTENNA__27605__A (.DIODE(net282));
 sky130_as_sc_hs__diode_2 ANTENNA__27606__B (.DIODE(net292));
 sky130_as_sc_hs__diode_2 ANTENNA__27607__A (.DIODE(net292));
 sky130_as_sc_hs__diode_2 ANTENNA__27608__A (.DIODE(net173));
 sky130_as_sc_hs__diode_2 ANTENNA__27609__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__27610__A (.DIODE(net153));
 sky130_as_sc_hs__diode_2 ANTENNA__27611__A (.DIODE(net250));
 sky130_as_sc_hs__diode_2 ANTENNA__27613__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__27616__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27619__A (.DIODE(net264));
 sky130_as_sc_hs__diode_2 ANTENNA__27620__A (.DIODE(net160));
 sky130_as_sc_hs__diode_2 ANTENNA__27623__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27626__A (.DIODE(net264));
 sky130_as_sc_hs__diode_2 ANTENNA__27627__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__27630__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27633__A (.DIODE(net264));
 sky130_as_sc_hs__diode_2 ANTENNA__27634__A (.DIODE(net160));
 sky130_as_sc_hs__diode_2 ANTENNA__27637__A (.DIODE(net264));
 sky130_as_sc_hs__diode_2 ANTENNA__27640__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27641__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__27642__A (.DIODE(net153));
 sky130_as_sc_hs__diode_2 ANTENNA__27643__A (.DIODE(net250));
 sky130_as_sc_hs__diode_2 ANTENNA__27645__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__27651__A (.DIODE(_19754_));
 sky130_as_sc_hs__diode_2 ANTENNA__27652__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__27655__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__27678__A (.DIODE(_19920_));
 sky130_as_sc_hs__diode_2 ANTENNA__27686__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__27689__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27692__A (.DIODE(net269));
 sky130_as_sc_hs__diode_2 ANTENNA__27693__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__27696__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27699__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__27700__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__27703__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27706__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__27707__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__27710__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__27713__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27714__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__27715__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__27716__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__27717__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__27720__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27723__A (.DIODE(net269));
 sky130_as_sc_hs__diode_2 ANTENNA__27724__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__27727__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27730__A (.DIODE(net269));
 sky130_as_sc_hs__diode_2 ANTENNA__27731__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__27734__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27737__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__27738__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__27741__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__27744__A (.DIODE(net172));
 sky130_as_sc_hs__diode_2 ANTENNA__27745__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__27746__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__27747__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__27748__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__27753__A (.DIODE(_19754_));
 sky130_as_sc_hs__diode_2 ANTENNA__27754__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__27757__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__27791__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27794__A (.DIODE(net264));
 sky130_as_sc_hs__diode_2 ANTENNA__27795__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__27798__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27801__A (.DIODE(net264));
 sky130_as_sc_hs__diode_2 ANTENNA__27802__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__27805__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27808__A (.DIODE(net264));
 sky130_as_sc_hs__diode_2 ANTENNA__27809__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__27812__A (.DIODE(net264));
 sky130_as_sc_hs__diode_2 ANTENNA__27815__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27816__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__27817__A (.DIODE(net153));
 sky130_as_sc_hs__diode_2 ANTENNA__27818__A (.DIODE(net250));
 sky130_as_sc_hs__diode_2 ANTENNA__27819__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__27822__A (.DIODE(net172));
 sky130_as_sc_hs__diode_2 ANTENNA__27825__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__27826__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__27829__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__27832__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__27833__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__27836__A (.DIODE(net172));
 sky130_as_sc_hs__diode_2 ANTENNA__27839__A (.DIODE(net269));
 sky130_as_sc_hs__diode_2 ANTENNA__27840__A (.DIODE(net165));
 sky130_as_sc_hs__diode_2 ANTENNA__27843__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__27846__A (.DIODE(net175));
 sky130_as_sc_hs__diode_2 ANTENNA__27847__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__27848__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__27849__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__27850__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__27856__A (.DIODE(_19754_));
 sky130_as_sc_hs__diode_2 ANTENNA__27857__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__27860__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__27889__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27892__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__27893__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__27896__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27899__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__27900__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__27903__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27906__A (.DIODE(net264));
 sky130_as_sc_hs__diode_2 ANTENNA__27907__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__27910__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__27913__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27914__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__27915__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__27916__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__27917__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__27920__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27923__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__27924__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__27927__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27930__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__27931__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__27934__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27937__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__27938__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__27941__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__27944__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__27945__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__27946__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__27947__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__27948__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__27950__A (.DIODE(_19754_));
 sky130_as_sc_hs__diode_2 ANTENNA__27950__B (.DIODE(_21440_));
 sky130_as_sc_hs__diode_2 ANTENNA__27953__A (.DIODE(_19754_));
 sky130_as_sc_hs__diode_2 ANTENNA__27954__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__27957__A (.DIODE(net502));
 sky130_as_sc_hs__diode_2 ANTENNA__27982__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__27984__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27985__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__27987__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__27988__A (.DIODE(net160));
 sky130_as_sc_hs__diode_2 ANTENNA__27989__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__27990__A (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__27991__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__27992__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__27994__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__27995__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__27996__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__27998__A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA__27999__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__28001__A (.DIODE(net264));
 sky130_as_sc_hs__diode_2 ANTENNA__28002__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__28003__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__28005__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__28006__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__28008__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__28009__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__28010__A (.DIODE(net153));
 sky130_as_sc_hs__diode_2 ANTENNA__28011__A (.DIODE(net250));
 sky130_as_sc_hs__diode_2 ANTENNA__28012__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__28013__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__28015__A (.DIODE(net175));
 sky130_as_sc_hs__diode_2 ANTENNA__28016__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__28017__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__28018__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__28019__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__28021__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__28022__A (.DIODE(net175));
 sky130_as_sc_hs__diode_2 ANTENNA__28023__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__28025__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__28026__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__28027__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__28029__A (.DIODE(net175));
 sky130_as_sc_hs__diode_2 ANTENNA__28030__A (.DIODE(net188));
 sky130_as_sc_hs__diode_2 ANTENNA__28032__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__28033__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__28035__A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA__28036__A (.DIODE(net271));
 sky130_as_sc_hs__diode_2 ANTENNA__28039__A (.DIODE(net175));
 sky130_as_sc_hs__diode_2 ANTENNA__28040__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__28041__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__28042__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__28043__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__28049__A (.DIODE(_19754_));
 sky130_as_sc_hs__diode_2 ANTENNA__28050__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__28052__A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA__28053__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__28055__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__28058__B (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__28059__A (.DIODE(\tholin_riscv.Bimm[4] ));
 sky130_as_sc_hs__diode_2 ANTENNA__28062__B (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__28063__A (.DIODE(\tholin_riscv.Bimm[3] ));
 sky130_as_sc_hs__diode_2 ANTENNA__28067__B (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__28068__A (.DIODE(\tholin_riscv.Bimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__28077__A (.DIODE(net145));
 sky130_as_sc_hs__diode_2 ANTENNA__28081__A (.DIODE(net502));
 sky130_as_sc_hs__diode_2 ANTENNA__28081__B (.DIODE(net145));
 sky130_as_sc_hs__diode_2 ANTENNA__28086__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__28087__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__28088__B (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__28089__A (.DIODE(\tholin_riscv.Bimm[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__28091__B (.DIODE(_21576_));
 sky130_as_sc_hs__diode_2 ANTENNA__28092__B (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__28093__A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA__28099__A (.DIODE(\tholin_riscv.instr[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__28099__B (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__28109__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28110__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__28116__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28117__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__28124__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__28131__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__28132__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__28133__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__28134__A (.DIODE(\tholin_riscv.Jimm[19] ));
 sky130_as_sc_hs__diode_2 ANTENNA__28140__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28141__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__28147__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28148__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__28154__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28155__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__28162__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__28163__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__28164__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__28165__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__28167__A (.DIODE(\tholin_riscv.Jimm[13] ));
 sky130_as_sc_hs__diode_2 ANTENNA__28167__B (.DIODE(\tholin_riscv.Jimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__28169__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__28170__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__28174__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__28177__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__28178__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__28181__A (.DIODE(net224));
 sky130_as_sc_hs__diode_2 ANTENNA__28184__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__28185__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__28188__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__28191__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__28192__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__28195__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__28198__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__28199__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__28200__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__28201__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__28202__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__28208__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28209__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__28215__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28216__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__28222__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28223__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__28230__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__28231__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__28232__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__28233__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__28235__A (.DIODE(net400));
 sky130_as_sc_hs__diode_2 ANTENNA__28237__A (.DIODE(net224));
 sky130_as_sc_hs__diode_2 ANTENNA__28238__A (.DIODE(net400));
 sky130_as_sc_hs__diode_2 ANTENNA__28241__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__28242__A (.DIODE(net400));
 sky130_as_sc_hs__diode_2 ANTENNA__28244__A (.DIODE(net224));
 sky130_as_sc_hs__diode_2 ANTENNA__28245__A (.DIODE(net400));
 sky130_as_sc_hs__diode_2 ANTENNA__28248__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__28251__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__28255__A (.DIODE(net239));
 sky130_as_sc_hs__diode_2 ANTENNA__28261__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__28262__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__28263__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__28264__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__28265__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__28269__A (.DIODE(net409));
 sky130_as_sc_hs__diode_2 ANTENNA__28271__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28272__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__28273__A (.DIODE(net409));
 sky130_as_sc_hs__diode_2 ANTENNA__28276__A (.DIODE(net409));
 sky130_as_sc_hs__diode_2 ANTENNA__28278__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28279__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__28285__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28286__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__28289__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__28293__A (.DIODE(net350));
 sky130_as_sc_hs__diode_2 ANTENNA__28294__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__28295__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__28296__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__28301__A (.DIODE(net230));
 sky130_as_sc_hs__diode_2 ANTENNA__28304__A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA__28305__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__28308__A (.DIODE(net230));
 sky130_as_sc_hs__diode_2 ANTENNA__28311__A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA__28312__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__28315__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__28318__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__28319__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__28322__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__28325__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__28326__A (.DIODE(net350));
 sky130_as_sc_hs__diode_2 ANTENNA__28327__A (.DIODE(net244));
 sky130_as_sc_hs__diode_2 ANTENNA__28328__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__28329__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__28332__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__28335__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__28336__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__28339__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__28342__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__28343__A (.DIODE(net350));
 sky130_as_sc_hs__diode_2 ANTENNA__28346__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__28349__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__28350__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__28353__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__28356__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__28357__A (.DIODE(net350));
 sky130_as_sc_hs__diode_2 ANTENNA__28358__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__28359__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__28360__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__28365__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28368__A (.DIODE(net358));
 sky130_as_sc_hs__diode_2 ANTENNA__28369__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__28372__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__28375__A (.DIODE(net358));
 sky130_as_sc_hs__diode_2 ANTENNA__28376__A (.DIODE(net345));
 sky130_as_sc_hs__diode_2 ANTENNA__28379__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28382__A (.DIODE(net358));
 sky130_as_sc_hs__diode_2 ANTENNA__28383__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__28386__A (.DIODE(net358));
 sky130_as_sc_hs__diode_2 ANTENNA__28389__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__28390__A (.DIODE(net345));
 sky130_as_sc_hs__diode_2 ANTENNA__28391__A (.DIODE(net241));
 sky130_as_sc_hs__diode_2 ANTENNA__28392__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__28393__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__28394__A (.DIODE(net409));
 sky130_as_sc_hs__diode_2 ANTENNA__28397__A (.DIODE(net409));
 sky130_as_sc_hs__diode_2 ANTENNA__28399__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28400__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__28402__A (.DIODE(net209));
 sky130_as_sc_hs__diode_2 ANTENNA__28403__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28404__A (.DIODE(net410));
 sky130_as_sc_hs__diode_2 ANTENNA__28406__A (.DIODE(net358));
 sky130_as_sc_hs__diode_2 ANTENNA__28407__A (.DIODE(net345));
 sky130_as_sc_hs__diode_2 ANTENNA__28408__A (.DIODE(net410));
 sky130_as_sc_hs__diode_2 ANTENNA__28410__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28413__A (.DIODE(net358));
 sky130_as_sc_hs__diode_2 ANTENNA__28414__A (.DIODE(net234));
 sky130_as_sc_hs__diode_2 ANTENNA__28417__A (.DIODE(net358));
 sky130_as_sc_hs__diode_2 ANTENNA__28420__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28421__A (.DIODE(net345));
 sky130_as_sc_hs__diode_2 ANTENNA__28422__A (.DIODE(net241));
 sky130_as_sc_hs__diode_2 ANTENNA__28423__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__28424__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__28426__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__28427__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28428__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__28429__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__28430__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28431__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__28432__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__28434__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28435__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__28436__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__28437__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28438__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__28439__A (.DIODE(net343));
 sky130_as_sc_hs__diode_2 ANTENNA__28440__A (.DIODE(net373));
 sky130_as_sc_hs__diode_2 ANTENNA__28441__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__28442__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__28443__A (.DIODE(net373));
 sky130_as_sc_hs__diode_2 ANTENNA__28444__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__28445__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__28446__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__28447__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__28448__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__28449__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__28450__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__28451__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28452__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__28453__A (.DIODE(net343));
 sky130_as_sc_hs__diode_2 ANTENNA__28454__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__28455__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__28456__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__28458__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28459__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__28461__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28462__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__28463__A (.DIODE(_19483_));
 sky130_as_sc_hs__diode_2 ANTENNA__28465__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28466__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__28468__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28469__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__28470__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__28473__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__28476__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__28477__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__28479__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__28480__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__28482__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__28483__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__28484__A (.DIODE(net343));
 sky130_as_sc_hs__diode_2 ANTENNA__28485__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__28486__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__28487__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__28489__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__28490__B (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__28491__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__28492__A (.DIODE(net373));
 sky130_as_sc_hs__diode_2 ANTENNA__28493__B (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28494__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__28495__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__28496__A (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28497__B (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28498__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__28499__A (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28500__B (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28501__A (.DIODE(net361));
 sky130_as_sc_hs__diode_2 ANTENNA__28502__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__28503__A (.DIODE(net373));
 sky130_as_sc_hs__diode_2 ANTENNA__28504__B (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__28505__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__28506__A (.DIODE(net373));
 sky130_as_sc_hs__diode_2 ANTENNA__28507__B (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28508__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__28509__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__28512__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__28515__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__28516__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__28517__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__28518__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__28519__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__28520__A (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28522__A (.DIODE(net224));
 sky130_as_sc_hs__diode_2 ANTENNA__28525__A (.DIODE(net361));
 sky130_as_sc_hs__diode_2 ANTENNA__28526__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__28527__A (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28528__B (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28529__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__28530__A (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28531__B (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28532__A (.DIODE(net361));
 sky130_as_sc_hs__diode_2 ANTENNA__28533__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__28536__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__28539__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__28540__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__28541__A (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28542__B (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28543__A (.DIODE(net361));
 sky130_as_sc_hs__diode_2 ANTENNA__28546__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__28547__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__28548__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__28549__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__28550__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__28555__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__28558__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__28559__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__28562__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__28565__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__28566__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__28569__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__28572__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__28573__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__28576__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__28579__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__28580__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__28581__A (.DIODE(net244));
 sky130_as_sc_hs__diode_2 ANTENNA__28582__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__28583__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__28585__B (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA__28586__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__28589__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__28590__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__28593__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__28596__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__28597__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__28600__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__28603__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__28604__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__28607__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__28610__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__28611__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__28612__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__28613__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__28614__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__28618__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__28621__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__28622__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__28625__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__28626__A (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA__28627__B (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA__28628__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__28629__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__28632__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__28635__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__28636__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__28637__A (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA__28638__B (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA__28639__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__28642__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__28643__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__28644__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__28645__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__28646__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__28649__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__28652__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__28653__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__28656__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__28657__A (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA__28658__B (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA__28659__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__28660__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__28663__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__28666__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__28667__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__28668__A (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA__28669__B (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA__28670__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__28673__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__28674__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__28675__A (.DIODE(net244));
 sky130_as_sc_hs__diode_2 ANTENNA__28676__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__28677__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__28682__A (.DIODE(_21977_));
 sky130_as_sc_hs__diode_2 ANTENNA__28685__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__28688__A (.DIODE(net361));
 sky130_as_sc_hs__diode_2 ANTENNA__28689__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__28692__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__28693__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__28695__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__28696__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__28699__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__28702__A (.DIODE(net361));
 sky130_as_sc_hs__diode_2 ANTENNA__28703__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__28706__A (.DIODE(net361));
 sky130_as_sc_hs__diode_2 ANTENNA__28707__A (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28709__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__28710__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__28711__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__28712__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__28713__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__28714__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__28716__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__28717__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__28720__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__28721__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__28724__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__28727__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__28728__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__28731__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__28734__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__28735__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__28738__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__28740__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__28741__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__28742__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__28743__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__28744__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__28751__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__28752__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28754__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__28755__A (.DIODE(net358));
 sky130_as_sc_hs__diode_2 ANTENNA__28756__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__28757__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__28758__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__28759__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__28761__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__28762__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__28763__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__28764__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__28765__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__28766__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__28768__A (.DIODE(net210));
 sky130_as_sc_hs__diode_2 ANTENNA__28769__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__28770__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__28771__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__28772__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__28773__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__28774__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__28775__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__28776__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__28777__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__28778__A (.DIODE(net241));
 sky130_as_sc_hs__diode_2 ANTENNA__28779__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__28780__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__28782__A (.DIODE(net209));
 sky130_as_sc_hs__diode_2 ANTENNA__28783__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28786__A (.DIODE(net358));
 sky130_as_sc_hs__diode_2 ANTENNA__28787__A (.DIODE(net234));
 sky130_as_sc_hs__diode_2 ANTENNA__28789__A (.DIODE(net209));
 sky130_as_sc_hs__diode_2 ANTENNA__28790__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28792__A (.DIODE(net209));
 sky130_as_sc_hs__diode_2 ANTENNA__28793__A (.DIODE(net358));
 sky130_as_sc_hs__diode_2 ANTENNA__28794__A (.DIODE(net345));
 sky130_as_sc_hs__diode_2 ANTENNA__28796__A (.DIODE(net209));
 sky130_as_sc_hs__diode_2 ANTENNA__28797__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28799__A (.DIODE(net209));
 sky130_as_sc_hs__diode_2 ANTENNA__28800__A (.DIODE(net358));
 sky130_as_sc_hs__diode_2 ANTENNA__28801__A (.DIODE(net234));
 sky130_as_sc_hs__diode_2 ANTENNA__28803__A (.DIODE(net209));
 sky130_as_sc_hs__diode_2 ANTENNA__28804__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__28806__A (.DIODE(net209));
 sky130_as_sc_hs__diode_2 ANTENNA__28807__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28808__A (.DIODE(net345));
 sky130_as_sc_hs__diode_2 ANTENNA__28809__A (.DIODE(net241));
 sky130_as_sc_hs__diode_2 ANTENNA__28810__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__28811__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__28814__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28815__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__28816__A (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__28818__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__28819__A (.DIODE(_19483_));
 sky130_as_sc_hs__diode_2 ANTENNA__28821__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28822__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__28824__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28825__A (.DIODE(net361));
 sky130_as_sc_hs__diode_2 ANTENNA__28826__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__28828__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28829__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__28831__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28832__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__28833__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__28836__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__28839__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__28840__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__28841__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__28842__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__28843__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__28845__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28846__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__28848__A (.DIODE(net204));
 sky130_as_sc_hs__diode_2 ANTENNA__28849__A (.DIODE(net361));
 sky130_as_sc_hs__diode_2 ANTENNA__28850__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__28853__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__28856__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__28857__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__28860__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__28863__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28864__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__28865__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__28867__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__28868__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__28871__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__28872__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__28873__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__28874__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__28877__A (.DIODE(_22301_));
 sky130_as_sc_hs__diode_2 ANTENNA__28881__A (.DIODE(net216));
 sky130_as_sc_hs__diode_2 ANTENNA__28882__A (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__28884__A (.DIODE(net356));
 sky130_as_sc_hs__diode_2 ANTENNA__28885__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__28888__A (.DIODE(net216));
 sky130_as_sc_hs__diode_2 ANTENNA__28889__A (.DIODE(net394));
 sky130_as_sc_hs__diode_2 ANTENNA__28890__B (.DIODE(net394));
 sky130_as_sc_hs__diode_2 ANTENNA__28891__A (.DIODE(net356));
 sky130_as_sc_hs__diode_2 ANTENNA__28892__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__28893__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__28895__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__28898__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__28899__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__28902__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__28905__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__28906__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__28907__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__28908__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__28909__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__28912__A (.DIODE(net218));
 sky130_as_sc_hs__diode_2 ANTENNA__28915__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__28916__A (.DIODE(net234));
 sky130_as_sc_hs__diode_2 ANTENNA__28919__A (.DIODE(net218));
 sky130_as_sc_hs__diode_2 ANTENNA__28922__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__28923__A (.DIODE(net345));
 sky130_as_sc_hs__diode_2 ANTENNA__28926__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__28928__B (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__28929__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__28930__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__28931__A (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__28932__B (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__28933__A (.DIODE(net356));
 sky130_as_sc_hs__diode_2 ANTENNA__28934__A (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__28936__A (.DIODE(net216));
 sky130_as_sc_hs__diode_2 ANTENNA__28937__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__28938__A (.DIODE(net241));
 sky130_as_sc_hs__diode_2 ANTENNA__28939__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__28940__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__28944__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28945__A (.DIODE(net394));
 sky130_as_sc_hs__diode_2 ANTENNA__28947__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__28948__A (.DIODE(net234));
 sky130_as_sc_hs__diode_2 ANTENNA__28951__A (.DIODE(net218));
 sky130_as_sc_hs__diode_2 ANTENNA__28954__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__28955__A (.DIODE(net345));
 sky130_as_sc_hs__diode_2 ANTENNA__28958__A (.DIODE(net218));
 sky130_as_sc_hs__diode_2 ANTENNA__28961__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__28962__A (.DIODE(net234));
 sky130_as_sc_hs__diode_2 ANTENNA__28965__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__28968__A (.DIODE(net218));
 sky130_as_sc_hs__diode_2 ANTENNA__28969__A (.DIODE(net345));
 sky130_as_sc_hs__diode_2 ANTENNA__28970__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__28971__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__28972__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__28975__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28978__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__28979__A (.DIODE(net234));
 sky130_as_sc_hs__diode_2 ANTENNA__28982__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28985__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__28986__A (.DIODE(net345));
 sky130_as_sc_hs__diode_2 ANTENNA__28989__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__28992__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__28993__A (.DIODE(net234));
 sky130_as_sc_hs__diode_2 ANTENNA__28996__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__28999__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__29000__A (.DIODE(net345));
 sky130_as_sc_hs__diode_2 ANTENNA__29001__A (.DIODE(net241));
 sky130_as_sc_hs__diode_2 ANTENNA__29002__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__29003__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__29006__A (.DIODE(_22430_));
 sky130_as_sc_hs__diode_2 ANTENNA__29009__A (.DIODE(net217));
 sky130_as_sc_hs__diode_2 ANTENNA__29012__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__29013__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__29016__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__29019__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__29020__A (.DIODE(net350));
 sky130_as_sc_hs__diode_2 ANTENNA__29022__B (.DIODE(net394));
 sky130_as_sc_hs__diode_2 ANTENNA__29023__A (.DIODE(net218));
 sky130_as_sc_hs__diode_2 ANTENNA__29026__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__29027__A (.DIODE(net234));
 sky130_as_sc_hs__diode_2 ANTENNA__29030__A (.DIODE(net358));
 sky130_as_sc_hs__diode_2 ANTENNA__29033__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__29034__A (.DIODE(net345));
 sky130_as_sc_hs__diode_2 ANTENNA__29035__A (.DIODE(net241));
 sky130_as_sc_hs__diode_2 ANTENNA__29036__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__29037__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__29040__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__29043__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__29044__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__29047__A (.DIODE(net230));
 sky130_as_sc_hs__diode_2 ANTENNA__29050__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__29051__A (.DIODE(net350));
 sky130_as_sc_hs__diode_2 ANTENNA__29054__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__29057__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__29058__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__29061__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__29064__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__29065__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__29066__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__29067__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__29068__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__29073__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__29076__A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA__29077__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__29080__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__29083__A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA__29084__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__29087__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__29090__A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA__29091__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__29094__A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA__29096__B (.DIODE(net408));
 sky130_as_sc_hs__diode_2 ANTENNA__29097__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__29098__A (.DIODE(net350));
 sky130_as_sc_hs__diode_2 ANTENNA__29099__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__29100__A (.DIODE(net341));
 sky130_as_sc_hs__diode_2 ANTENNA__29101__A (.DIODE(\tholin_riscv.Jimm[19] ));
 sky130_as_sc_hs__diode_2 ANTENNA__29104__A (.DIODE(net230));
 sky130_as_sc_hs__diode_2 ANTENNA__29107__A (.DIODE(net370));
 sky130_as_sc_hs__diode_2 ANTENNA__29108__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__29111__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__29114__A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA__29115__A (.DIODE(net350));
 sky130_as_sc_hs__diode_2 ANTENNA__29116__A (.DIODE(net408));
 sky130_as_sc_hs__diode_2 ANTENNA__29118__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__29121__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__29122__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__29125__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__29128__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__29129__A (.DIODE(net350));
 sky130_as_sc_hs__diode_2 ANTENNA__29130__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__29131__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__29132__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__29134__B (.DIODE(_22622_));
 sky130_as_sc_hs__diode_2 ANTENNA__29137__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__29138__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__29140__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__29141__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__29142__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__29143__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__29144__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__29145__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__29146__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__29147__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__29148__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__29149__A (.DIODE(net343));
 sky130_as_sc_hs__diode_2 ANTENNA__29150__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__29151__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__29152__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__29153__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__29154__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__29155__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__29156__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__29158__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__29159__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__29161__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__29162__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__29163__A (.DIODE(net343));
 sky130_as_sc_hs__diode_2 ANTENNA__29164__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__29165__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__29166__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__29167__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__29169__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__29172__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__29173__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__29176__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__29179__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__29180__A (.DIODE(net343));
 sky130_as_sc_hs__diode_2 ANTENNA__29181__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__29183__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__29184__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__29186__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__29187__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__29188__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__29190__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__29191__A (.DIODE(net372));
 sky130_as_sc_hs__diode_2 ANTENNA__29193__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__29194__A (.DIODE(net343));
 sky130_as_sc_hs__diode_2 ANTENNA__29195__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__29196__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__29197__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__29200__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__29201__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__29203__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__29204__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__29205__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__29207__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__29208__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__29210__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__29211__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__29212__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__29213__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__29214__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__29215__A (.DIODE(net219));
 sky130_as_sc_hs__diode_2 ANTENNA__29217__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__29218__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__29219__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__29220__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__29221__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__29222__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__29224__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__29225__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__29226__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__29227__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__29228__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__29229__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__29230__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__29231__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__29232__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__29233__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__29234__A (.DIODE(net210));
 sky130_as_sc_hs__diode_2 ANTENNA__29235__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__29236__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__29237__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__29238__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__29239__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__29240__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__29241__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__29242__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__29243__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__29244__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__29245__A (.DIODE(net201));
 sky130_as_sc_hs__diode_2 ANTENNA__29246__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__29248__A (.DIODE(net210));
 sky130_as_sc_hs__diode_2 ANTENNA__29249__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__29250__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__29252__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__29253__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__29255__A (.DIODE(net203));
 sky130_as_sc_hs__diode_2 ANTENNA__29256__A (.DIODE(net219));
 sky130_as_sc_hs__diode_2 ANTENNA__29257__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__29258__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__29259__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__29260__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__29264__A (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__29265__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__29266__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__29267__A (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__29268__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__29269__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__29270__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__29271__A (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__29272__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__29273__A (.DIODE(net216));
 sky130_as_sc_hs__diode_2 ANTENNA__29274__A (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__29275__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__29276__A (.DIODE(net356));
 sky130_as_sc_hs__diode_2 ANTENNA__29277__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__29278__A (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__29279__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__29280__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__29281__A (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__29282__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__29283__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__29284__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__29285__A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA__29286__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__29287__A (.DIODE(net355));
 sky130_as_sc_hs__diode_2 ANTENNA__29288__A (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__29289__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__29290__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__29291__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__29292__A (.DIODE(net241));
 sky130_as_sc_hs__diode_2 ANTENNA__29293__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__29294__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__29295__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29296__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29297__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__29298__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29299__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29300__A (.DIODE(net356));
 sky130_as_sc_hs__diode_2 ANTENNA__29301__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__29302__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29303__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29304__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__29305__A (.DIODE(net394));
 sky130_as_sc_hs__diode_2 ANTENNA__29306__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29307__A (.DIODE(net356));
 sky130_as_sc_hs__diode_2 ANTENNA__29308__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__29309__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29310__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29311__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__29312__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29313__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29314__A (.DIODE(net356));
 sky130_as_sc_hs__diode_2 ANTENNA__29315__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__29316__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29317__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__29318__A (.DIODE(net356));
 sky130_as_sc_hs__diode_2 ANTENNA__29319__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29320__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29321__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__29322__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__29323__A (.DIODE(net241));
 sky130_as_sc_hs__diode_2 ANTENNA__29324__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__29325__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__29328__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29329__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29330__A (.DIODE(net215));
 sky130_as_sc_hs__diode_2 ANTENNA__29331__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29332__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29333__A (.DIODE(net356));
 sky130_as_sc_hs__diode_2 ANTENNA__29334__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__29335__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29336__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29337__A (.DIODE(net216));
 sky130_as_sc_hs__diode_2 ANTENNA__29338__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29339__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29340__A (.DIODE(net356));
 sky130_as_sc_hs__diode_2 ANTENNA__29341__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__29342__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29343__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29344__A (.DIODE(net216));
 sky130_as_sc_hs__diode_2 ANTENNA__29345__A (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__29346__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__29347__A (.DIODE(net356));
 sky130_as_sc_hs__diode_2 ANTENNA__29348__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__29349__A (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA__29350__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__29351__A (.DIODE(net356));
 sky130_as_sc_hs__diode_2 ANTENNA__29352__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29353__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29354__A (.DIODE(net216));
 sky130_as_sc_hs__diode_2 ANTENNA__29355__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__29356__A (.DIODE(net241));
 sky130_as_sc_hs__diode_2 ANTENNA__29357__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__29358__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__29359__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29360__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29361__A (.DIODE(net218));
 sky130_as_sc_hs__diode_2 ANTENNA__29363__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__29364__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__29365__A (.DIODE(net234));
 sky130_as_sc_hs__diode_2 ANTENNA__29366__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29367__A (.DIODE(net209));
 sky130_as_sc_hs__diode_2 ANTENNA__29368__A (.DIODE(net216));
 sky130_as_sc_hs__diode_2 ANTENNA__29369__A (.DIODE(net389));
 sky130_as_sc_hs__diode_2 ANTENNA__29370__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29371__A (.DIODE(net356));
 sky130_as_sc_hs__diode_2 ANTENNA__29372__A (.DIODE(net344));
 sky130_as_sc_hs__diode_2 ANTENNA__29374__A (.DIODE(net207));
 sky130_as_sc_hs__diode_2 ANTENNA__29375__A (.DIODE(net218));
 sky130_as_sc_hs__diode_2 ANTENNA__29377__A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA__29378__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__29379__A (.DIODE(net233));
 sky130_as_sc_hs__diode_2 ANTENNA__29381__A (.DIODE(net209));
 sky130_as_sc_hs__diode_2 ANTENNA__29382__A (.DIODE(net357));
 sky130_as_sc_hs__diode_2 ANTENNA__29384__A (.DIODE(net209));
 sky130_as_sc_hs__diode_2 ANTENNA__29385__A (.DIODE(net218));
 sky130_as_sc_hs__diode_2 ANTENNA__29386__A (.DIODE(net345));
 sky130_as_sc_hs__diode_2 ANTENNA__29387__A (.DIODE(net241));
 sky130_as_sc_hs__diode_2 ANTENNA__29388__A (.DIODE(net338));
 sky130_as_sc_hs__diode_2 ANTENNA__29389__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__29392__A (.DIODE(_22624_));
 sky130_as_sc_hs__diode_2 ANTENNA__29396__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29400__A (.DIODE(net239));
 sky130_as_sc_hs__diode_2 ANTENNA__29403__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29407__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__29410__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__29414__A (.DIODE(net239));
 sky130_as_sc_hs__diode_2 ANTENNA__29420__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__29421__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__29422__A (.DIODE(net244));
 sky130_as_sc_hs__diode_2 ANTENNA__29423__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__29424__A (.DIODE(\tholin_riscv.Jimm[19] ));
 sky130_as_sc_hs__diode_2 ANTENNA__29427__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__29430__A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA__29431__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__29434__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__29437__A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA__29438__A (.DIODE(net350));
 sky130_as_sc_hs__diode_2 ANTENNA__29441__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__29444__A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA__29445__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__29448__A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA__29449__A (.DIODE(net408));
 sky130_as_sc_hs__diode_2 ANTENNA__29451__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__29452__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__29453__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__29454__A (.DIODE(net341));
 sky130_as_sc_hs__diode_2 ANTENNA__29455__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__29462__A (.DIODE(net224));
 sky130_as_sc_hs__diode_2 ANTENNA__29463__A (.DIODE(net400));
 sky130_as_sc_hs__diode_2 ANTENNA__29465__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__29466__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__29469__A (.DIODE(net224));
 sky130_as_sc_hs__diode_2 ANTENNA__29470__A (.DIODE(net400));
 sky130_as_sc_hs__diode_2 ANTENNA__29472__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__29473__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__29476__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__29479__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__29480__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__29483__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__29486__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__29487__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__29488__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__29489__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__29490__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__29494__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__29497__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__29500__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29504__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__29510__A (.DIODE(net370));
 sky130_as_sc_hs__diode_2 ANTENNA__29511__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__29518__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__29519__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__29520__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__29526__A (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA__29528__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__29529__A (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA__29531__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__29532__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__29535__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__29538__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__29539__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__29542__A (.DIODE(net224));
 sky130_as_sc_hs__diode_2 ANTENNA__29545__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__29546__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__29549__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__29552__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__29553__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__29554__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__29555__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__29556__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__29557__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__29560__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__29562__A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA__29563__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__29566__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29569__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29570__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__29571__A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA__29573__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29576__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29577__A (.DIODE(net239));
 sky130_as_sc_hs__diode_2 ANTENNA__29580__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29583__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29584__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__29585__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__29586__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__29587__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__29592__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__29595__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__29596__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__29599__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__29602__A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA__29603__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__29606__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__29609__A (.DIODE(net361));
 sky130_as_sc_hs__diode_2 ANTENNA__29610__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__29613__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__29616__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__29617__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__29618__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__29619__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__29620__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__29621__A (.DIODE(net375));
 sky130_as_sc_hs__diode_2 ANTENNA__29623__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__29626__A (.DIODE(net361));
 sky130_as_sc_hs__diode_2 ANTENNA__29627__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__29630__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__29633__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__29634__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__29637__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__29640__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__29641__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__29644__A (.DIODE(net361));
 sky130_as_sc_hs__diode_2 ANTENNA__29647__A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA__29648__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__29649__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__29650__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__29651__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__29655__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29658__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29659__A (.DIODE(net239));
 sky130_as_sc_hs__diode_2 ANTENNA__29662__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29665__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29666__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__29669__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29672__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29673__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__29676__A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA__29679__A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA__29680__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__29681__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__29682__A (.DIODE(net341));
 sky130_as_sc_hs__diode_2 ANTENNA__29683__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__29686__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__29689__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__29690__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__29693__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__29696__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__29697__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__29700__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__29703__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__29704__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__29707__A (.DIODE(net366));
 sky130_as_sc_hs__diode_2 ANTENNA__29710__A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA__29711__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__29712__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__29713__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__29714__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__29719__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29722__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29723__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__29726__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29729__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29730__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__29733__A (.DIODE(net224));
 sky130_as_sc_hs__diode_2 ANTENNA__29734__A (.DIODE(net400));
 sky130_as_sc_hs__diode_2 ANTENNA__29736__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29737__A (.DIODE(net239));
 sky130_as_sc_hs__diode_2 ANTENNA__29740__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29743__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__29744__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__29745__A (.DIODE(net243));
 sky130_as_sc_hs__diode_2 ANTENNA__29746__A (.DIODE(net341));
 sky130_as_sc_hs__diode_2 ANTENNA__29747__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__29750__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__29753__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__29754__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__29757__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__29760__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__29761__A (.DIODE(\tholin_riscv.Jimm[17] ));
 sky130_as_sc_hs__diode_2 ANTENNA__29764__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__29767__A (.DIODE(net362));
 sky130_as_sc_hs__diode_2 ANTENNA__29768__A (.DIODE(net235));
 sky130_as_sc_hs__diode_2 ANTENNA__29771__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29774__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__29775__A (.DIODE(net346));
 sky130_as_sc_hs__diode_2 ANTENNA__29776__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__29777__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__29778__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__29781__A (.DIODE(_23141_));
 sky130_as_sc_hs__diode_2 ANTENNA__29785__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__29789__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__29792__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__29795__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29796__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__29799__A (.DIODE(net220));
 sky130_as_sc_hs__diode_2 ANTENNA__29803__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__29809__A (.DIODE(net222));
 sky130_as_sc_hs__diode_2 ANTENNA__29810__A (.DIODE(net348));
 sky130_as_sc_hs__diode_2 ANTENNA__29811__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__29812__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__29813__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__29816__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29819__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29820__A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA__29823__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29826__A (.DIODE(net367));
 sky130_as_sc_hs__diode_2 ANTENNA__29827__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__29834__A (.DIODE(net237));
 sky130_as_sc_hs__diode_2 ANTENNA__29840__A (.DIODE(net228));
 sky130_as_sc_hs__diode_2 ANTENNA__29841__A (.DIODE(net349));
 sky130_as_sc_hs__diode_2 ANTENNA__29842__A (.DIODE(net244));
 sky130_as_sc_hs__diode_2 ANTENNA__29843__A (.DIODE(net339));
 sky130_as_sc_hs__diode_2 ANTENNA__29844__A (.DIODE(net245));
 sky130_as_sc_hs__diode_2 ANTENNA__29848__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__29852__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__29855__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__29859__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__29862__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__29865__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__29866__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__29869__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__29872__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__29873__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__29874__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__29875__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__29876__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__29879__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__29883__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__29886__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__29889__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__29890__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__29893__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__29896__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__29897__A (.DIODE(net236));
 sky130_as_sc_hs__diode_2 ANTENNA__29900__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__29903__A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA__29904__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__29905__A (.DIODE(net242));
 sky130_as_sc_hs__diode_2 ANTENNA__29906__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__29907__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__29916__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__29923__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__29930__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__29936__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__29937__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__29938__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__29939__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__29940__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__29947__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__29954__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__29961__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__29968__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__29969__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__29970__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__29971__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__29976__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__29980__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__29983__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__29987__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__29990__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__29994__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__30000__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__30001__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__30002__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__30003__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__30004__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__30007__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__30011__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__30014__A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA__30018__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__30021__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__30025__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__30028__A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA__30031__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__30032__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__30033__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__30034__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__30035__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__30044__A (.DIODE(_21659_));
 sky130_as_sc_hs__diode_2 ANTENNA__30046__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__30046__B (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA__30052__A (.DIODE(net274));
 sky130_as_sc_hs__diode_2 ANTENNA__30053__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__30060__A (.DIODE(net259));
 sky130_as_sc_hs__diode_2 ANTENNA__30066__A (.DIODE(net274));
 sky130_as_sc_hs__diode_2 ANTENNA__30067__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__30070__A (.DIODE(net274));
 sky130_as_sc_hs__diode_2 ANTENNA__30074__A (.DIODE(net259));
 sky130_as_sc_hs__diode_2 ANTENNA__30075__A (.DIODE(net153));
 sky130_as_sc_hs__diode_2 ANTENNA__30076__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__30077__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__30084__A (.DIODE(net160));
 sky130_as_sc_hs__diode_2 ANTENNA__30091__A (.DIODE(net259));
 sky130_as_sc_hs__diode_2 ANTENNA__30098__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__30105__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__30106__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__30107__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__30108__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__30110__B (.DIODE(\tholin_riscv.Jimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__30112__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__30113__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__30114__A (.DIODE(\tholin_riscv.Jimm[13] ));
 sky130_as_sc_hs__diode_2 ANTENNA__30114__B (.DIODE(\tholin_riscv.Jimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__30115__A (.DIODE(\tholin_riscv.Jimm[13] ));
 sky130_as_sc_hs__diode_2 ANTENNA__30115__B (.DIODE(\tholin_riscv.Jimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__30116__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__30117__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__30117__B (.DIODE(\tholin_riscv.Jimm[13] ));
 sky130_as_sc_hs__diode_2 ANTENNA__30118__A (.DIODE(_23598_));
 sky130_as_sc_hs__diode_2 ANTENNA__30122__A (.DIODE(_21140_));
 sky130_as_sc_hs__diode_2 ANTENNA__30125__A (.DIODE(_21343_));
 sky130_as_sc_hs__diode_2 ANTENNA__30125__B (.DIODE(_21440_));
 sky130_as_sc_hs__diode_2 ANTENNA__30141__B (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__30143__A (.DIODE(_21440_));
 sky130_as_sc_hs__diode_2 ANTENNA__30155__B (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__30162__B (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__30169__B (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__30181__A (.DIODE(_21659_));
 sky130_as_sc_hs__diode_2 ANTENNA__30186__B (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__30192__B (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__30201__A (.DIODE(_21659_));
 sky130_as_sc_hs__diode_2 ANTENNA__30203__A (.DIODE(net115));
 sky130_as_sc_hs__diode_2 ANTENNA__30203__B (.DIODE(net121));
 sky130_as_sc_hs__diode_2 ANTENNA__30214__A (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__30214__B (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__30226__A (.DIODE(net172));
 sky130_as_sc_hs__diode_2 ANTENNA__30229__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30230__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__30233__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__30237__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__30240__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30243__A (.DIODE(net269));
 sky130_as_sc_hs__diode_2 ANTENNA__30244__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__30247__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30250__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30251__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__30252__A (.DIODE(net156));
 sky130_as_sc_hs__diode_2 ANTENNA__30253__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__30254__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__30257__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30260__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30261__A (.DIODE(net165));
 sky130_as_sc_hs__diode_2 ANTENNA__30264__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30266__A (.DIODE(net306));
 sky130_as_sc_hs__diode_2 ANTENNA__30267__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30268__A (.DIODE(_00002_));
 sky130_as_sc_hs__diode_2 ANTENNA__30271__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30274__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30275__A (.DIODE(net165));
 sky130_as_sc_hs__diode_2 ANTENNA__30278__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30281__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30282__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__30283__A (.DIODE(net156));
 sky130_as_sc_hs__diode_2 ANTENNA__30284__A (.DIODE(net253));
 sky130_as_sc_hs__diode_2 ANTENNA__30285__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__30290__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30293__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30294__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__30296__A (.DIODE(net306));
 sky130_as_sc_hs__diode_2 ANTENNA__30297__A (.DIODE(net172));
 sky130_as_sc_hs__diode_2 ANTENNA__30299__A (.DIODE(net306));
 sky130_as_sc_hs__diode_2 ANTENNA__30300__A (.DIODE(net269));
 sky130_as_sc_hs__diode_2 ANTENNA__30301__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__30304__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30307__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30308__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__30310__A (.DIODE(net306));
 sky130_as_sc_hs__diode_2 ANTENNA__30311__A (.DIODE(net269));
 sky130_as_sc_hs__diode_2 ANTENNA__30313__A (.DIODE(net306));
 sky130_as_sc_hs__diode_2 ANTENNA__30314__A (.DIODE(net172));
 sky130_as_sc_hs__diode_2 ANTENNA__30315__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__30316__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__30317__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__30318__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__30321__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__30324__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__30325__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__30328__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__30331__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__30332__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__30334__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__30335__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__30338__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__30339__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__30341__A (.DIODE(net333));
 sky130_as_sc_hs__diode_2 ANTENNA__30342__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__30345__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__30346__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__30347__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__30348__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__30349__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__30353__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30356__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30357__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__30360__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30363__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30364__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__30367__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30370__A (.DIODE(net269));
 sky130_as_sc_hs__diode_2 ANTENNA__30371__A (.DIODE(net165));
 sky130_as_sc_hs__diode_2 ANTENNA__30374__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30377__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30378__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__30379__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__30380__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__30381__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__30384__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__30387__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__30388__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__30391__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__30393__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__30394__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__30395__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__30397__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__30398__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__30400__A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA__30401__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__30402__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__30405__A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA__30408__A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA__30409__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__30410__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__30411__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__30412__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__30421__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__30427__A (.DIODE(net281));
 sky130_as_sc_hs__diode_2 ANTENNA__30428__A (.DIODE(net262));
 sky130_as_sc_hs__diode_2 ANTENNA__30435__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__30438__A (.DIODE(net281));
 sky130_as_sc_hs__diode_2 ANTENNA__30441__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__30442__A (.DIODE(net262));
 sky130_as_sc_hs__diode_2 ANTENNA__30443__A (.DIODE(net156));
 sky130_as_sc_hs__diode_2 ANTENNA__30444__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__30445__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__30448__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__30451__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__30452__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__30455__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__30458__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__30459__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__30462__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__30466__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__30469__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__30472__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__30473__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__30474__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__30475__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__30476__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__30480__A (.DIODE(_20622_));
 sky130_as_sc_hs__diode_2 ANTENNA__30480__B (.DIODE(_20707_));
 sky130_as_sc_hs__diode_2 ANTENNA__30488__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__30492__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__30495__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__30499__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__30502__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__30506__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__30512__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__30513__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__30514__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__30515__A (.DIODE(net253));
 sky130_as_sc_hs__diode_2 ANTENNA__30516__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__30519__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__30522__A (.DIODE(net281));
 sky130_as_sc_hs__diode_2 ANTENNA__30523__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__30526__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__30529__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__30530__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__30533__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__30536__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__30537__A (.DIODE(net165));
 sky130_as_sc_hs__diode_2 ANTENNA__30540__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__30543__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__30544__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__30545__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__30546__A (.DIODE(net253));
 sky130_as_sc_hs__diode_2 ANTENNA__30547__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__30559__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__30559__B (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__30561__A (.DIODE(_21977_));
 sky130_as_sc_hs__diode_2 ANTENNA__30567__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__30571__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__30574__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__30578__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__30581__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__30585__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__30592__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__30593__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__30594__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__30595__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__30598__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__30601__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__30602__A (.DIODE(net165));
 sky130_as_sc_hs__diode_2 ANTENNA__30605__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__30608__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__30609__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__30616__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__30619__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__30622__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__30623__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__30624__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__30625__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__30626__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__30635__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__30635__B (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__30636__A (.DIODE(_21659_));
 sky130_as_sc_hs__diode_2 ANTENNA__30642__A (.DIODE(net169));
 sky130_as_sc_hs__diode_2 ANTENNA__30645__A (.DIODE(net266));
 sky130_as_sc_hs__diode_2 ANTENNA__30646__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__30649__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30652__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30653__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__30656__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30659__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30660__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__30663__A (.DIODE(net266));
 sky130_as_sc_hs__diode_2 ANTENNA__30666__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__30667__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__30668__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__30669__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__30670__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__30673__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__30677__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__30680__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__30684__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__30687__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__30691__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__30697__A (.DIODE(net180));
 sky130_as_sc_hs__diode_2 ANTENNA__30698__A (.DIODE(net262));
 sky130_as_sc_hs__diode_2 ANTENNA__30699__A (.DIODE(net156));
 sky130_as_sc_hs__diode_2 ANTENNA__30700__A (.DIODE(net253));
 sky130_as_sc_hs__diode_2 ANTENNA__30701__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__30710__A (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__30711__B (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__30711__C (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__30722__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__30722__B (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__30726__A (.DIODE(_21659_));
 sky130_as_sc_hs__diode_2 ANTENNA__30733__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__30733__B (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__30739__A (.DIODE(_21659_));
 sky130_as_sc_hs__diode_2 ANTENNA__30746__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__30746__B (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__30756__C (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__30759__A (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__30759__B (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__30766__A (.DIODE(_21659_));
 sky130_as_sc_hs__diode_2 ANTENNA__30768__A (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__30768__B (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__30769__A (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__30769__B (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__30770__A (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__30770__B (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__30784__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__30787__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__30788__A (.DIODE(net332));
 sky130_as_sc_hs__diode_2 ANTENNA__30789__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__30790__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__30791__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__30794__A (.DIODE(net196));
 sky130_as_sc_hs__diode_2 ANTENNA__30796__A (.DIODE(net281));
 sky130_as_sc_hs__diode_2 ANTENNA__30797__A (.DIODE(net260));
 sky130_as_sc_hs__diode_2 ANTENNA__30800__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__30803__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__30804__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__30806__A (.DIODE(net332));
 sky130_as_sc_hs__diode_2 ANTENNA__30807__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__30810__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__30811__A (.DIODE(net262));
 sky130_as_sc_hs__diode_2 ANTENNA__30812__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__30813__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__30815__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__30816__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__30818__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__30819__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__30821__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__30822__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__30823__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__30824__A (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__30825__A (.DIODE(net166));
 sky130_as_sc_hs__diode_2 ANTENNA__30826__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__30828__A (.DIODE(net263));
 sky130_as_sc_hs__diode_2 ANTENNA__30829__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__30830__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__30831__A (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__30832__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__30833__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__30834__A (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__30835__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__30836__A (.DIODE(net157));
 sky130_as_sc_hs__diode_2 ANTENNA__30837__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__30838__A (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__30839__A (.DIODE(net270));
 sky130_as_sc_hs__diode_2 ANTENNA__30840__A (.DIODE(net187));
 sky130_as_sc_hs__diode_2 ANTENNA__30841__A (.DIODE(net308));
 sky130_as_sc_hs__diode_2 ANTENNA__30842__A (.DIODE(net174));
 sky130_as_sc_hs__diode_2 ANTENNA__30843__A (.DIODE(net257));
 sky130_as_sc_hs__diode_2 ANTENNA__30844__A (.DIODE(net153));
 sky130_as_sc_hs__diode_2 ANTENNA__30845__A (.DIODE(net250));
 sky130_as_sc_hs__diode_2 ANTENNA__30847__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__30854__A (.DIODE(net169));
 sky130_as_sc_hs__diode_2 ANTENNA__30857__A (.DIODE(net266));
 sky130_as_sc_hs__diode_2 ANTENNA__30858__A (.DIODE(net162));
 sky130_as_sc_hs__diode_2 ANTENNA__30861__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__30864__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__30865__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__30868__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__30871__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__30872__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__30875__A (.DIODE(net265));
 sky130_as_sc_hs__diode_2 ANTENNA__30878__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__30879__A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA__30880__A (.DIODE(net154));
 sky130_as_sc_hs__diode_2 ANTENNA__30881__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__30882__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__30885__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__30888__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__30889__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__30892__A (.DIODE(net171));
 sky130_as_sc_hs__diode_2 ANTENNA__30895__A (.DIODE(net268));
 sky130_as_sc_hs__diode_2 ANTENNA__30896__A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA__30899__A (.DIODE(net170));
 sky130_as_sc_hs__diode_2 ANTENNA__30902__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__30903__A (.DIODE(net161));
 sky130_as_sc_hs__diode_2 ANTENNA__30906__A (.DIODE(net267));
 sky130_as_sc_hs__diode_2 ANTENNA__30909__A (.DIODE(net168));
 sky130_as_sc_hs__diode_2 ANTENNA__30910__A (.DIODE(net254));
 sky130_as_sc_hs__diode_2 ANTENNA__30911__A (.DIODE(net156));
 sky130_as_sc_hs__diode_2 ANTENNA__30912__A (.DIODE(net251));
 sky130_as_sc_hs__diode_2 ANTENNA__30913__A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA__30926__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__30929__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__30932__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__30933__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__30935__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__30936__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__30940__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__30946__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__30947__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__30948__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__30949__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__30950__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__30952__A (.DIODE(net320));
 sky130_as_sc_hs__diode_2 ANTENNA__30954__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__30957__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__30958__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__30960__A (.DIODE(net179));
 sky130_as_sc_hs__diode_2 ANTENNA__30962__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__30964__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__30967__A (.DIODE(net179));
 sky130_as_sc_hs__diode_2 ANTENNA__30970__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__30971__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__30974__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__30977__A (.DIODE(net179));
 sky130_as_sc_hs__diode_2 ANTENNA__30978__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__30979__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__30980__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__30981__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__30985__A (.DIODE(_24337_));
 sky130_as_sc_hs__diode_2 ANTENNA__30986__A (.DIODE(_24337_));
 sky130_as_sc_hs__diode_2 ANTENNA__30991__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__30991__B (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__30992__A (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__30992__B (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__30994__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__31007__B (.DIODE(_22622_));
 sky130_as_sc_hs__diode_2 ANTENNA__31008__B (.DIODE(_22622_));
 sky130_as_sc_hs__diode_2 ANTENNA__31013__A (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__31013__B (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__31014__A (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__31014__B (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__31015__A (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__31015__B (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__31039__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__31039__B (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__31043__A (.DIODE(_20622_));
 sky130_as_sc_hs__diode_2 ANTENNA__31044__B (.DIODE(_20707_));
 sky130_as_sc_hs__diode_2 ANTENNA__31047__A (.DIODE(_20707_));
 sky130_as_sc_hs__diode_2 ANTENNA__31048__B (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__31049__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__31049__C (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__31050__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__31057__A (.DIODE(_20622_));
 sky130_as_sc_hs__diode_2 ANTENNA__31060__A (.DIODE(_20622_));
 sky130_as_sc_hs__diode_2 ANTENNA__31062__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__31062__B (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__31073__A (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__31073__B (.DIODE(net455));
 sky130_as_sc_hs__diode_2 ANTENNA__31074__B (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__31074__C (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__31085__A (.DIODE(_22430_));
 sky130_as_sc_hs__diode_2 ANTENNA__31097__A (.DIODE(net453));
 sky130_as_sc_hs__diode_2 ANTENNA__31097__B (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__31098__A (.DIODE(_22430_));
 sky130_as_sc_hs__diode_2 ANTENNA__31101__A (.DIODE(_21659_));
 sky130_as_sc_hs__diode_2 ANTENNA__31101__B (.DIODE(_22430_));
 sky130_as_sc_hs__diode_2 ANTENNA__31108__A (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__31108__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__31116__A (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__31116__B (.DIODE(net86));
 sky130_as_sc_hs__diode_2 ANTENNA__31117__B (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__31117__C (.DIODE(net455));
 sky130_as_sc_hs__diode_2 ANTENNA__31134__A (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__31134__B (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__31135__A (.DIODE(net453));
 sky130_as_sc_hs__diode_2 ANTENNA__31135__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__31150__A (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__31150__B (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__31151__A (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__31151__B (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__31153__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__31168__A (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__31168__B (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__31169__A (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__31169__B (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__31170__A (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__31170__B (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__31192__A (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__31192__B (.DIODE(net453));
 sky130_as_sc_hs__diode_2 ANTENNA__31193__B (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__31193__C (.DIODE(net86));
 sky130_as_sc_hs__diode_2 ANTENNA__31208__A (.DIODE(_21659_));
 sky130_as_sc_hs__diode_2 ANTENNA__31210__A (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__31210__B (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__31211__A (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__31211__B (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__31235__A (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__31235__B (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__31241__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__31241__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__31248__A (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__31248__B (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__31254__A (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__31254__B (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__31259__A (.DIODE(net455));
 sky130_as_sc_hs__diode_2 ANTENNA__31259__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__31260__A (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__31260__B (.DIODE(net86));
 sky130_as_sc_hs__diode_2 ANTENNA__31265__A (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__31265__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__31266__A (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__31266__B (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__31280__A (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__31280__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__31286__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__31286__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__31292__A (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__31292__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__31299__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__31299__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__31300__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__31300__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__31307__A (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__31307__B (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__31316__A (.DIODE(_21140_));
 sky130_as_sc_hs__diode_2 ANTENNA__31320__A (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__31320__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__31326__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__31326__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__31332__A (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__31333__A (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__31333__C (.DIODE(net437));
 sky130_as_sc_hs__diode_2 ANTENNA__31345__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__31345__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__31346__A (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__31353__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__31359__A (.DIODE(net281));
 sky130_as_sc_hs__diode_2 ANTENNA__31360__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__31363__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__31366__A (.DIODE(net281));
 sky130_as_sc_hs__diode_2 ANTENNA__31367__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__31370__A (.DIODE(net281));
 sky130_as_sc_hs__diode_2 ANTENNA__31373__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__31374__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__31375__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__31376__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__31377__A (.DIODE(net247));
 sky130_as_sc_hs__diode_2 ANTENNA__31380__A (.DIODE(net179));
 sky130_as_sc_hs__diode_2 ANTENNA__31383__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__31384__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__31387__A (.DIODE(net179));
 sky130_as_sc_hs__diode_2 ANTENNA__31390__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__31391__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__31394__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__31397__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__31398__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__31401__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__31404__A (.DIODE(net179));
 sky130_as_sc_hs__diode_2 ANTENNA__31405__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__31406__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__31407__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__31408__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__31434__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__31434__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__31435__A (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__31435__B (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__31436__A (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__31436__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__31446__A (.DIODE(_23141_));
 sky130_as_sc_hs__diode_2 ANTENNA__31449__A (.DIODE(_21659_));
 sky130_as_sc_hs__diode_2 ANTENNA__31449__B (.DIODE(_23141_));
 sky130_as_sc_hs__diode_2 ANTENNA__31451__A (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__31451__B (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__31452__A (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__31452__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__31453__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__31454__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__31454__B (.DIODE(net437));
 sky130_as_sc_hs__diode_2 ANTENNA__31476__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__31478__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__31479__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__31481__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__31482__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__31483__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__31485__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__31486__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__31487__A (.DIODE(net332));
 sky130_as_sc_hs__diode_2 ANTENNA__31488__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__31489__A (.DIODE(net262));
 sky130_as_sc_hs__diode_2 ANTENNA__31490__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__31492__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__31493__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__31495__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__31496__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__31497__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__31498__A (.DIODE(net332));
 sky130_as_sc_hs__diode_2 ANTENNA__31499__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__31500__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__31501__A (.DIODE(net332));
 sky130_as_sc_hs__diode_2 ANTENNA__31502__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__31503__A (.DIODE(net262));
 sky130_as_sc_hs__diode_2 ANTENNA__31504__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__31505__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__31506__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__31509__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__31512__A (.DIODE(net275));
 sky130_as_sc_hs__diode_2 ANTENNA__31513__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__31516__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__31517__A (.DIODE(net195));
 sky130_as_sc_hs__diode_2 ANTENNA__31519__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__31520__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__31523__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__31524__A (.DIODE(net195));
 sky130_as_sc_hs__diode_2 ANTENNA__31526__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__31527__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__31528__A (.DIODE(net195));
 sky130_as_sc_hs__diode_2 ANTENNA__31530__A (.DIODE(net272));
 sky130_as_sc_hs__diode_2 ANTENNA__31531__A (.DIODE(net195));
 sky130_as_sc_hs__diode_2 ANTENNA__31533__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__31534__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__31535__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__31536__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__31537__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__31547__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__31547__B (.DIODE(_25035_));
 sky130_as_sc_hs__diode_2 ANTENNA__31548__A (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__31548__B (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__31552__A (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__31552__B (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__31553__C (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__31569__A (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__31569__B (.DIODE(net455));
 sky130_as_sc_hs__diode_2 ANTENNA__31570__A (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__31570__B (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__31571__A (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__31571__B (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__31592__A (.DIODE(_24550_));
 sky130_as_sc_hs__diode_2 ANTENNA__31592__B (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__31593__B (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__31593__C (.DIODE(net453));
 sky130_as_sc_hs__diode_2 ANTENNA__31605__A (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__31605__B (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__31606__A (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__31606__B (.DIODE(net443));
 sky130_as_sc_hs__diode_2 ANTENNA__31628__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__31628__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__31629__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__31629__B (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__31630__A (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__31630__B (.DIODE(net435));
 sky130_as_sc_hs__diode_2 ANTENNA__31652__A (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__31652__B (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__31653__A (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__31653__B (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__31654__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__31655__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__31655__B (.DIODE(net437));
 sky130_as_sc_hs__diode_2 ANTENNA__31661__A (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__31661__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__31662__A (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__31662__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__31663__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__31663__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__31692__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__31692__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__31693__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__31693__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__31700__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__31700__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__31701__A (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__31701__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__31702__A (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__31703__A (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__31703__B (.DIODE(net437));
 sky130_as_sc_hs__diode_2 ANTENNA__31717__A (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__31717__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__31723__A (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__31723__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__31730__A (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__31730__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__31731__A (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__31731__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__31737__A (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__31737__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__31738__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__31739__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__31739__B (.DIODE(net437));
 sky130_as_sc_hs__diode_2 ANTENNA__31740__A (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__31740__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__31748__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__31748__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__31749__A (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__31749__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__31767__A (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__31767__B (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__31768__A (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__31768__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__31787__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__31787__B (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__31793__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__31793__B (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__31796__B (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__31797__B (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__31807__B (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__31808__B (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__31811__A (.DIODE(net115));
 sky130_as_sc_hs__diode_2 ANTENNA__31811__B (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__31829__A (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__31829__B (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__31830__A (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__31830__B (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__31849__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__31849__B (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__31873__A (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__31873__B (.DIODE(_25035_));
 sky130_as_sc_hs__diode_2 ANTENNA__31874__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__31874__B (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__31881__A (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__31881__B (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__31882__C (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__31898__A (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__31898__B (.DIODE(net86));
 sky130_as_sc_hs__diode_2 ANTENNA__31899__A (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__31899__B (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__31900__A (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__31900__B (.DIODE(net455));
 sky130_as_sc_hs__diode_2 ANTENNA__31921__A (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__31921__B (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__31922__B (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__31922__C (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__31934__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__31934__B (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__31935__A (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__31936__A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA__31938__A (.DIODE(net186));
 sky130_as_sc_hs__diode_2 ANTENNA__31941__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__31942__A (.DIODE(net164));
 sky130_as_sc_hs__diode_2 ANTENNA__31945__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__31948__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__31949__A (.DIODE(net262));
 sky130_as_sc_hs__diode_2 ANTENNA__31952__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__31955__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__31956__A (.DIODE(net165));
 sky130_as_sc_hs__diode_2 ANTENNA__31959__A (.DIODE(net280));
 sky130_as_sc_hs__diode_2 ANTENNA__31962__A (.DIODE(net185));
 sky130_as_sc_hs__diode_2 ANTENNA__31963__A (.DIODE(net262));
 sky130_as_sc_hs__diode_2 ANTENNA__31964__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__31965__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__31966__A (.DIODE(_00004_));
 sky130_as_sc_hs__diode_2 ANTENNA__31969__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__31972__A (.DIODE(net275));
 sky130_as_sc_hs__diode_2 ANTENNA__31973__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__31976__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__31979__A (.DIODE(net275));
 sky130_as_sc_hs__diode_2 ANTENNA__31980__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__31983__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__31986__A (.DIODE(net275));
 sky130_as_sc_hs__diode_2 ANTENNA__31987__A (.DIODE(net158));
 sky130_as_sc_hs__diode_2 ANTENNA__31990__A (.DIODE(net275));
 sky130_as_sc_hs__diode_2 ANTENNA__31993__A (.DIODE(net176));
 sky130_as_sc_hs__diode_2 ANTENNA__31994__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__31995__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__31996__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__31997__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__32031__A (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__32031__B (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__32032__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__32032__B (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__32033__A (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__32033__B (.DIODE(net435));
 sky130_as_sc_hs__diode_2 ANTENNA__32050__A (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__32050__B (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__32051__A (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__32051__B (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__32052__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__32053__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__32053__B (.DIODE(net437));
 sky130_as_sc_hs__diode_2 ANTENNA__32059__A (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__32059__B (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__32060__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__32060__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__32061__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__32061__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__32096__A (.DIODE(net121));
 sky130_as_sc_hs__diode_2 ANTENNA__32096__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__32097__A (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__32097__B (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__32142__A (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__32142__B (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__32143__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__32143__B (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__32150__A (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__32150__B (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__32151__C (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__32167__A (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__32167__B (.DIODE(net453));
 sky130_as_sc_hs__diode_2 ANTENNA__32168__A (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__32168__B (.DIODE(net455));
 sky130_as_sc_hs__diode_2 ANTENNA__32169__A (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__32169__B (.DIODE(net86));
 sky130_as_sc_hs__diode_2 ANTENNA__32190__A (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__32190__B (.DIODE(net443));
 sky130_as_sc_hs__diode_2 ANTENNA__32192__B (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__32192__C (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__32203__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__32203__B (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__32204__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__32204__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__32205__A (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__32205__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__32231__A (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__32231__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__32232__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__32232__B (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__32233__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__32233__B (.DIODE(net435));
 sky130_as_sc_hs__diode_2 ANTENNA__32250__A (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__32250__B (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__32252__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__32259__A (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__32259__B (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__32260__A (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__32260__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__32261__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__32261__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__32295__A (.DIODE(net121));
 sky130_as_sc_hs__diode_2 ANTENNA__32295__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__32296__A (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA__32296__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__32316__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__32316__B (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__32323__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__32330__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__32333__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__32336__A (.DIODE(net359));
 sky130_as_sc_hs__diode_2 ANTENNA__32337__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__32340__A (.DIODE(net359));
 sky130_as_sc_hs__diode_2 ANTENNA__32343__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__32344__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__32345__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__32346__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__32347__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__32350__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__32353__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__32354__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__32357__A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA__32360__A (.DIODE(net359));
 sky130_as_sc_hs__diode_2 ANTENNA__32361__A (.DIODE(net343));
 sky130_as_sc_hs__diode_2 ANTENNA__32367__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__32368__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__32371__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__32375__A (.DIODE(net343));
 sky130_as_sc_hs__diode_2 ANTENNA__32376__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__32377__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__32378__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__32386__A (.DIODE(net115));
 sky130_as_sc_hs__diode_2 ANTENNA__32386__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__32387__B (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__32388__B (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__32395__A (.DIODE(net165));
 sky130_as_sc_hs__diode_2 ANTENNA__32402__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__32403__A (.DIODE(net198));
 sky130_as_sc_hs__diode_2 ANTENNA__32406__A (.DIODE(net198));
 sky130_as_sc_hs__diode_2 ANTENNA__32409__A (.DIODE(net165));
 sky130_as_sc_hs__diode_2 ANTENNA__32412__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__32413__A (.DIODE(net198));
 sky130_as_sc_hs__diode_2 ANTENNA__32416__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__32417__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__32418__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__32419__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__32420__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__32421__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__32424__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__32425__A (.DIODE(net274));
 sky130_as_sc_hs__diode_2 ANTENNA__32426__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__32428__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__32431__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__32433__A (.DIODE(net259));
 sky130_as_sc_hs__diode_2 ANTENNA__32435__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__32438__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__32440__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__32441__A (.DIODE(net193));
 sky130_as_sc_hs__diode_2 ANTENNA__32442__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__32445__A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA__32447__A (.DIODE(net259));
 sky130_as_sc_hs__diode_2 ANTENNA__32448__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__32449__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__32450__A (.DIODE(net150));
 sky130_as_sc_hs__diode_2 ANTENNA__32459__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__32459__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__32505__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__32505__B (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__32506__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__32506__B (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__32508__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__32508__B (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__32513__A (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__32513__B (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__32514__A (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__32515__A (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__32515__B (.DIODE(net467));
 sky130_as_sc_hs__diode_2 ANTENNA__32516__B (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__32535__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__32535__B (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__32536__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__32536__C (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__32537__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__32537__B (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__32538__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__32538__B (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__32570__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__32570__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__32571__A (.DIODE(net455));
 sky130_as_sc_hs__diode_2 ANTENNA__32571__B (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__32576__A (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__32576__B (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__32577__A (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__32577__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__32606__A (.DIODE(net443));
 sky130_as_sc_hs__diode_2 ANTENNA__32606__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__32607__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__32607__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__32621__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__32621__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__32622__A (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__32622__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__32627__A (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__32627__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__32628__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__32628__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__32643__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__32643__B (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__32646__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__32647__B (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__32652__A (.DIODE(net115));
 sky130_as_sc_hs__diode_2 ANTENNA__32652__B (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__32699__A (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__32699__B (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__32700__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__32700__B (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__32702__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__32702__B (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__32707__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__32707__B (.DIODE(net469));
 sky130_as_sc_hs__diode_2 ANTENNA__32708__A (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__32708__B (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__32724__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__32724__B (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__32725__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__32725__C (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__32726__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__32726__B (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__32727__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__32727__B (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__32759__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__32759__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__32760__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__32760__B (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__32765__A (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__32765__B (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__32766__A (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__32766__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__32795__A (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__32795__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__32796__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__32796__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__32810__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__32810__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__32811__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__32811__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__32816__A (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__32816__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__32817__A (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__32817__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__32832__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__32832__B (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__32835__B (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__32836__B (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__32841__A (.DIODE(net115));
 sky130_as_sc_hs__diode_2 ANTENNA__32841__B (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__32892__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__32892__B (.DIODE(_25035_));
 sky130_as_sc_hs__diode_2 ANTENNA__32893__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__32893__B (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__32900__A (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__32900__B (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__32901__A (.DIODE(net467));
 sky130_as_sc_hs__diode_2 ANTENNA__32901__B (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__32902__A (.DIODE(net469));
 sky130_as_sc_hs__diode_2 ANTENNA__32902__B (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__32917__A (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__32917__B (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__32918__A (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__32918__B (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__32919__A (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__32919__B (.DIODE(net453));
 sky130_as_sc_hs__diode_2 ANTENNA__32940__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__32940__B (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__32941__A (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__32941__B (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__32942__A (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__32942__B (.DIODE(net443));
 sky130_as_sc_hs__diode_2 ANTENNA__32953__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__32953__B (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__32954__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__32954__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__32955__A (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__32955__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__32981__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__32981__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__32982__A (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__32982__B (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__32983__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__32983__B (.DIODE(net435));
 sky130_as_sc_hs__diode_2 ANTENNA__33000__A (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__33000__B (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__33001__A (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__33001__B (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__33002__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__33002__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__33014__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__33018__A (.DIODE(net121));
 sky130_as_sc_hs__diode_2 ANTENNA__33018__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__33045__A (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__33045__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__33046__A (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA__33046__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__33049__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__33052__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__33053__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__33056__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__33059__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__33060__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__33063__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__33066__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__33067__A (.DIODE(net163));
 sky130_as_sc_hs__diode_2 ANTENNA__33070__A (.DIODE(net278));
 sky130_as_sc_hs__diode_2 ANTENNA__33073__A (.DIODE(net183));
 sky130_as_sc_hs__diode_2 ANTENNA__33074__A (.DIODE(net261));
 sky130_as_sc_hs__diode_2 ANTENNA__33075__A (.DIODE(net155));
 sky130_as_sc_hs__diode_2 ANTENNA__33076__A (.DIODE(net252));
 sky130_as_sc_hs__diode_2 ANTENNA__33077__A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA__33084__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__33091__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__33098__A (.DIODE(net159));
 sky130_as_sc_hs__diode_2 ANTENNA__33105__A (.DIODE(net258));
 sky130_as_sc_hs__diode_2 ANTENNA__33106__A (.DIODE(net152));
 sky130_as_sc_hs__diode_2 ANTENNA__33107__A (.DIODE(net249));
 sky130_as_sc_hs__diode_2 ANTENNA__33108__A (.DIODE(_19538_));
 sky130_as_sc_hs__diode_2 ANTENNA__33116__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__33116__B (.DIODE(net129));
 sky130_as_sc_hs__diode_2 ANTENNA__33139__A (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__33139__B (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__33146__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__33153__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__33156__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__33159__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__33160__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__33163__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__33167__A (.DIODE(net343));
 sky130_as_sc_hs__diode_2 ANTENNA__33168__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__33169__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__33170__A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__33173__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__33176__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__33177__A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA__33180__A (.DIODE(net211));
 sky130_as_sc_hs__diode_2 ANTENNA__33183__A (.DIODE(net351));
 sky130_as_sc_hs__diode_2 ANTENNA__33184__A (.DIODE(net343));
 sky130_as_sc_hs__diode_2 ANTENNA__33191__A (.DIODE(net231));
 sky130_as_sc_hs__diode_2 ANTENNA__33198__A (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__33199__A (.DIODE(net240));
 sky130_as_sc_hs__diode_2 ANTENNA__33200__A (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__33201__A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA__33210__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__33210__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__33211__B (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__33212__B (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__33213__A (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__33213__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__33266__A (.DIODE(net467));
 sky130_as_sc_hs__diode_2 ANTENNA__33266__B (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__33267__A (.DIODE(net469));
 sky130_as_sc_hs__diode_2 ANTENNA__33267__B (.DIODE(net455));
 sky130_as_sc_hs__diode_2 ANTENNA__33271__A (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__33271__B (.DIODE(net86));
 sky130_as_sc_hs__diode_2 ANTENNA__33275__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__33275__B (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__33276__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__33278__A (.DIODE(_23598_));
 sky130_as_sc_hs__diode_2 ANTENNA__33279__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__33279__B (.DIODE(_23598_));
 sky130_as_sc_hs__diode_2 ANTENNA__33297__A (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__33297__B (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__33298__A (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__33298__B (.DIODE(net453));
 sky130_as_sc_hs__diode_2 ANTENNA__33299__A (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__33299__B (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__33320__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__33320__B (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__33321__A (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__33321__B (.DIODE(net443));
 sky130_as_sc_hs__diode_2 ANTENNA__33322__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__33333__A (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__33333__B (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__33334__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__33334__B (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__33335__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__33335__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__33361__A (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__33361__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__33362__A (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__33362__B (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__33363__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__33363__B (.DIODE(net435));
 sky130_as_sc_hs__diode_2 ANTENNA__33385__A (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA__33385__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__33389__A (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__33389__B (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__33390__A (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__33390__B (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__33391__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__33391__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__33426__A (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__33426__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__33427__A (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__33427__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__33428__A (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__33428__B (.DIODE(net129));
 sky130_as_sc_hs__diode_2 ANTENNA__33451__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__33451__B (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__33453__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__33454__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__33454__B (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA__33455__B (.DIODE(_23643_));
 sky130_as_sc_hs__diode_2 ANTENNA__33456__B (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__33457__A (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__33457__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__33519__A (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__33519__B (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__33520__A (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__33520__B (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__33522__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__33522__B (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__33536__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__33536__B (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__33537__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__33537__C (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__33538__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__33539__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__33539__B (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__33570__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__33570__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__33571__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__33571__B (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__33576__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__33576__B (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__33577__A (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__33577__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__33608__A (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__33608__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__33609__A (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__33609__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__33623__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__33623__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__33624__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__33624__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__33629__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__33629__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__33630__A (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__33630__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__33643__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__33643__B (.DIODE(net443));
 sky130_as_sc_hs__diode_2 ANTENNA__33648__B (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__33649__B (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__33652__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__33652__B (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__33697__A (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__33697__B (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__33698__A (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__33698__B (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__33699__A (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__33701__A (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__33701__B (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__33717__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__33717__B (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__33718__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__33718__C (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__33719__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__33720__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__33720__B (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__33751__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__33751__B (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__33752__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__33752__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__33757__A (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__33757__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__33758__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__33758__B (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__33787__A (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__33787__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__33788__A (.DIODE(net453));
 sky130_as_sc_hs__diode_2 ANTENNA__33788__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__33802__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__33802__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__33803__A (.DIODE(net443));
 sky130_as_sc_hs__diode_2 ANTENNA__33803__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__33808__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__33808__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__33809__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__33809__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__33824__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__33824__B (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__33829__B (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__33830__B (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__33833__A (.DIODE(net115));
 sky130_as_sc_hs__diode_2 ANTENNA__33833__B (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__33880__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__33880__C (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__33883__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__33883__B (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__33899__A (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__33899__B (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__33900__A (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__33900__B (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__33920__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__33920__B (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__33921__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__33921__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__33928__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__33928__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__33929__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__33929__B (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__33958__A (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__33958__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__33959__A (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__33959__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__33973__A (.DIODE(net443));
 sky130_as_sc_hs__diode_2 ANTENNA__33973__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__33974__A (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__33974__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__33979__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__33979__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__33980__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__33980__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__33993__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__33993__B (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__33998__B (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__33999__B (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__34002__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__34002__B (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__34048__A (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__34048__C (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__34051__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__34051__B (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__34076__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__34076__B (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__34077__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__34082__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__34082__B (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__34083__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__34083__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__34113__A (.DIODE(net455));
 sky130_as_sc_hs__diode_2 ANTENNA__34113__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__34114__A (.DIODE(net453));
 sky130_as_sc_hs__diode_2 ANTENNA__34114__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__34128__A (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__34128__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__34129__A (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__34129__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__34134__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__34134__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__34135__C (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__34136__A (.DIODE(net443));
 sky130_as_sc_hs__diode_2 ANTENNA__34136__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__34146__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__34146__B (.DIODE(net453));
 sky130_as_sc_hs__diode_2 ANTENNA__34151__B (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__34152__B (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__34155__A (.DIODE(net115));
 sky130_as_sc_hs__diode_2 ANTENNA__34155__B (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__34206__A (.DIODE(net116));
 sky130_as_sc_hs__diode_2 ANTENNA__34206__B (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__34207__B (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__34208__B (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__34210__B (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__34211__B (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__34221__B (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__34222__B (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__34227__A (.DIODE(net116));
 sky130_as_sc_hs__diode_2 ANTENNA__34227__B (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__34239__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__34239__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__34240__A (.DIODE(net455));
 sky130_as_sc_hs__diode_2 ANTENNA__34240__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__34244__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__34244__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__34245__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__34245__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__34249__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__34249__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__34250__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__34250__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__34258__A (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__34258__B (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__34259__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__34259__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__34263__A (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__34263__B (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__34264__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__34264__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__34266__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__34266__B (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__34267__A (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__34267__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__34279__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__34279__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__34280__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__34280__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__34284__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__34284__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__34285__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__34285__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__34299__A (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__34299__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__34300__A (.DIODE(net86));
 sky130_as_sc_hs__diode_2 ANTENNA__34300__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__34305__A (.DIODE(net86));
 sky130_as_sc_hs__diode_2 ANTENNA__34305__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__34306__A (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__34306__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__34313__A (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__34313__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__34314__A (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__34314__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__34334__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__34334__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__34335__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__34335__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__34340__A (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__34340__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__34341__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__34341__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__34364__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__34364__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__34365__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__34365__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__34379__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__34379__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__34380__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__34380__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__34387__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__34387__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__34388__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__34388__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__34405__B (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__34406__B (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__34409__A (.DIODE(net116));
 sky130_as_sc_hs__diode_2 ANTENNA__34409__B (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__34424__A (.DIODE(net455));
 sky130_as_sc_hs__diode_2 ANTENNA__34424__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__34425__A (.DIODE(net86));
 sky130_as_sc_hs__diode_2 ANTENNA__34425__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__34429__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__34429__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__34430__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__34430__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__34440__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__34440__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__34441__A (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__34441__B (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__34444__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__34444__B (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__34445__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__34445__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__34465__A (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__34465__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__34466__A (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__34466__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__34488__A (.DIODE(net116));
 sky130_as_sc_hs__diode_2 ANTENNA__34488__B (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__34489__B (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__34490__B (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__34519__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__34519__B (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__34520__A (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__34520__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__34521__A (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__34521__B (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__34529__A (.DIODE(net86));
 sky130_as_sc_hs__diode_2 ANTENNA__34529__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__34530__A (.DIODE(net453));
 sky130_as_sc_hs__diode_2 ANTENNA__34530__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__34534__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__34534__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__34535__A (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__34535__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__34545__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__34545__B (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__34546__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__34546__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__34569__A (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__34569__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__34570__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__34570__B (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__34574__A (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__34575__A (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__34575__B (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__34618__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__34618__B (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__34642__A (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__34642__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__34643__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__34643__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__34657__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__34657__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__34658__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__34658__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__34663__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__34663__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__34664__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__34664__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__34681__B (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__34682__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__34685__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__34685__B (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__34719__A (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__34719__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__34735__A (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__34735__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__34736__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__34736__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__34750__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__34750__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__34751__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__34751__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__34756__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__34756__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__34757__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__34757__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__34772__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__34772__B (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__34810__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__34810__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__34826__A (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__34826__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__34827__A (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__34827__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__34841__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__34841__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__34842__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__34842__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__34847__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__34847__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__34848__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__34848__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__34859__B (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__34860__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__34860__B (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__34913__A (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__34913__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__34914__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__34914__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__34919__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__34919__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__34920__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__34920__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__34931__B (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__34932__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__34932__B (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__34971__A (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__34971__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__34980__A (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__34980__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__34981__A (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__34981__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__34986__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__34986__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__34987__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__34987__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__34998__B (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__34999__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__34999__B (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__35017__B (.DIODE(_04288_));
 sky130_as_sc_hs__diode_2 ANTENNA__35038__A (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__35038__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__35049__A (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__35049__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__35050__A (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__35050__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__35054__A (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__35054__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__35055__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__35055__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__35065__A (.DIODE(net112));
 sky130_as_sc_hs__diode_2 ANTENNA__35066__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__35066__B (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__35103__A (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__35103__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__35104__A (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__35104__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__35138__A (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__35138__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__35139__A (.DIODE(net459));
 sky130_as_sc_hs__diode_2 ANTENNA__35139__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__35152__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__35152__B (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__35181__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__35181__B (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__35225__A (.DIODE(net116));
 sky130_as_sc_hs__diode_2 ANTENNA__35225__B (.DIODE(net91));
 sky130_as_sc_hs__diode_2 ANTENNA__35292__A (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__35292__C (.DIODE(_24536_));
 sky130_as_sc_hs__diode_2 ANTENNA__35295__A (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__35295__B (.DIODE(net87));
 sky130_as_sc_hs__diode_2 ANTENNA__35320__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__35320__B (.DIODE(net448));
 sky130_as_sc_hs__diode_2 ANTENNA__35321__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__35321__B (.DIODE(net450));
 sky130_as_sc_hs__diode_2 ANTENNA__35326__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__35326__B (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__35327__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__35327__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__35357__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__35357__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__35358__A (.DIODE(net86));
 sky130_as_sc_hs__diode_2 ANTENNA__35358__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__35372__A (.DIODE(net453));
 sky130_as_sc_hs__diode_2 ANTENNA__35372__B (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__35373__A (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__35373__B (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__35378__A (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__35378__B (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__35379__A (.DIODE(net443));
 sky130_as_sc_hs__diode_2 ANTENNA__35379__B (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__35390__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__35390__B (.DIODE(net86));
 sky130_as_sc_hs__diode_2 ANTENNA__35395__B (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__35396__B (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__35399__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__35399__B (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__35446__A (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__35446__B (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__35524__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__35524__B (.DIODE(net455));
 sky130_as_sc_hs__diode_2 ANTENNA__35529__B (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__35530__B (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__35533__A (.DIODE(net114));
 sky130_as_sc_hs__diode_2 ANTENNA__35533__B (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__35628__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__35628__B (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__35634__A (.DIODE(net116));
 sky130_as_sc_hs__diode_2 ANTENNA__35634__B (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__35702__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__35702__B (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__35856__B (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__35857__B (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__35858__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__35858__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__35873__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__35873__B (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__35886__A (.DIODE(_25205_));
 sky130_as_sc_hs__diode_2 ANTENNA__35886__B (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA__35922__A (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__35922__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__35926__A (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__35926__B (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__35927__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__35927__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__35931__A (.DIODE(net121));
 sky130_as_sc_hs__diode_2 ANTENNA__35931__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__35944__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__35944__B (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__35945__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__35945__B (.DIODE(net435));
 sky130_as_sc_hs__diode_2 ANTENNA__35949__A (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__35949__B (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__35974__A (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__35974__B (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__35975__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__35975__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__35979__A (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__35979__B (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__35983__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__35983__B (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__35984__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__35984__B (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__35988__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__35988__B (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__36007__A (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__36007__B (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__36008__A (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__36008__B (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__36012__A (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__36012__B (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__36022__A (.DIODE(net467));
 sky130_as_sc_hs__diode_2 ANTENNA__36022__B (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__36023__A (.DIODE(net469));
 sky130_as_sc_hs__diode_2 ANTENNA__36023__B (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__36027__A (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__36027__B (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__36031__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__36031__B (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__36032__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__36033__A (.DIODE(_23598_));
 sky130_as_sc_hs__diode_2 ANTENNA__36033__B (.DIODE(net458));
 sky130_as_sc_hs__diode_2 ANTENNA__36094__A (.DIODE(_05123_));
 sky130_as_sc_hs__diode_2 ANTENNA__36125__A (.DIODE(net116));
 sky130_as_sc_hs__diode_2 ANTENNA__36125__B (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__36185__B (.DIODE(_05456_));
 sky130_as_sc_hs__diode_2 ANTENNA__36237__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__36239__C (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__36240__A (.DIODE(\tholin_riscv.Jimm[13] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36243__A (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__36243__B (.DIODE(net417));
 sky130_as_sc_hs__diode_2 ANTENNA__36244__A (.DIODE(_23598_));
 sky130_as_sc_hs__diode_2 ANTENNA__36259__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36268__B (.DIODE(_05518_));
 sky130_as_sc_hs__diode_2 ANTENNA__36297__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36303__A (.DIODE(_24337_));
 sky130_as_sc_hs__diode_2 ANTENNA__36306__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36312__B (.DIODE(net417));
 sky130_as_sc_hs__diode_2 ANTENNA__36315__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__36330__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__36331__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36336__A (.DIODE(_05606_));
 sky130_as_sc_hs__diode_2 ANTENNA__36338__B (.DIODE(net417));
 sky130_as_sc_hs__diode_2 ANTENNA__36340__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36341__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36348__B (.DIODE(net417));
 sky130_as_sc_hs__diode_2 ANTENNA__36350__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36351__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36360__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__36361__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36370__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36371__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36380__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36381__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36389__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__36390__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36395__A (.DIODE(_20707_));
 sky130_as_sc_hs__diode_2 ANTENNA__36399__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__36405__A (.DIODE(_20622_));
 sky130_as_sc_hs__diode_2 ANTENNA__36419__B (.DIODE(_05518_));
 sky130_as_sc_hs__diode_2 ANTENNA__36429__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36447__A (.DIODE(\tholin_riscv.Bimm[10] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36447__B (.DIODE(net417));
 sky130_as_sc_hs__diode_2 ANTENNA__36458__A (.DIODE(\tholin_riscv.Bimm[9] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36458__B (.DIODE(net417));
 sky130_as_sc_hs__diode_2 ANTENNA__36470__B (.DIODE(net417));
 sky130_as_sc_hs__diode_2 ANTENNA__36475__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__36476__A (.DIODE(_22301_));
 sky130_as_sc_hs__diode_2 ANTENNA__36478__B (.DIODE(net417));
 sky130_as_sc_hs__diode_2 ANTENNA__36479__B (.DIODE(net417));
 sky130_as_sc_hs__diode_2 ANTENNA__36517__A (.DIODE(\tholin_riscv.Bimm[4] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36524__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__36525__A (.DIODE(_21977_));
 sky130_as_sc_hs__diode_2 ANTENNA__36531__A (.DIODE(\tholin_riscv.Bimm[3] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36543__A (.DIODE(\tholin_riscv.Iimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36546__A (.DIODE(\tholin_riscv.Bimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36553__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__36554__B (.DIODE(net126));
 sky130_as_sc_hs__diode_2 ANTENNA__36559__B (.DIODE(\tholin_riscv.Bimm[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36565__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__36566__A (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__36570__A (.DIODE(\tholin_riscv.Iimm[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36573__A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36652__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__36659__A (.DIODE(\tholin_riscv.Bimm[10] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36666__B (.DIODE(_21036_));
 sky130_as_sc_hs__diode_2 ANTENNA__36667__A (.DIODE(\tholin_riscv.Iimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36671__B (.DIODE(_20931_));
 sky130_as_sc_hs__diode_2 ANTENNA__36672__A (.DIODE(\tholin_riscv.Iimm[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36675__B (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__36676__B (.DIODE(net116));
 sky130_as_sc_hs__diode_2 ANTENNA__36677__A (.DIODE(\tholin_riscv.Iimm[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36694__A (.DIODE(_05926_));
 sky130_as_sc_hs__diode_2 ANTENNA__36695__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__36734__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__36738__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__36758__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__36779__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__36806__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__36870__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__36877__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__36893__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__36894__A (.DIODE(\tholin_riscv.Jimm[13] ));
 sky130_as_sc_hs__diode_2 ANTENNA__36897__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__36915__B (.DIODE(net121));
 sky130_as_sc_hs__diode_2 ANTENNA__36916__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__36916__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__36920__B (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__36931__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__36931__B (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__36939__A (.DIODE(_25211_));
 sky130_as_sc_hs__diode_2 ANTENNA__36939__B (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA__36940__A (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__36940__B (.DIODE(net129));
 sky130_as_sc_hs__diode_2 ANTENNA__36972__A (.DIODE(net455));
 sky130_as_sc_hs__diode_2 ANTENNA__36976__A (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__36976__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__36980__A (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__36980__B (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__36981__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__36981__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__36985__A (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA__36985__B (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__36998__A (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__36998__B (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__36999__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__36999__B (.DIODE(net435));
 sky130_as_sc_hs__diode_2 ANTENNA__37003__A (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__37003__B (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__37028__A (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__37028__B (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__37029__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__37029__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__37033__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__37033__B (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__37037__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__37037__B (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__37038__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__37038__B (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__37042__A (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__37042__B (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__37061__A (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__37061__B (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__37062__A (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__37062__B (.DIODE(net443));
 sky130_as_sc_hs__diode_2 ANTENNA__37066__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__37066__B (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__37076__A (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__37076__B (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__37077__A (.DIODE(net467));
 sky130_as_sc_hs__diode_2 ANTENNA__37077__B (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__37078__A (.DIODE(net469));
 sky130_as_sc_hs__diode_2 ANTENNA__37078__B (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__37085__A (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__37085__B (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__37086__A (.DIODE(_23598_));
 sky130_as_sc_hs__diode_2 ANTENNA__37086__B (.DIODE(net90));
 sky130_as_sc_hs__diode_2 ANTENNA__37087__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__37154__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__37178__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__37182__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__37190__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__37199__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__37213__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__37225__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__37233__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__37249__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__37251__A (.DIODE(_05968_));
 sky130_as_sc_hs__diode_2 ANTENNA__37256__B (.DIODE(\tholin_riscv.Bimm[10] ));
 sky130_as_sc_hs__diode_2 ANTENNA__37261__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__37266__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__37273__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__37275__A (.DIODE(_23598_));
 sky130_as_sc_hs__diode_2 ANTENNA__37277__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__37281__B (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__37288__B (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__37292__C (.DIODE(net109));
 sky130_as_sc_hs__diode_2 ANTENNA__37298__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__37307__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__37317__A (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA__37318__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__37318__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__37322__B (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__37333__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__37333__B (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__37340__A (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__37340__B (.DIODE(net129));
 sky130_as_sc_hs__diode_2 ANTENNA__37368__A (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__37368__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__37369__A (.DIODE(net86));
 sky130_as_sc_hs__diode_2 ANTENNA__37369__B (.DIODE(net437));
 sky130_as_sc_hs__diode_2 ANTENNA__37373__A (.DIODE(_24808_));
 sky130_as_sc_hs__diode_2 ANTENNA__37373__B (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA__37377__A (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__37377__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__37378__C (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__37395__A (.DIODE(net445));
 sky130_as_sc_hs__diode_2 ANTENNA__37395__B (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__37396__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__37396__B (.DIODE(net435));
 sky130_as_sc_hs__diode_2 ANTENNA__37400__A (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__37400__B (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__37425__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__37425__B (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__37426__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__37426__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__37430__A (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__37430__B (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__37434__A (.DIODE(net477));
 sky130_as_sc_hs__diode_2 ANTENNA__37434__B (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__37435__A (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__37435__B (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__37439__B (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__37458__A (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__37458__B (.DIODE(net443));
 sky130_as_sc_hs__diode_2 ANTENNA__37459__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__37459__B (.DIODE(net462));
 sky130_as_sc_hs__diode_2 ANTENNA__37463__B (.DIODE(net461));
 sky130_as_sc_hs__diode_2 ANTENNA__37473__A (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__37473__B (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__37474__A (.DIODE(net467));
 sky130_as_sc_hs__diode_2 ANTENNA__37474__B (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__37475__A (.DIODE(net469));
 sky130_as_sc_hs__diode_2 ANTENNA__37475__B (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__37482__A (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__37482__B (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__37483__A (.DIODE(_23598_));
 sky130_as_sc_hs__diode_2 ANTENNA__37483__B (.DIODE(_24053_));
 sky130_as_sc_hs__diode_2 ANTENNA__37484__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__37557__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__37559__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__37567__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__37569__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__37570__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__37575__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__37582__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__37594__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__37595__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__37606__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__37611__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__37614__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__37617__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__37620__A (.DIODE(net109));
 sky130_as_sc_hs__diode_2 ANTENNA__37624__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__37631__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__37634__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__37647__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__37648__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__37659__B (.DIODE(_25874_));
 sky130_as_sc_hs__diode_2 ANTENNA__37660__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__37660__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__37664__B (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__37675__A (.DIODE(net121));
 sky130_as_sc_hs__diode_2 ANTENNA__37675__B (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__37682__A (.DIODE(_24216_));
 sky130_as_sc_hs__diode_2 ANTENNA__37682__B (.DIODE(net129));
 sky130_as_sc_hs__diode_2 ANTENNA__37707__A (.DIODE(_24814_));
 sky130_as_sc_hs__diode_2 ANTENNA__37707__B (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA__37708__A (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__37708__B (.DIODE(net437));
 sky130_as_sc_hs__diode_2 ANTENNA__37712__A (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA__37712__B (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__37713__A (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__37713__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__37717__A (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__37717__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__37730__A (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__37730__B (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__37731__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__37731__B (.DIODE(net435));
 sky130_as_sc_hs__diode_2 ANTENNA__37735__A (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__37735__B (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__37760__B (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__37761__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__37761__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__37765__A (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__37765__B (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__37769__A (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__37769__B (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__37770__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__37770__B (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__37774__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__37774__B (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__37793__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__37793__B (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__37794__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__37794__B (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__37798__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__37798__B (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__37808__A (.DIODE(net467));
 sky130_as_sc_hs__diode_2 ANTENNA__37808__B (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__37809__A (.DIODE(net469));
 sky130_as_sc_hs__diode_2 ANTENNA__37809__B (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__37813__A (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__37813__B (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__37817__A (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__37817__B (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__37818__A (.DIODE(_23598_));
 sky130_as_sc_hs__diode_2 ANTENNA__37818__B (.DIODE(_23712_));
 sky130_as_sc_hs__diode_2 ANTENNA__37819__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__37887__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__37890__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__37893__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__37903__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__37908__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__37911__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__37912__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__37914__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__37917__A (.DIODE(net109));
 sky130_as_sc_hs__diode_2 ANTENNA__37921__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__37934__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__37936__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__37937__A (.DIODE(net82));
 sky130_as_sc_hs__diode_2 ANTENNA__37942__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__37949__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__37961__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__37962__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__37981__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__37982__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__37993__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__37994__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__37994__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__37998__B (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__38009__A (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA__38009__B (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__38014__A (.DIODE(_24229_));
 sky130_as_sc_hs__diode_2 ANTENNA__38014__B (.DIODE(net129));
 sky130_as_sc_hs__diode_2 ANTENNA__38039__A (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__38039__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__38040__A (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__38040__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__38044__A (.DIODE(_24768_));
 sky130_as_sc_hs__diode_2 ANTENNA__38044__B (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA__38052__A (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA__38052__B (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__38058__A (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__38058__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__38059__A (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__38059__B (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__38063__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__38063__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__38088__A (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__38088__B (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__38089__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__38089__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__38093__A (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__38093__B (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__38097__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__38097__B (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__38098__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__38098__B (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__38102__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__38102__B (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__38121__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__38121__B (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__38122__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__38122__B (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__38126__A (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__38126__B (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__38136__A (.DIODE(net467));
 sky130_as_sc_hs__diode_2 ANTENNA__38136__B (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__38137__A (.DIODE(net469));
 sky130_as_sc_hs__diode_2 ANTENNA__38137__B (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__38141__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__38141__B (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__38145__A (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__38145__B (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__38223__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__38226__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__38229__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__38239__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__38242__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__38246__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__38251__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__38253__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__38261__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__38266__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__38269__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__38270__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__38272__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__38275__A (.DIODE(net109));
 sky130_as_sc_hs__diode_2 ANTENNA__38279__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__38292__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__38293__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__38302__B (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA__38303__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__38303__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__38307__B (.DIODE(net121));
 sky130_as_sc_hs__diode_2 ANTENNA__38318__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__38318__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__38323__A (.DIODE(_24256_));
 sky130_as_sc_hs__diode_2 ANTENNA__38323__B (.DIODE(net129));
 sky130_as_sc_hs__diode_2 ANTENNA__38345__A (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__38345__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__38346__A (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__38346__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__38354__A (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__38354__B (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__38360__A (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__38360__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__38361__A (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__38361__B (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__38365__A (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA__38365__B (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__38390__A (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__38390__B (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__38391__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__38391__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__38395__A (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__38395__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__38399__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__38399__B (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__38400__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__38400__B (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__38404__A (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__38404__B (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__38423__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__38423__B (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__38424__A (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__38424__B (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__38428__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__38428__B (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__38438__A (.DIODE(net467));
 sky130_as_sc_hs__diode_2 ANTENNA__38438__B (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__38439__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__38439__B (.DIODE(net469));
 sky130_as_sc_hs__diode_2 ANTENNA__38443__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__38443__B (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__38447__A (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__38447__B (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__38516__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__38522__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__38532__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__38535__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__38539__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__38544__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__38546__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__38554__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__38556__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__38559__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__38563__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__38565__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__38568__A (.DIODE(net109));
 sky130_as_sc_hs__diode_2 ANTENNA__38572__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__38584__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__38585__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__38595__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__38595__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__38596__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__38596__B (.DIODE(_23624_));
 sky130_as_sc_hs__diode_2 ANTENNA__38608__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__38608__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__38613__A (.DIODE(_24501_));
 sky130_as_sc_hs__diode_2 ANTENNA__38613__B (.DIODE(net129));
 sky130_as_sc_hs__diode_2 ANTENNA__38632__A (.DIODE(_24774_));
 sky130_as_sc_hs__diode_2 ANTENNA__38632__B (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA__38633__A (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__38633__B (.DIODE(net441));
 sky130_as_sc_hs__diode_2 ANTENNA__38640__A (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__38640__B (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__38651__A (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__38651__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__38676__A (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__38676__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__38677__A (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__38677__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__38681__A (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__38681__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__38685__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__38685__B (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__38686__A (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__38686__B (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__38690__A (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__38690__B (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__38709__A (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__38709__B (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__38710__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__38710__B (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__38714__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__38714__B (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__38724__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__38724__B (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__38725__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__38725__B (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__38729__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__38729__B (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__38733__A (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__38733__B (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__38809__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__38810__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__38813__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__38823__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__38826__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__38830__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__38835__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__38837__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__38845__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__38847__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__38850__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__38854__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__38856__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__38859__A (.DIODE(net109));
 sky130_as_sc_hs__diode_2 ANTENNA__38863__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__38876__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__38877__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__38888__A (.DIODE(_23702_));
 sky130_as_sc_hs__diode_2 ANTENNA__38888__B (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA__38889__A (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__38889__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__38890__A (.DIODE(_23624_));
 sky130_as_sc_hs__diode_2 ANTENNA__38890__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__38902__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__38902__B (.DIODE(net129));
 sky130_as_sc_hs__diode_2 ANTENNA__38922__A (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__38924__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__38924__B (.DIODE(net437));
 sky130_as_sc_hs__diode_2 ANTENNA__38930__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__38930__B (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__38931__A (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__38931__B (.DIODE(net435));
 sky130_as_sc_hs__diode_2 ANTENNA__38935__A (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__38935__B (.DIODE(_02481_));
 sky130_as_sc_hs__diode_2 ANTENNA__38960__A (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__38960__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__38961__A (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__38961__B (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__38965__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__38965__B (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__38969__A (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__38969__B (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__38970__A (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__38970__B (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__38974__A (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__38974__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__38993__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__38993__B (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__38994__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__38994__B (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__38998__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__38998__B (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__39008__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__39008__B (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__39009__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__39009__B (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__39013__A (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__39013__B (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__39017__A (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__39017__B (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__39088__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__39089__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__39092__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__39102__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__39110__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__39114__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__39119__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__39121__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__39124__A (.DIODE(_05968_));
 sky130_as_sc_hs__diode_2 ANTENNA__39126__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__39129__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__39133__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__39135__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__39142__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__39155__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__39156__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__39173__A (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__39173__B (.DIODE(net129));
 sky130_as_sc_hs__diode_2 ANTENNA__39180__A (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__39180__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__39181__A (.DIODE(_23624_));
 sky130_as_sc_hs__diode_2 ANTENNA__39181__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__39201__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__39201__B (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__39202__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__39202__B (.DIODE(net437));
 sky130_as_sc_hs__diode_2 ANTENNA__39208__A (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__39208__B (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__39209__A (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA__39209__B (.DIODE(net435));
 sky130_as_sc_hs__diode_2 ANTENNA__39213__A (.DIODE(_24729_));
 sky130_as_sc_hs__diode_2 ANTENNA__39213__B (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA__39238__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__39238__B (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__39239__A (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__39239__B (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__39243__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__39243__B (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__39247__A (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__39247__B (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__39248__A (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__39248__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__39252__A (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__39252__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__39271__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__39271__B (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__39272__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__39272__B (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__39276__A (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__39276__B (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__39286__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__39286__B (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__39287__A (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__39287__B (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__39291__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__39291__B (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__39295__A (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__39295__B (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__39296__A (.DIODE(_24545_));
 sky130_as_sc_hs__diode_2 ANTENNA__39296__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__39297__A (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__39297__B (.DIODE(_25035_));
 sky130_as_sc_hs__diode_2 ANTENNA__39372__A (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__39378__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__39381__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__39391__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__39395__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__39397__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__39400__A (.DIODE(_05968_));
 sky130_as_sc_hs__diode_2 ANTENNA__39402__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__39405__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__39409__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__39411__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__39418__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__39431__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__39432__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__39442__A (.DIODE(net85));
 sky130_as_sc_hs__diode_2 ANTENNA__39442__B (.DIODE(net129));
 sky130_as_sc_hs__diode_2 ANTENNA__39449__A (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__39449__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__39450__A (.DIODE(_23624_));
 sky130_as_sc_hs__diode_2 ANTENNA__39450__B (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA__39470__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__39470__B (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__39471__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__39471__B (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__39477__A (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__39477__B (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__39478__A (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__39478__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__39508__A (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__39508__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__39512__A (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__39512__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__39513__A (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__39513__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__39517__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__39517__B (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__39536__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__39536__B (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__39537__A (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__39537__B (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__39541__A (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__39541__B (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__39551__A (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__39551__B (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__39552__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__39552__B (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__39556__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__39556__B (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__39560__A (.DIODE(net454));
 sky130_as_sc_hs__diode_2 ANTENNA__39560__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__39561__A (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__39561__B (.DIODE(_25035_));
 sky130_as_sc_hs__diode_2 ANTENNA__39565__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__39565__B (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__39627__A (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__39630__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__39631__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__39634__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__39646__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__39647__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__39648__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__39653__A (.DIODE(_05926_));
 sky130_as_sc_hs__diode_2 ANTENNA__39655__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__39658__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__39663__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__39667__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__39671__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__39683__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__39684__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__39695__A (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__39702__A (.DIODE(net452));
 sky130_as_sc_hs__diode_2 ANTENNA__39702__B (.DIODE(net129));
 sky130_as_sc_hs__diode_2 ANTENNA__39720__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__39720__B (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__39721__A (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__39721__B (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__39726__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__39726__B (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__39727__A (.DIODE(net444));
 sky130_as_sc_hs__diode_2 ANTENNA__39727__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__39752__A (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__39752__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__39753__A (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__39753__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__39757__A (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__39757__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__39766__A (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA__39766__B (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__39785__A (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__39785__B (.DIODE(net84));
 sky130_as_sc_hs__diode_2 ANTENNA__39786__A (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__39786__B (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__39790__A (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__39790__B (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__39801__C (.DIODE(_25035_));
 sky130_as_sc_hs__diode_2 ANTENNA__39805__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__39805__B (.DIODE(_24479_));
 sky130_as_sc_hs__diode_2 ANTENNA__39813__A (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA__39813__B (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__39814__A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA__39814__B (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__39818__A (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__39818__B (.DIODE(net470));
 sky130_as_sc_hs__diode_2 ANTENNA__39885__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__39886__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__39889__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__39899__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__39902__A (.DIODE(_05926_));
 sky130_as_sc_hs__diode_2 ANTENNA__39903__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__39905__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__39906__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__39910__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__39914__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__39917__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__39919__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__39926__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__39938__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__39939__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__39954__A (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__39954__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__39972__A (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__39972__B (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__39973__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__39973__B (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__39977__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__39977__B (.DIODE(net435));
 sky130_as_sc_hs__diode_2 ANTENNA__40000__A (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__40000__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__40001__A (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__40001__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__40005__A (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA__40005__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__40014__A (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__40014__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__40036__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__40036__B (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__40044__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__40044__B (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__40045__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__40045__B (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__40049__A (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__40049__B (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__40062__A (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__40062__B (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__40063__A (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__40063__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__40067__A (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__40067__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__40123__A (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__40127__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__40143__A (.DIODE(_05926_));
 sky130_as_sc_hs__diode_2 ANTENNA__40144__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__40146__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__40147__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__40151__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__40153__A (.DIODE(_05714_));
 sky130_as_sc_hs__diode_2 ANTENNA__40155__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__40158__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__40160__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__40167__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__40179__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__40180__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__40190__A (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__40190__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__40197__A (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__40197__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__40209__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__40209__B (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__40210__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__40210__B (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__40214__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__40214__B (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__40232__A (.DIODE(net446));
 sky130_as_sc_hs__diode_2 ANTENNA__40232__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__40233__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__40233__B (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__40237__A (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__40237__B (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__40245__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__40245__B (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__40246__A (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__40246__B (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__40250__A (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__40250__B (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__40263__A (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__40263__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__40264__A (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__40264__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__40268__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__40268__B (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__40287__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__40287__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__40288__A (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA__40288__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__40292__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__40292__B (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__40293__A (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__40293__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__40297__A (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__40297__B (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__40361__A (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__40365__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__40366__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__40369__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__40378__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__40379__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__40381__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__40382__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__40387__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__40389__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__40392__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__40397__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__40401__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__40404__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__40417__A (.DIODE(\tholin_riscv.Jimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__40420__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__40421__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__40440__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__40440__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__40450__A (.DIODE(net78));
 sky130_as_sc_hs__diode_2 ANTENNA__40450__B (.DIODE(_02550_));
 sky130_as_sc_hs__diode_2 ANTENNA__40451__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__40451__B (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__40455__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__40455__B (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__40468__A (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__40468__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__40481__A (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__40481__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__40482__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__40482__B (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__40486__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__40486__B (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__40505__A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA__40505__B (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA__40506__A (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__40506__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__40507__A (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__40507__B (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__40511__A (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA__40511__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__40537__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__40537__B (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__40538__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__40538__B (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__40601__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__40602__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__40604__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__40605__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__40610__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__40612__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__40615__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__40617__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__40624__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__40627__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__40640__B (.DIODE(\tholin_riscv.Jimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__40642__B (.DIODE(\tholin_riscv.Jimm[13] ));
 sky130_as_sc_hs__diode_2 ANTENNA__40646__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__40647__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__40649__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__40657__A (.DIODE(net442));
 sky130_as_sc_hs__diode_2 ANTENNA__40657__B (.DIODE(_02550_));
 sky130_as_sc_hs__diode_2 ANTENNA__40658__A (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__40658__B (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__40662__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__40662__B (.DIODE(net456));
 sky130_as_sc_hs__diode_2 ANTENNA__40670__A (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__40670__B (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__40671__A (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__40671__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__40675__A (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__40675__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__40688__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__40688__B (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__40689__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__40689__B (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__40693__A (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__40693__B (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA__40712__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__40712__B (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__40713__A (.DIODE(_24527_));
 sky130_as_sc_hs__diode_2 ANTENNA__40713__B (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__40714__A (.DIODE(net89));
 sky130_as_sc_hs__diode_2 ANTENNA__40714__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__40740__A (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA__40740__B (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__40741__A (.DIODE(net437));
 sky130_as_sc_hs__diode_2 ANTENNA__40741__B (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__40745__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__40745__B (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__40767__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__40767__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__40774__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__40774__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__40816__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__40828__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__40829__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__40831__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__40832__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__40837__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__40839__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__40844__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__40847__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__40851__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__40854__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__40866__A (.DIODE(\tholin_riscv.Jimm[14] ));
 sky130_as_sc_hs__diode_2 ANTENNA__40869__B (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__40873__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__40876__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__40884__A (.DIODE(_23674_));
 sky130_as_sc_hs__diode_2 ANTENNA__40884__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__40885__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__40885__B (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__40889__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__40889__B (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__40897__A (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__40897__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__40898__A (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__40898__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__40902__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__40902__B (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__40915__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__40915__B (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__40916__A (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__40916__B (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__40920__A (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__40920__B (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__40939__A (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__40939__B (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__40960__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__40960__B (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__40961__A (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__40961__B (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__40962__A (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__40962__B (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__40984__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__40984__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__40991__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__40991__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__41029__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__41032__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__41041__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__41042__A (.DIODE(_05935_));
 sky130_as_sc_hs__diode_2 ANTENNA__41044__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__41045__A (.DIODE(_05929_));
 sky130_as_sc_hs__diode_2 ANTENNA__41050__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__41052__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__41055__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__41057__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__41064__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__41067__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__41083__B (.DIODE(net373));
 sky130_as_sc_hs__diode_2 ANTENNA__41087__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__41090__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__41097__A (.DIODE(net360));
 sky130_as_sc_hs__diode_2 ANTENNA__41097__B (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__41105__A (.DIODE(_05123_));
 sky130_as_sc_hs__diode_2 ANTENNA__41114__A (.DIODE(net480));
 sky130_as_sc_hs__diode_2 ANTENNA__41114__B (.DIODE(_02550_));
 sky130_as_sc_hs__diode_2 ANTENNA__41115__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__41115__B (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__41119__A (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__41119__B (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__41127__A (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__41127__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__41128__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__41128__B (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__41132__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__41132__B (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__41145__A (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__41145__B (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__41146__A (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA__41146__B (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__41150__A (.DIODE(net460));
 sky130_as_sc_hs__diode_2 ANTENNA__41150__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__41168__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__41168__B (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__41184__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__41184__B (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__41185__A (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__41185__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__41186__A (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__41186__B (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__41208__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__41208__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__41215__A (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__41215__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__41248__A (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__41252__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__41264__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__41266__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__41268__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__41273__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__41276__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__41280__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__41283__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__41303__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__41306__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__41311__A (.DIODE(net347));
 sky130_as_sc_hs__diode_2 ANTENNA__41311__B (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__41315__A (.DIODE(net476));
 sky130_as_sc_hs__diode_2 ANTENNA__41315__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__41316__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__41316__B (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__41320__A (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__41320__B (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__41328__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__41328__B (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__41329__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__41329__B (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__41333__A (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__41333__B (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__41346__A (.DIODE(net464));
 sky130_as_sc_hs__diode_2 ANTENNA__41346__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__41364__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__41364__B (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__41377__A (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__41377__B (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__41378__A (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__41378__B (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__41379__A (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__41379__B (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__41401__A (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA__41401__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__41408__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__41408__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__41446__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__41456__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__41458__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__41460__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__41463__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__41465__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__41472__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__41475__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__41491__B (.DIODE(net342));
 sky130_as_sc_hs__diode_2 ANTENNA__41495__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__41498__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__41503__A (.DIODE(net340));
 sky130_as_sc_hs__diode_2 ANTENNA__41503__B (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__41506__A (.DIODE(net438));
 sky130_as_sc_hs__diode_2 ANTENNA__41506__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__41507__A (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__41507__B (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__41511__A (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__41511__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__41519__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__41519__B (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__41520__A (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__41520__B (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__41524__A (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__41524__B (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__41536__A (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA__41536__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__41548__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__41548__B (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__41560__A (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__41560__B (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__41561__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__41561__B (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__41562__A (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__41562__B (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__41584__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__41584__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__41591__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__41591__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__41628__A (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__41633__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__41647__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__41649__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__41651__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__41654__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__41656__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__41662__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__41666__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__41669__C (.DIODE(_10922_));
 sky130_as_sc_hs__diode_2 ANTENNA__41682__B (.DIODE(net337));
 sky130_as_sc_hs__diode_2 ANTENNA__41686__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__41689__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__41694__A (.DIODE(net335));
 sky130_as_sc_hs__diode_2 ANTENNA__41694__B (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__41698__A (.DIODE(net472));
 sky130_as_sc_hs__diode_2 ANTENNA__41698__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__41699__A (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__41699__B (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__41703__A (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__41703__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__41711__A (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__41711__B (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__41712__A (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__41712__B (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__41716__A (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA__41716__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__41735__A (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__41735__B (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__41748__A (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__41748__B (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__41749__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__41749__B (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__41750__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__41750__B (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__41772__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__41772__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__41779__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__41779__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__41811__A (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__41815__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__41816__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__41828__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__41830__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__41832__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__41837__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__41840__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__41843__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__41847__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__41863__B (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA__41867__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__41869__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__41871__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__41876__A (.DIODE(\tholin_riscv.Iimm[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__41876__B (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__41885__A (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__41885__B (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__41886__A (.DIODE(net478));
 sky130_as_sc_hs__diode_2 ANTENNA__41886__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__41887__A (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__41887__B (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__41891__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__41891__B (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__41899__A (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__41899__B (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__41900__A (.DIODE(net468));
 sky130_as_sc_hs__diode_2 ANTENNA__41900__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__41926__A (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__41926__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__41927__A (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__41927__B (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__41928__A (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA__41928__B (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__41950__A (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__41950__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__41951__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__41951__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__41995__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__42007__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__42008__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__42011__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__42016__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__42019__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__42022__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__42026__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__42038__A (.DIODE(\tholin_riscv.Iimm[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42042__B (.DIODE(\tholin_riscv.Iimm[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42046__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__42049__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__42054__A (.DIODE(\tholin_riscv.Iimm[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42054__B (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__42058__A (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__42058__B (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__42059__A (.DIODE(net466));
 sky130_as_sc_hs__diode_2 ANTENNA__42059__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__42060__A (.DIODE(net474));
 sky130_as_sc_hs__diode_2 ANTENNA__42060__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__42061__A (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__42061__B (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__42065__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__42065__B (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__42094__A (.DIODE(net121));
 sky130_as_sc_hs__diode_2 ANTENNA__42094__B (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__42095__A (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__42095__B (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__42096__A (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__42096__B (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__42115__A (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA__42115__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__42116__A (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__42116__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__42169__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__42171__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__42174__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__42176__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__42182__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__42186__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__42199__B (.DIODE(\tholin_riscv.Iimm[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42203__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__42211__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__42216__A (.DIODE(\tholin_riscv.Iimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42216__B (.DIODE(\tholin_riscv.io_size[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42219__A (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__42219__B (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__42220__A (.DIODE(net83));
 sky130_as_sc_hs__diode_2 ANTENNA__42220__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__42221__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__42221__B (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__42225__A (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__42225__B (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__42248__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__42248__B (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__42249__A (.DIODE(net436));
 sky130_as_sc_hs__diode_2 ANTENNA__42249__B (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA__42250__A (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__42250__B (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__42268__A (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA__42268__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__42269__A (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__42269__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__42312__A (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__42322__A (.DIODE(_05606_));
 sky130_as_sc_hs__diode_2 ANTENNA__42322__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__42326__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__42332__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__42335__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__42337__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__42352__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__42358__B (.DIODE(\tholin_riscv.Iimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42362__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__42363__A (.DIODE(\tholin_riscv.Iimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42370__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__42375__B (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__42379__A (.DIODE(net121));
 sky130_as_sc_hs__diode_2 ANTENNA__42379__B (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__42380__A (.DIODE(net431));
 sky130_as_sc_hs__diode_2 ANTENNA__42380__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__42381__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__42381__B (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__42385__A (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__42385__B (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__42404__A (.DIODE(net440));
 sky130_as_sc_hs__diode_2 ANTENNA__42404__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__42405__A (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__42405__B (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__42420__A (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__42420__B (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA__42421__A (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__42421__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__42461__A (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__42467__A (.DIODE(_05456_));
 sky130_as_sc_hs__diode_2 ANTENNA__42477__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__42478__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__42482__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__42485__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__42491__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__42496__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__42499__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__42511__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__42518__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__42520__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__42525__B (.DIODE(\tholin_riscv.io_size[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42534__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__42534__B (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__42535__A (.DIODE(net429));
 sky130_as_sc_hs__diode_2 ANTENNA__42535__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__42536__A (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__42536__B (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__42540__A (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA__42540__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__42562__A (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__42574__A (.DIODE(net121));
 sky130_as_sc_hs__diode_2 ANTENNA__42574__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__42575__A (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA__42610__A (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__42614__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__42626__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__42628__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__42631__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__42633__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__42637__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__42642__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__42645__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__42659__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__42667__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__42672__A (.DIODE(\tholin_riscv.Bimm[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42672__B (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__42676__A (.DIODE(net434));
 sky130_as_sc_hs__diode_2 ANTENNA__42676__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__42677__A (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__42677__B (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__42678__A (.DIODE(net427));
 sky130_as_sc_hs__diode_2 ANTENNA__42678__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__42679__A (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__42679__B (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__42708__A (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA__42708__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__42709__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__42709__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__42757__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__42759__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__42762__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__42764__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__42768__A (.DIODE(_05968_));
 sky130_as_sc_hs__diode_2 ANTENNA__42773__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__42776__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__42785__B (.DIODE(\tholin_riscv.Bimm[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42791__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__42798__A (.DIODE(_21569_));
 sky130_as_sc_hs__diode_2 ANTENNA__42800__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__42805__A (.DIODE(\tholin_riscv.Bimm[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42805__B (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__42808__A (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__42808__B (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__42810__A (.DIODE(net120));
 sky130_as_sc_hs__diode_2 ANTENNA__42810__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__42811__A (.DIODE(net433));
 sky130_as_sc_hs__diode_2 ANTENNA__42811__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__42834__A (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA__42834__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__42835__A (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__42835__B (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__42868__A (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__42873__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__42887__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__42889__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__42892__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__42894__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__42898__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__42903__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__42906__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__42916__B (.DIODE(\tholin_riscv.Bimm[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42920__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__42921__A (.DIODE(\tholin_riscv.Bimm[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42928__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__42933__B (.DIODE(\tholin_riscv.io_size[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__42937__A (.DIODE(net425));
 sky130_as_sc_hs__diode_2 ANTENNA__42937__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__42941__A (.DIODE(net122));
 sky130_as_sc_hs__diode_2 ANTENNA__42961__A (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__42961__B (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__42962__A (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__42962__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__42989__A (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__42994__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__43008__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__43010__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__43013__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__43015__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__43019__A (.DIODE(_05968_));
 sky130_as_sc_hs__diode_2 ANTENNA__43024__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__43027__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__43051__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__43056__B (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__43060__A (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__43060__B (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__43072__A (.DIODE(net128));
 sky130_as_sc_hs__diode_2 ANTENNA__43072__B (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA__43073__A (.DIODE(net421));
 sky130_as_sc_hs__diode_2 ANTENNA__43073__B (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA__43109__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__43113__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__43124__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__43126__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__43131__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__43134__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__43135__A (.DIODE(net140));
 sky130_as_sc_hs__diode_2 ANTENNA__43140__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__43143__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__43156__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__43164__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__43169__A (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__43170__A (.DIODE(net423));
 sky130_as_sc_hs__diode_2 ANTENNA__43171__A (.DIODE(net419));
 sky130_as_sc_hs__diode_2 ANTENNA__43219__A (.DIODE(net118));
 sky130_as_sc_hs__diode_2 ANTENNA__43221__A (.DIODE(net414));
 sky130_as_sc_hs__diode_2 ANTENNA__43224__A (.DIODE(net110));
 sky130_as_sc_hs__diode_2 ANTENNA__43226__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__43230__A (.DIODE(_05968_));
 sky130_as_sc_hs__diode_2 ANTENNA__43235__B (.DIODE(_06161_));
 sky130_as_sc_hs__diode_2 ANTENNA__43238__A (.DIODE(net412));
 sky130_as_sc_hs__diode_2 ANTENNA__43249__B (.DIODE(\tholin_riscv.Bimm[9] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43253__A (.DIODE(net117));
 sky130_as_sc_hs__diode_2 ANTENNA__43258__A (.DIODE(\tholin_riscv.Bimm[9] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43261__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__43262__A (.DIODE(\tholin_riscv.Bimm[9] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43262__B (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__43271__A (.DIODE(net418));
 sky130_as_sc_hs__diode_2 ANTENNA__43271__B (.DIODE(net74));
 sky130_as_sc_hs__diode_2 ANTENNA__43293__A (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__43297__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__43302__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__43305__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__43307__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__43311__A (.DIODE(_05968_));
 sky130_as_sc_hs__diode_2 ANTENNA__43318__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__43336__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__43342__B (.DIODE(\tholin_riscv.Bimm[10] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43351__A (.DIODE(\tholin_riscv.Bimm[10] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43354__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__43355__A (.DIODE(\tholin_riscv.Bimm[10] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43355__B (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__43362__A (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__43362__B (.DIODE(\tholin_riscv.io_size[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43375__A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA__43384__A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA__43385__B (.DIODE(_05505_));
 sky130_as_sc_hs__diode_2 ANTENNA__43389__A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA__43391__A (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__43394__A (.DIODE(net109));
 sky130_as_sc_hs__diode_2 ANTENNA__43396__A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA__43399__A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA__43400__B (.DIODE(_05968_));
 sky130_as_sc_hs__diode_2 ANTENNA__43407__A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA__43418__B (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__43425__A (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__43432__A (.DIODE(_21546_));
 sky130_as_sc_hs__diode_2 ANTENNA__43439__A (.DIODE(_21576_));
 sky130_as_sc_hs__diode_2 ANTENNA__43939__A (.DIODE(\tholin_riscv.Jimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43941__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__43968__A (.DIODE(\tholin_riscv.Bimm[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43968__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__43972__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__43973__B (.DIODE(\tholin_riscv.Bimm[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43974__A (.DIODE(\tholin_riscv.Bimm[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43976__A (.DIODE(\tholin_riscv.Bimm[9] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43977__A (.DIODE(\tholin_riscv.Iimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43977__B (.DIODE(\tholin_riscv.Iimm[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__43983__C (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__43989__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__43990__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__43999__A (.DIODE(net502));
 sky130_as_sc_hs__diode_2 ANTENNA__44593__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44594__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44595__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44596__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44597__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44598__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44599__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44600__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44601__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44602__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44603__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44604__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44605__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44606__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44607__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44608__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44609__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44610__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44611__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44612__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44613__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44614__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44615__B (.DIODE(_13479_));
 sky130_as_sc_hs__diode_2 ANTENNA__44616__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44617__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44618__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44619__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44620__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44621__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44622__B (.DIODE(net76));
 sky130_as_sc_hs__diode_2 ANTENNA__44623__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44624__B (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA__44725__B (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__44725__C (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__44734__A (.DIODE(net502));
 sky130_as_sc_hs__diode_2 ANTENNA__46263__B (.DIODE(net12));
 sky130_as_sc_hs__diode_2 ANTENNA__46293__B (.DIODE(_14629_));
 sky130_as_sc_hs__diode_2 ANTENNA__46531__A (.DIODE(net526));
 sky130_as_sc_hs__diode_2 ANTENNA__46536__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__46540__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__46552__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__46564__A (.DIODE(_00988_));
 sky130_as_sc_hs__diode_2 ANTENNA__46568__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__46575__B (.DIODE(_14629_));
 sky130_as_sc_hs__diode_2 ANTENNA__46576__A (.DIODE(\tholin_riscv.instr[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__46581__B (.DIODE(_14629_));
 sky130_as_sc_hs__diode_2 ANTENNA__46582__A (.DIODE(\tholin_riscv.instr[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__46587__B (.DIODE(_14629_));
 sky130_as_sc_hs__diode_2 ANTENNA__46593__B (.DIODE(_14629_));
 sky130_as_sc_hs__diode_2 ANTENNA__46599__B (.DIODE(_14629_));
 sky130_as_sc_hs__diode_2 ANTENNA__46605__B (.DIODE(_14629_));
 sky130_as_sc_hs__diode_2 ANTENNA__46611__B (.DIODE(_14629_));
 sky130_as_sc_hs__diode_2 ANTENNA__46617__B (.DIODE(_14629_));
 sky130_as_sc_hs__diode_2 ANTENNA__46618__A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA__46623__B (.DIODE(_14629_));
 sky130_as_sc_hs__diode_2 ANTENNA__46624__A (.DIODE(_19528_));
 sky130_as_sc_hs__diode_2 ANTENNA__46630__A (.DIODE(_00988_));
 sky130_as_sc_hs__diode_2 ANTENNA__46645__A (.DIODE(_00988_));
 sky130_as_sc_hs__diode_2 ANTENNA__46646__B (.DIODE(_14629_));
 sky130_as_sc_hs__diode_2 ANTENNA__46651__B (.DIODE(net12));
 sky130_as_sc_hs__diode_2 ANTENNA__46652__A (.DIODE(_19528_));
 sky130_as_sc_hs__diode_2 ANTENNA__46665__A (.DIODE(net526));
 sky130_as_sc_hs__diode_2 ANTENNA__46677__A (.DIODE(net526));
 sky130_as_sc_hs__diode_2 ANTENNA__46687__A (.DIODE(net12));
 sky130_as_sc_hs__diode_2 ANTENNA__46728__A (.DIODE(net522));
 sky130_as_sc_hs__diode_2 ANTENNA__46893__A (.DIODE(_19528_));
 sky130_as_sc_hs__diode_2 ANTENNA__46897__A (.DIODE(_19528_));
 sky130_as_sc_hs__diode_2 ANTENNA__46923__A (.DIODE(\tholin_riscv.instr[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__46927__A (.DIODE(\tholin_riscv.instr[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__46937__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__46943__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__46963__A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA__46979__A (.DIODE(net522));
 sky130_as_sc_hs__diode_2 ANTENNA__46983__A (.DIODE(net522));
 sky130_as_sc_hs__diode_2 ANTENNA__46987__A (.DIODE(net522));
 sky130_as_sc_hs__diode_2 ANTENNA__47005__A (.DIODE(net1168));
 sky130_as_sc_hs__diode_2 ANTENNA__47009__A (.DIODE(net1374));
 sky130_as_sc_hs__diode_2 ANTENNA__47013__A (.DIODE(net1343));
 sky130_as_sc_hs__diode_2 ANTENNA__47025__A (.DIODE(net1032));
 sky130_as_sc_hs__diode_2 ANTENNA__47069__A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA__47072__A (.DIODE(net1710));
 sky130_as_sc_hs__diode_2 ANTENNA__47075__A (.DIODE(net1168));
 sky130_as_sc_hs__diode_2 ANTENNA__47078__A (.DIODE(net1374));
 sky130_as_sc_hs__diode_2 ANTENNA__47085__A (.DIODE(net145));
 sky130_as_sc_hs__diode_2 ANTENNA__47085__B (.DIODE(net134));
 sky130_as_sc_hs__diode_2 ANTENNA__47089__C (.DIODE(net134));
 sky130_as_sc_hs__diode_2 ANTENNA__47092__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__47099__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__47106__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__47113__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__47120__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__47232__B (.DIODE(net116));
 sky130_as_sc_hs__diode_2 ANTENNA__47275__A (.DIODE(_20622_));
 sky130_as_sc_hs__diode_2 ANTENNA__47280__A (.DIODE(_20707_));
 sky130_as_sc_hs__diode_2 ANTENNA__47332__B (.DIODE(_15529_));
 sky130_as_sc_hs__diode_2 ANTENNA__47387__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__47391__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__47395__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__47399__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__47403__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__47407__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__47411__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__47415__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__47419__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__47423__A (.DIODE(net496));
 sky130_as_sc_hs__diode_2 ANTENNA__47427__A (.DIODE(net496));
 sky130_as_sc_hs__diode_2 ANTENNA__47431__A (.DIODE(net496));
 sky130_as_sc_hs__diode_2 ANTENNA__47455__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__47459__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__47463__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__47467__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__47499__A (.DIODE(net496));
 sky130_as_sc_hs__diode_2 ANTENNA__47503__A (.DIODE(net496));
 sky130_as_sc_hs__diode_2 ANTENNA__47505__A (.DIODE(net145));
 sky130_as_sc_hs__diode_2 ANTENNA__47505__B (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA__47507__A (.DIODE(net526));
 sky130_as_sc_hs__diode_2 ANTENNA__47510__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47512__A (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47513__B (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47516__B (.DIODE(_06548_));
 sky130_as_sc_hs__diode_2 ANTENNA__47519__A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA__47522__B (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47523__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__47526__A (.DIODE(_21977_));
 sky130_as_sc_hs__diode_2 ANTENNA__47526__B (.DIODE(_06548_));
 sky130_as_sc_hs__diode_2 ANTENNA__47527__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47535__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47537__A (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47538__B (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47542__B (.DIODE(_06548_));
 sky130_as_sc_hs__diode_2 ANTENNA__47543__A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA__47545__A (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47546__B (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47547__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__47551__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47558__C (.DIODE(_06548_));
 sky130_as_sc_hs__diode_2 ANTENNA__47564__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__47567__A (.DIODE(_22622_));
 sky130_as_sc_hs__diode_2 ANTENNA__47567__B (.DIODE(_06548_));
 sky130_as_sc_hs__diode_2 ANTENNA__47568__A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA__47572__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__47576__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47580__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__47584__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47586__A (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47587__B (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47591__A (.DIODE(_22430_));
 sky130_as_sc_hs__diode_2 ANTENNA__47591__B (.DIODE(_06548_));
 sky130_as_sc_hs__diode_2 ANTENNA__47592__A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA__47595__B (.DIODE(_15290_));
 sky130_as_sc_hs__diode_2 ANTENNA__47596__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__47600__A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA__47602__A (.DIODE(_15290_));
 sky130_as_sc_hs__diode_2 ANTENNA__47604__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__47608__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47610__A (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47611__B (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47615__B (.DIODE(_06548_));
 sky130_as_sc_hs__diode_2 ANTENNA__47616__A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA__47620__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__47624__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47632__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47640__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47642__A (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47643__B (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47648__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47656__A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA__47660__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__47664__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47672__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47676__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__47680__A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA__47684__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__47687__A (.DIODE(_23141_));
 sky130_as_sc_hs__diode_2 ANTENNA__47687__B (.DIODE(_06548_));
 sky130_as_sc_hs__diode_2 ANTENNA__47688__A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA__47692__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__47696__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47704__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47706__A (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47707__B (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47712__A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA__47716__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__47719__B (.DIODE(_06548_));
 sky130_as_sc_hs__diode_2 ANTENNA__47720__A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA__47724__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__47727__B (.DIODE(_06548_));
 sky130_as_sc_hs__diode_2 ANTENNA__47728__A (.DIODE(net143));
 sky130_as_sc_hs__diode_2 ANTENNA__47736__A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA__47740__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__47744__A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA__47748__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__47751__A (.DIODE(net145));
 sky130_as_sc_hs__diode_2 ANTENNA__47751__B (.DIODE(_21655_));
 sky130_as_sc_hs__diode_2 ANTENNA__47753__A (.DIODE(net102));
 sky130_as_sc_hs__diode_2 ANTENNA__47758__A (.DIODE(net116));
 sky130_as_sc_hs__diode_2 ANTENNA__47758__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47761__A (.DIODE(net134));
 sky130_as_sc_hs__diode_2 ANTENNA__47763__A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__47767__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47769__A (.DIODE(net134));
 sky130_as_sc_hs__diode_2 ANTENNA__47771__A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__47776__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47777__A (.DIODE(net134));
 sky130_as_sc_hs__diode_2 ANTENNA__47779__A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__47785__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47786__A (.DIODE(net134));
 sky130_as_sc_hs__diode_2 ANTENNA__47788__A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__47794__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47796__A (.DIODE(net134));
 sky130_as_sc_hs__diode_2 ANTENNA__47798__A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__47805__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47806__A (.DIODE(net134));
 sky130_as_sc_hs__diode_2 ANTENNA__47808__A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__47815__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47817__A (.DIODE(net134));
 sky130_as_sc_hs__diode_2 ANTENNA__47819__A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__47824__A (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47825__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47826__A (.DIODE(net134));
 sky130_as_sc_hs__diode_2 ANTENNA__47835__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47846__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47856__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47865__A (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47866__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47877__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47885__A (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47886__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47897__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47905__A (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47906__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47917__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47927__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47938__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47946__A (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47947__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47958__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47966__A (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47967__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47978__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47988__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__47999__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__48009__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__48020__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__48028__A (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__48029__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__48040__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__48050__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__48061__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__48069__B (.DIODE(_15574_));
 sky130_as_sc_hs__diode_2 ANTENNA__48072__A (.DIODE(net496));
 sky130_as_sc_hs__diode_2 ANTENNA__48272__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48273__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48274__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48275__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48276__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48277__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48278__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48279__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48280__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48281__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48282__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48283__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48284__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48285__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48286__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48287__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48288__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48289__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48290__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48291__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48292__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48293__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48294__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48295__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48296__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48298__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48299__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48300__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48301__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48302__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48303__B (.DIODE(_16371_));
 sky130_as_sc_hs__diode_2 ANTENNA__48309__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__48314__A (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__48314__B (.DIODE(_19755_));
 sky130_as_sc_hs__diode_2 ANTENNA__48315__A (.DIODE(_19750_));
 sky130_as_sc_hs__diode_2 ANTENNA__48320__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__48324__B (.DIODE(net134));
 sky130_as_sc_hs__diode_2 ANTENNA__48328__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__48330__A (.DIODE(_19755_));
 sky130_as_sc_hs__diode_2 ANTENNA__48330__B (.DIODE(_19761_));
 sky130_as_sc_hs__diode_2 ANTENNA__48331__A (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48338__A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__48341__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__48342__A (.DIODE(\tholin_riscv.Bimm[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__48344__B (.DIODE(\tholin_riscv.Iimm[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__48345__A (.DIODE(\tholin_riscv.Iimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__48345__B (.DIODE(\tholin_riscv.Iimm[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__48349__A (.DIODE(net145));
 sky130_as_sc_hs__diode_2 ANTENNA__48358__A (.DIODE(net502));
 sky130_as_sc_hs__diode_2 ANTENNA__48369__A (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48369__B (.DIODE(_16428_));
 sky130_as_sc_hs__diode_2 ANTENNA__48372__A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__48379__A (.DIODE(net371));
 sky130_as_sc_hs__diode_2 ANTENNA__48379__B (.DIODE(_16428_));
 sky130_as_sc_hs__diode_2 ANTENNA__48387__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48388__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48402__B (.DIODE(_20005_));
 sky130_as_sc_hs__diode_2 ANTENNA__48403__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__48405__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48410__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48411__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48425__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__48426__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48429__A (.DIODE(net526));
 sky130_as_sc_hs__diode_2 ANTENNA__48432__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48433__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48447__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__48448__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48451__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__48454__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48455__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48468__B (.DIODE(_20005_));
 sky130_as_sc_hs__diode_2 ANTENNA__48469__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__48470__A (.DIODE(_16512_));
 sky130_as_sc_hs__diode_2 ANTENNA__48471__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48474__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__48476__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48477__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48492__A (.DIODE(_16533_));
 sky130_as_sc_hs__diode_2 ANTENNA__48493__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48496__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__48498__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48499__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48513__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__48514__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48517__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__48520__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48521__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48534__B (.DIODE(_20005_));
 sky130_as_sc_hs__diode_2 ANTENNA__48535__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__48536__A (.DIODE(_16575_));
 sky130_as_sc_hs__diode_2 ANTENNA__48537__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48542__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48543__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48557__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__48558__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48561__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__48564__A (.DIODE(net20));
 sky130_as_sc_hs__diode_2 ANTENNA__48564__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48565__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48579__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__48580__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48583__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__48586__A (.DIODE(net21));
 sky130_as_sc_hs__diode_2 ANTENNA__48586__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48587__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48600__B (.DIODE(_20005_));
 sky130_as_sc_hs__diode_2 ANTENNA__48601__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__48603__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48606__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__48608__A (.DIODE(net4));
 sky130_as_sc_hs__diode_2 ANTENNA__48608__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48609__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48625__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48630__A (.DIODE(net5));
 sky130_as_sc_hs__diode_2 ANTENNA__48630__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48631__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48645__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__48646__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48649__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__48652__A (.DIODE(net6));
 sky130_as_sc_hs__diode_2 ANTENNA__48652__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48653__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48666__B (.DIODE(_20005_));
 sky130_as_sc_hs__diode_2 ANTENNA__48667__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__48669__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48672__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__48674__A (.DIODE(net7));
 sky130_as_sc_hs__diode_2 ANTENNA__48674__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48675__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48691__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48695__A (.DIODE(_19750_));
 sky130_as_sc_hs__diode_2 ANTENNA__48696__A (.DIODE(net8));
 sky130_as_sc_hs__diode_2 ANTENNA__48696__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48697__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48710__B (.DIODE(_20005_));
 sky130_as_sc_hs__diode_2 ANTENNA__48711__A (.DIODE(net137));
 sky130_as_sc_hs__diode_2 ANTENNA__48713__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48717__A (.DIODE(_19750_));
 sky130_as_sc_hs__diode_2 ANTENNA__48717__B (.DIODE(_23598_));
 sky130_as_sc_hs__diode_2 ANTENNA__48718__A (.DIODE(net9));
 sky130_as_sc_hs__diode_2 ANTENNA__48718__B (.DIODE(_19751_));
 sky130_as_sc_hs__diode_2 ANTENNA__48719__A (.DIODE(_19759_));
 sky130_as_sc_hs__diode_2 ANTENNA__48735__A (.DIODE(_16445_));
 sky130_as_sc_hs__diode_2 ANTENNA__48743__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48746__B (.DIODE(_16428_));
 sky130_as_sc_hs__diode_2 ANTENNA__48747__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__48750__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48753__B (.DIODE(_16428_));
 sky130_as_sc_hs__diode_2 ANTENNA__48754__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__48764__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48771__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48778__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48785__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48792__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48799__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48806__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48813__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48820__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48827__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48834__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48841__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48848__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48855__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48862__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48869__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48876__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48883__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48890__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48897__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48904__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48911__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48918__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48925__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48932__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48939__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48946__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48953__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48960__B (.DIODE(_19937_));
 sky130_as_sc_hs__diode_2 ANTENNA__48966__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__48970__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__48974__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__48978__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__48982__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__48986__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__48987__A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA__48987__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__48990__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__48991__A (.DIODE(net1260));
 sky130_as_sc_hs__diode_2 ANTENNA__48991__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__48994__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__48995__A (.DIODE(net1780));
 sky130_as_sc_hs__diode_2 ANTENNA__48995__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__48998__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__48999__A (.DIODE(net1791));
 sky130_as_sc_hs__diode_2 ANTENNA__48999__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__49002__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__49003__A (.DIODE(net1792));
 sky130_as_sc_hs__diode_2 ANTENNA__49003__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__49006__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__49010__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__49014__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__49015__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__49015__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__49018__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__49022__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__49024__A (.DIODE(net499));
 sky130_as_sc_hs__diode_2 ANTENNA__49026__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__49030__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__49034__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__49036__A (.DIODE(net499));
 sky130_as_sc_hs__diode_2 ANTENNA__49038__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__49039__A (.DIODE(\tholin_riscv.Iimm[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49039__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__49042__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__49046__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__49047__A (.DIODE(\tholin_riscv.Iimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49047__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__49050__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__49054__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__49058__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__49059__A (.DIODE(\tholin_riscv.Bimm[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49059__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__49062__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__49063__A (.DIODE(\tholin_riscv.Bimm[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49063__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__49066__B (.DIODE(net105));
 sky130_as_sc_hs__diode_2 ANTENNA__49070__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__49072__A (.DIODE(net499));
 sky130_as_sc_hs__diode_2 ANTENNA__49074__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__49075__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__49076__A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__49078__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__49079__A (.DIODE(\tholin_riscv.Bimm[10] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49079__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__49082__B (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA__49083__A (.DIODE(\tholin_riscv.Bimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49083__B (.DIODE(_19931_));
 sky130_as_sc_hs__diode_2 ANTENNA__49282__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49283__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49284__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49285__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49286__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49287__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49288__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49289__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49290__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49291__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49292__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49293__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49294__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49295__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49296__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49297__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49298__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49299__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49300__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49301__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49302__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49303__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49304__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49305__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49306__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49308__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49309__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49310__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49311__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49312__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49313__B (.DIODE(_17261_));
 sky130_as_sc_hs__diode_2 ANTENNA__49451__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49456__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49457__C (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49459__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49460__A (.DIODE(\tholin_riscv.instr[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49460__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49467__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49469__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49475__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49477__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49479__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49485__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49487__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49489__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49497__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49499__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49505__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49507__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49509__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49515__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49517__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49519__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49520__A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49520__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49526__A (.DIODE(net98));
 sky130_as_sc_hs__diode_2 ANTENNA__49527__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49529__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49530__A (.DIODE(net1260));
 sky130_as_sc_hs__diode_2 ANTENNA__49530__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49531__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__49535__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49536__A (.DIODE(net98));
 sky130_as_sc_hs__diode_2 ANTENNA__49537__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49539__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49540__A (.DIODE(\tholin_riscv.Bimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49540__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49541__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__49545__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49546__A (.DIODE(net98));
 sky130_as_sc_hs__diode_2 ANTENNA__49547__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49549__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49550__A (.DIODE(net1791));
 sky130_as_sc_hs__diode_2 ANTENNA__49550__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49551__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__49557__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49559__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49560__A (.DIODE(net1792));
 sky130_as_sc_hs__diode_2 ANTENNA__49560__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49567__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49569__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49577__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49579__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49587__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49589__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49590__A (.DIODE(net1796));
 sky130_as_sc_hs__diode_2 ANTENNA__49590__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49595__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49597__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49599__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49605__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49607__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49609__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49617__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49619__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49625__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49627__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49629__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49635__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49637__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49639__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49647__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49649__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49650__A (.DIODE(\tholin_riscv.Iimm[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49650__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49657__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49659__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49666__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49668__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49669__A (.DIODE(\tholin_riscv.Iimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49669__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49676__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49678__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49683__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49685__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49687__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49692__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49694__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49696__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49697__A (.DIODE(\tholin_riscv.Bimm[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49697__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49703__A (.DIODE(net98));
 sky130_as_sc_hs__diode_2 ANTENNA__49704__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49706__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49707__A (.DIODE(\tholin_riscv.Bimm[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49707__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49711__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49712__B (.DIODE(net98));
 sky130_as_sc_hs__diode_2 ANTENNA__49713__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49715__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49720__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49721__B (.DIODE(net98));
 sky130_as_sc_hs__diode_2 ANTENNA__49722__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49724__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49726__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__49731__A (.DIODE(net98));
 sky130_as_sc_hs__diode_2 ANTENNA__49732__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49734__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49735__A (.DIODE(\tholin_riscv.Bimm[9] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49735__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49739__B (.DIODE(net81));
 sky130_as_sc_hs__diode_2 ANTENNA__49740__B (.DIODE(net98));
 sky130_as_sc_hs__diode_2 ANTENNA__49741__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49743__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49744__A (.DIODE(\tholin_riscv.Bimm[10] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49744__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49750__A (.DIODE(net98));
 sky130_as_sc_hs__diode_2 ANTENNA__49751__A (.DIODE(_16370_));
 sky130_as_sc_hs__diode_2 ANTENNA__49753__A (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49754__A (.DIODE(\tholin_riscv.Bimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49754__B (.DIODE(_17264_));
 sky130_as_sc_hs__diode_2 ANTENNA__49780__A (.DIODE(net509));
 sky130_as_sc_hs__diode_2 ANTENNA__49783__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__49786__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__49789__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__49816__A (.DIODE(net509));
 sky130_as_sc_hs__diode_2 ANTENNA__49834__A (.DIODE(net509));
 sky130_as_sc_hs__diode_2 ANTENNA__49843__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__49849__A (.DIODE(net509));
 sky130_as_sc_hs__diode_2 ANTENNA__49948__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__49950__A (.DIODE(\tholin_riscv.instr[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49950__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__49954__A (.DIODE(net1684));
 sky130_as_sc_hs__diode_2 ANTENNA__49954__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__49955__A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA__49959__A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA__49963__A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA__49967__A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA__49971__A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA__49975__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__49978__A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA__49978__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__49979__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__49982__A (.DIODE(net1260));
 sky130_as_sc_hs__diode_2 ANTENNA__49982__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__49986__A (.DIODE(net1168));
 sky130_as_sc_hs__diode_2 ANTENNA__49986__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__49990__A (.DIODE(net1374));
 sky130_as_sc_hs__diode_2 ANTENNA__49990__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__49994__A (.DIODE(net1343));
 sky130_as_sc_hs__diode_2 ANTENNA__49994__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__50005__A (.DIODE(net1032));
 sky130_as_sc_hs__diode_2 ANTENNA__50005__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__50006__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__50010__A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA__50014__A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA__50018__A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA__50022__A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA__50026__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__50029__A (.DIODE(\tholin_riscv.Iimm[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50029__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__50030__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__50034__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__50037__A (.DIODE(\tholin_riscv.Iimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50037__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__50038__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__50042__A (.DIODE(net512));
 sky130_as_sc_hs__diode_2 ANTENNA__50049__A (.DIODE(\tholin_riscv.Bimm[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50049__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__50053__A (.DIODE(\tholin_riscv.Bimm[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50053__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__50065__A (.DIODE(\tholin_riscv.Bimm[9] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50065__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__50069__A (.DIODE(\tholin_riscv.Bimm[10] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50069__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__50073__A (.DIODE(\tholin_riscv.Bimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50073__B (.DIODE(_19962_));
 sky130_as_sc_hs__diode_2 ANTENNA__50078__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50079__A (.DIODE(\tholin_riscv.instr[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50080__A (.DIODE(net523));
 sky130_as_sc_hs__diode_2 ANTENNA__50082__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50083__A (.DIODE(net1684));
 sky130_as_sc_hs__diode_2 ANTENNA__50086__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50088__A (.DIODE(net523));
 sky130_as_sc_hs__diode_2 ANTENNA__50090__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50092__A (.DIODE(net523));
 sky130_as_sc_hs__diode_2 ANTENNA__50094__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50098__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50107__A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50108__A (.DIODE(net522));
 sky130_as_sc_hs__diode_2 ANTENNA__50111__A (.DIODE(net1260));
 sky130_as_sc_hs__diode_2 ANTENNA__50112__A (.DIODE(net522));
 sky130_as_sc_hs__diode_2 ANTENNA__50115__A (.DIODE(net1168));
 sky130_as_sc_hs__diode_2 ANTENNA__50116__A (.DIODE(net522));
 sky130_as_sc_hs__diode_2 ANTENNA__50119__A (.DIODE(net1374));
 sky130_as_sc_hs__diode_2 ANTENNA__50123__A (.DIODE(net1343));
 sky130_as_sc_hs__diode_2 ANTENNA__50126__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50130__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50132__A (.DIODE(net523));
 sky130_as_sc_hs__diode_2 ANTENNA__50134__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50135__A (.DIODE(net1032));
 sky130_as_sc_hs__diode_2 ANTENNA__50140__A (.DIODE(net523));
 sky130_as_sc_hs__diode_2 ANTENNA__50141__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50143__A (.DIODE(net523));
 sky130_as_sc_hs__diode_2 ANTENNA__50145__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50147__A (.DIODE(net523));
 sky130_as_sc_hs__diode_2 ANTENNA__50149__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50151__A (.DIODE(net523));
 sky130_as_sc_hs__diode_2 ANTENNA__50153__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50157__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50158__A (.DIODE(\tholin_riscv.Iimm[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50161__B (.DIODE(net95));
 sky130_as_sc_hs__diode_2 ANTENNA__50166__A (.DIODE(\tholin_riscv.Iimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50178__A (.DIODE(\tholin_riscv.Bimm[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50198__A (.DIODE(\tholin_riscv.Bimm[10] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50199__A (.DIODE(net522));
 sky130_as_sc_hs__diode_2 ANTENNA__50202__A (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__50341__B (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50342__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50347__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50348__C (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50350__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50351__A (.DIODE(\tholin_riscv.instr[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50351__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50358__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50360__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50366__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50368__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50370__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50376__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50378__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50380__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50388__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50390__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50396__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50398__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50400__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50406__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50408__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50410__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50411__A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50411__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50417__A (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50418__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50420__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50421__A (.DIODE(net1260));
 sky130_as_sc_hs__diode_2 ANTENNA__50421__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50427__A (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50428__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50430__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50431__A (.DIODE(net1780));
 sky130_as_sc_hs__diode_2 ANTENNA__50431__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50437__A (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50438__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50440__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50441__A (.DIODE(net1791));
 sky130_as_sc_hs__diode_2 ANTENNA__50441__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50448__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50450__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50451__A (.DIODE(net1792));
 sky130_as_sc_hs__diode_2 ANTENNA__50451__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50458__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50460__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50466__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50468__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50470__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50478__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50480__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50481__A (.DIODE(net1796));
 sky130_as_sc_hs__diode_2 ANTENNA__50481__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50486__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50487__A (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50488__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50490__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50496__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50498__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50500__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50507__A (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50508__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50510__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50516__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50518__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50520__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50526__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50528__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50530__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50532__A (.DIODE(net509));
 sky130_as_sc_hs__diode_2 ANTENNA__50537__A (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50538__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50540__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50541__A (.DIODE(\tholin_riscv.Iimm[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50541__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50547__A (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50548__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50550__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50555__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50557__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50559__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50560__A (.DIODE(\tholin_riscv.Iimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50560__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50567__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50569__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50574__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50575__B (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50576__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50578__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50583__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50585__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50587__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50588__A (.DIODE(\tholin_riscv.Bimm[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50588__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50594__A (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50595__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50597__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50598__A (.DIODE(\tholin_riscv.Bimm[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50598__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50599__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__50602__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50603__B (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50604__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50606__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50608__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__50611__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50612__B (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50613__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50615__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50622__A (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50623__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50625__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50626__A (.DIODE(\tholin_riscv.Bimm[9] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50626__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50627__A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__50630__B (.DIODE(net80));
 sky130_as_sc_hs__diode_2 ANTENNA__50631__B (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50632__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50634__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50635__A (.DIODE(\tholin_riscv.Bimm[10] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50635__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50641__A (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA__50642__A (.DIODE(_17260_));
 sky130_as_sc_hs__diode_2 ANTENNA__50644__A (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50645__A (.DIODE(\tholin_riscv.Bimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50645__B (.DIODE(_17995_));
 sky130_as_sc_hs__diode_2 ANTENNA__50650__A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA__50650__B (.DIODE(_16398_));
 sky130_as_sc_hs__diode_2 ANTENNA__50843__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__50843__B (.DIODE(net14));
 sky130_as_sc_hs__diode_2 ANTENNA__50848__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__50853__A (.DIODE(net526));
 sky130_as_sc_hs__diode_2 ANTENNA__50855__B (.DIODE(net14));
 sky130_as_sc_hs__diode_2 ANTENNA__50857__B (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA__50859__B (.DIODE(net98));
 sky130_as_sc_hs__diode_2 ANTENNA__50861__B (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__50863__B (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__50868__A (.DIODE(net1597));
 sky130_as_sc_hs__diode_2 ANTENNA__50869__A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__50873__A (.DIODE(net500));
 sky130_as_sc_hs__diode_2 ANTENNA__50876__A (.DIODE(\tholin_riscv.instr[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50877__A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__50881__B (.DIODE(_18595_));
 sky130_as_sc_hs__diode_2 ANTENNA__50882__A (.DIODE(\tholin_riscv.instr[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50883__A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA__50885__B (.DIODE(_18595_));
 sky130_as_sc_hs__diode_2 ANTENNA__50886__A (.DIODE(net1597));
 sky130_as_sc_hs__diode_2 ANTENNA__50887__A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA__50889__B (.DIODE(_18595_));
 sky130_as_sc_hs__diode_2 ANTENNA__50891__A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA__50893__B (.DIODE(_18595_));
 sky130_as_sc_hs__diode_2 ANTENNA__50895__A (.DIODE(net524));
 sky130_as_sc_hs__diode_2 ANTENNA__50897__B (.DIODE(_18595_));
 sky130_as_sc_hs__diode_2 ANTENNA__50899__A (.DIODE(net524));
 sky130_as_sc_hs__diode_2 ANTENNA__50901__B (.DIODE(_18595_));
 sky130_as_sc_hs__diode_2 ANTENNA__50903__A (.DIODE(net524));
 sky130_as_sc_hs__diode_2 ANTENNA__50908__A (.DIODE(\tholin_riscv.instr[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__50909__A (.DIODE(net523));
 sky130_as_sc_hs__diode_2 ANTENNA__50912__A (.DIODE(net1597));
 sky130_as_sc_hs__diode_2 ANTENNA__50913__A (.DIODE(net523));
 sky130_as_sc_hs__diode_2 ANTENNA__50917__A (.DIODE(net22));
 sky130_as_sc_hs__diode_2 ANTENNA__50921__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__50925__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__50929__A (.DIODE(net527));
 sky130_as_sc_hs__diode_2 ANTENNA__51032__A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA__51039__A (.DIODE(_19528_));
 sky130_as_sc_hs__diode_2 ANTENNA__51137__A (.DIODE(\tholin_riscv.Iimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__51138__A (.DIODE(\tholin_riscv.Bimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA__51138__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__51145__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51152__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51154__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51156__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__51160__A (.DIODE(\tholin_riscv.Bimm[3] ));
 sky130_as_sc_hs__diode_2 ANTENNA__51160__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__51169__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51176__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51178__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51179__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51180__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__51184__A (.DIODE(\tholin_riscv.Bimm[4] ));
 sky130_as_sc_hs__diode_2 ANTENNA__51184__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__51200__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51202__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51203__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51204__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__51208__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51209__B (.DIODE(\tholin_riscv.Bimm[5] ));
 sky130_as_sc_hs__diode_2 ANTENNA__51215__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51223__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51224__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51225__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__51228__B (.DIODE(\tholin_riscv.Bimm[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA__51235__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51241__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51242__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51244__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51245__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51246__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__51256__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51263__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51265__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51266__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51267__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__51277__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51284__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51286__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51287__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51288__A (.DIODE(net502));
 sky130_as_sc_hs__diode_2 ANTENNA__51292__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51294__B (.DIODE(\tholin_riscv.Bimm[9] ));
 sky130_as_sc_hs__diode_2 ANTENNA__51300__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51308__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51309__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51310__A (.DIODE(net502));
 sky130_as_sc_hs__diode_2 ANTENNA__51313__B (.DIODE(\tholin_riscv.Bimm[10] ));
 sky130_as_sc_hs__diode_2 ANTENNA__51320__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51327__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51329__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51330__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51331__A (.DIODE(net502));
 sky130_as_sc_hs__diode_2 ANTENNA__51334__A (.DIODE(\tholin_riscv.Iimm[0] ));
 sky130_as_sc_hs__diode_2 ANTENNA__51335__A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA__51335__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__51344__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51351__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51353__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51354__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51355__A (.DIODE(net502));
 sky130_as_sc_hs__diode_2 ANTENNA__51358__A (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__51358__B (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA__51373__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51376__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51378__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51379__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51391__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51395__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51398__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51400__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51401__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51405__A (.DIODE(net411));
 sky130_as_sc_hs__diode_2 ANTENNA__51419__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51422__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51424__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51425__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51426__A (.DIODE(net499));
 sky130_as_sc_hs__diode_2 ANTENNA__51437__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51441__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51444__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51446__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51447__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51465__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51468__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51470__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51471__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51472__A (.DIODE(net499));
 sky130_as_sc_hs__diode_2 ANTENNA__51483__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51487__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51490__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51492__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51493__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51494__A (.DIODE(net499));
 sky130_as_sc_hs__diode_2 ANTENNA__51506__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51510__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51513__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51515__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51516__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51517__A (.DIODE(net499));
 sky130_as_sc_hs__diode_2 ANTENNA__51529__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51536__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51538__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51539__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51540__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__51543__B (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__51550__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51554__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51556__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51557__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51559__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51560__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51561__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__51564__B (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__51576__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51579__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51581__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51582__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51583__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__51586__B (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__51593__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51597__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51599__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51600__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51602__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51603__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51604__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__51607__B (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__51616__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51622__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51623__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51625__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51626__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51627__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__51630__B (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__51637__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51641__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51643__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51644__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51646__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51647__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51648__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__51651__B (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__51666__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51667__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51669__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51670__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51671__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__51674__B (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__51681__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51685__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51687__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51688__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51690__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51691__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51692__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__51695__B (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__51704__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51710__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51711__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51713__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51714__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51715__A (.DIODE(net503));
 sky130_as_sc_hs__diode_2 ANTENNA__51718__B (.DIODE(\tholin_riscv.Bimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__51725__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51729__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51731__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51732__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51734__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51735__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51736__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__51739__B (.DIODE(\tholin_riscv.Bimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA__51752__B (.DIODE(net125));
 sky130_as_sc_hs__diode_2 ANTENNA__51754__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51755__A (.DIODE(_19942_));
 sky130_as_sc_hs__diode_2 ANTENNA__51757__A (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51758__B (.DIODE(_19944_));
 sky130_as_sc_hs__diode_2 ANTENNA__51759__A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA__51763__B (.DIODE(net334));
 sky130_as_sc_hs__diode_2 ANTENNA__51770__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51776__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51777__A (.DIODE(net145));
 sky130_as_sc_hs__diode_2 ANTENNA__51785__A (.DIODE(_13046_));
 sky130_as_sc_hs__diode_2 ANTENNA__51792__A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA__51793__A (.DIODE(net145));
 sky130_as_sc_hs__diode_2 ANTENNA__51894__A (.DIODE(net524));
 sky130_as_sc_hs__diode_2 ANTENNA__52416__CLK (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA__52882__D (.DIODE(_00988_));
 sky130_as_sc_hs__diode_2 ANTENNA__52990__CLK (.DIODE(clknet_4_0__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA__53011__CLK (.DIODE(clknet_4_0__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA__53202__CLK (.DIODE(clknet_4_2__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA__53547__CLK (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA__53629__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53630__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53631__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53632__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53633__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53634__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53635__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53636__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53637__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53638__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53639__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53640__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53641__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53642__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53643__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA__53644__A (.DIODE(net124));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_2_0_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_2_1_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_2_2_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_2_3_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_0__f_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_10__f_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_11__f_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_12__f_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_13__f_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_14__f_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_15__f_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_1__f_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_2__f_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_3__f_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_4__f_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_5__f_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_6__f_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_7__f_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_8__f_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_4_9__f_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_100_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_101_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_102_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_103_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_104_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_105_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_106_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_107_wb_clk_i_A (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_108_wb_clk_i_A (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_109_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_110_wb_clk_i_A (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_111_wb_clk_i_A (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_112_wb_clk_i_A (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_113_wb_clk_i_A (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_114_wb_clk_i_A (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_115_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_116_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_117_wb_clk_i_A (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_118_wb_clk_i_A (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_119_wb_clk_i_A (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_120_wb_clk_i_A (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_121_wb_clk_i_A (.DIODE(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_122_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_123_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_124_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_125_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_126_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_127_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_128_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_129_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_130_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_131_wb_clk_i_A (.DIODE(clknet_4_3__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_132_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_133_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_134_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_135_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_136_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_137_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_138_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_139_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_140_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_141_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_142_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_143_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_144_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_145_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_146_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_147_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_148_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_149_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_150_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_151_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_152_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_153_wb_clk_i_A (.DIODE(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_154_wb_clk_i_A (.DIODE(clknet_4_5__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_155_wb_clk_i_A (.DIODE(clknet_4_5__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_156_wb_clk_i_A (.DIODE(clknet_4_5__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_157_wb_clk_i_A (.DIODE(clknet_4_5__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_158_wb_clk_i_A (.DIODE(clknet_4_5__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_159_wb_clk_i_A (.DIODE(clknet_4_5__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_160_wb_clk_i_A (.DIODE(clknet_4_5__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_161_wb_clk_i_A (.DIODE(clknet_4_5__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_162_wb_clk_i_A (.DIODE(clknet_4_5__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_163_wb_clk_i_A (.DIODE(clknet_4_5__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_164_wb_clk_i_A (.DIODE(clknet_4_5__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_165_wb_clk_i_A (.DIODE(clknet_4_5__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_166_wb_clk_i_A (.DIODE(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_167_wb_clk_i_A (.DIODE(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_168_wb_clk_i_A (.DIODE(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_169_wb_clk_i_A (.DIODE(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_170_wb_clk_i_A (.DIODE(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_171_wb_clk_i_A (.DIODE(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_172_wb_clk_i_A (.DIODE(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_173_wb_clk_i_A (.DIODE(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_174_wb_clk_i_A (.DIODE(clknet_4_1__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_175_wb_clk_i_A (.DIODE(clknet_4_1__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_176_wb_clk_i_A (.DIODE(clknet_4_1__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_177_wb_clk_i_A (.DIODE(clknet_4_1__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_178_wb_clk_i_A (.DIODE(clknet_4_1__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_179_wb_clk_i_A (.DIODE(clknet_4_1__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_180_wb_clk_i_A (.DIODE(clknet_4_1__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_181_wb_clk_i_A (.DIODE(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_182_wb_clk_i_A (.DIODE(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_183_wb_clk_i_A (.DIODE(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_184_wb_clk_i_A (.DIODE(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_185_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_186_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_187_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_188_wb_clk_i_A (.DIODE(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_189_wb_clk_i_A (.DIODE(clknet_4_3__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_190_wb_clk_i_A (.DIODE(clknet_4_3__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_191_wb_clk_i_A (.DIODE(clknet_4_3__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_192_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_193_wb_clk_i_A (.DIODE(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_194_wb_clk_i_A (.DIODE(clknet_4_3__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_195_wb_clk_i_A (.DIODE(clknet_4_3__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_196_wb_clk_i_A (.DIODE(clknet_4_3__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_197_wb_clk_i_A (.DIODE(clknet_4_3__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_198_wb_clk_i_A (.DIODE(clknet_4_2__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_199_wb_clk_i_A (.DIODE(clknet_4_3__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_4_2__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_200_wb_clk_i_A (.DIODE(clknet_4_2__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_202_wb_clk_i_A (.DIODE(clknet_4_2__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_203_wb_clk_i_A (.DIODE(clknet_4_2__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_204_wb_clk_i_A (.DIODE(clknet_4_2__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_205_wb_clk_i_A (.DIODE(clknet_4_0__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_206_wb_clk_i_A (.DIODE(clknet_4_0__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_207_wb_clk_i_A (.DIODE(clknet_4_0__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_208_wb_clk_i_A (.DIODE(clknet_4_1__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_209_wb_clk_i_A (.DIODE(clknet_4_1__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_210_wb_clk_i_A (.DIODE(clknet_4_1__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_211_wb_clk_i_A (.DIODE(clknet_4_1__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_212_wb_clk_i_A (.DIODE(clknet_4_1__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_213_wb_clk_i_A (.DIODE(clknet_4_0__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_214_wb_clk_i_A (.DIODE(clknet_4_0__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_215_wb_clk_i_A (.DIODE(clknet_4_0__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_216_wb_clk_i_A (.DIODE(clknet_4_0__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_218_wb_clk_i_A (.DIODE(clknet_4_0__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_27_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_28_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_29_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_4_2__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_30_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_31_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_32_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_33_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_34_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_35_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_36_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_37_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_38_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_39_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_4_2__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_40_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_41_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_42_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_43_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_44_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_45_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_46_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_47_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_48_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_49_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_4_2__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_50_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_51_wb_clk_i_A (.DIODE(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_52_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_53_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_54_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_55_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_56_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_57_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_58_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_59_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_4_3__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_60_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_61_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_62_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_63_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_64_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_65_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_66_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_67_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_68_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_69_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_70_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_71_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_72_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_73_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_74_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_75_wb_clk_i_A (.DIODE(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_77_wb_clk_i_A (.DIODE(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_78_wb_clk_i_A (.DIODE(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_79_wb_clk_i_A (.DIODE(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_80_wb_clk_i_A (.DIODE(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_81_wb_clk_i_A (.DIODE(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_82_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_83_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_84_wb_clk_i_A (.DIODE(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_85_wb_clk_i_A (.DIODE(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_86_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_87_wb_clk_i_A (.DIODE(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_88_wb_clk_i_A (.DIODE(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_89_wb_clk_i_A (.DIODE(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_90_wb_clk_i_A (.DIODE(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_91_wb_clk_i_A (.DIODE(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_92_wb_clk_i_A (.DIODE(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_93_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_94_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_96_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_97_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_98_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_99_wb_clk_i_A (.DIODE(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout100_A (.DIODE(_15290_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout101_A (.DIODE(_15290_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout102_A (.DIODE(_15290_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout105_A (.DIODE(net106));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout107_A (.DIODE(net109));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout108_A (.DIODE(net109));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout110_A (.DIODE(net111));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout112_A (.DIODE(net113));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout113_A (.DIODE(_22167_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout114_A (.DIODE(net115));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout115_A (.DIODE(net116));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout116_A (.DIODE(_20825_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout118_A (.DIODE(net119));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout120_A (.DIODE(net121));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout122_A (.DIODE(net123));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout124_A (.DIODE(net29));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout126_A (.DIODE(net127));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout127_A (.DIODE(_05518_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout128_A (.DIODE(_02387_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout129_A (.DIODE(_02387_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout131_A (.DIODE(_16428_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout132_A (.DIODE(net134));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout133_A (.DIODE(net134));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout135_A (.DIODE(net136));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout138_A (.DIODE(net139));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout140_A (.DIODE(_05926_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout141_A (.DIODE(net142));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout143_A (.DIODE(net144));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout144_A (.DIODE(net145));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout150_A (.DIODE(net151));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout151_A (.DIODE(_19538_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout152_A (.DIODE(net153));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout153_A (.DIODE(net156));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout154_A (.DIODE(net156));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout155_A (.DIODE(net156));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout157_A (.DIODE(net160));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout158_A (.DIODE(net160));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout159_A (.DIODE(net160));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout161_A (.DIODE(net165));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout162_A (.DIODE(net165));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout163_A (.DIODE(net165));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout164_A (.DIODE(net165));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout166_A (.DIODE(net167));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout167_A (.DIODE(net173));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout168_A (.DIODE(net173));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout169_A (.DIODE(net173));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout170_A (.DIODE(net172));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout171_A (.DIODE(net172));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout172_A (.DIODE(net173));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout173_A (.DIODE(_19535_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout174_A (.DIODE(net186));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout175_A (.DIODE(net186));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout176_A (.DIODE(net179));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout178_A (.DIODE(net179));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout179_A (.DIODE(net186));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout180_A (.DIODE(net186));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout181_A (.DIODE(net182));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout182_A (.DIODE(net186));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout183_A (.DIODE(net186));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout184_A (.DIODE(net186));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout185_A (.DIODE(net186));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout186_A (.DIODE(_19535_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout187_A (.DIODE(net190));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout188_A (.DIODE(net190));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout189_A (.DIODE(net190));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout190_A (.DIODE(_19534_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout191_A (.DIODE(net195));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout192_A (.DIODE(net195));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout193_A (.DIODE(net195));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout195_A (.DIODE(_19534_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout196_A (.DIODE(_19534_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout197_A (.DIODE(net198));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout198_A (.DIODE(_19534_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout199_A (.DIODE(net200));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout200_A (.DIODE(_19534_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout201_A (.DIODE(net210));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout202_A (.DIODE(net210));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout203_A (.DIODE(net210));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout206_A (.DIODE(net210));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout207_A (.DIODE(net208));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout208_A (.DIODE(net209));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout209_A (.DIODE(net210));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout211_A (.DIODE(net219));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout212_A (.DIODE(net213));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout213_A (.DIODE(net214));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout214_A (.DIODE(net219));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout215_A (.DIODE(net219));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout216_A (.DIODE(net219));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout217_A (.DIODE(net219));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout218_A (.DIODE(net219));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout219_A (.DIODE(net230));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout220_A (.DIODE(net221));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout221_A (.DIODE(net224));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout222_A (.DIODE(net223));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout223_A (.DIODE(net224));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout224_A (.DIODE(net230));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout225_A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout226_A (.DIODE(net227));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout227_A (.DIODE(net230));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout228_A (.DIODE(net229));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout229_A (.DIODE(net230));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout231_A (.DIODE(net232));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout232_A (.DIODE(_19483_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout233_A (.DIODE(_19483_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout234_A (.DIODE(_19483_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout235_A (.DIODE(net239));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout236_A (.DIODE(net239));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout237_A (.DIODE(net238));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout238_A (.DIODE(net239));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout239_A (.DIODE(_19483_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout240_A (.DIODE(net244));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout241_A (.DIODE(net244));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout242_A (.DIODE(net244));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout243_A (.DIODE(net244));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout245_A (.DIODE(net246));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout247_A (.DIODE(net248));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout248_A (.DIODE(_00004_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout249_A (.DIODE(net250));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout250_A (.DIODE(_00003_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout251_A (.DIODE(net253));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout252_A (.DIODE(net253));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout253_A (.DIODE(_00003_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout254_A (.DIODE(net255));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout255_A (.DIODE(net256));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout256_A (.DIODE(_00002_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout257_A (.DIODE(net259));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout258_A (.DIODE(net259));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout259_A (.DIODE(_00002_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout260_A (.DIODE(net262));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout261_A (.DIODE(net262));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout262_A (.DIODE(_00002_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout263_A (.DIODE(net282));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout264_A (.DIODE(net282));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout265_A (.DIODE(net282));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout266_A (.DIODE(net282));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout267_A (.DIODE(net269));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout268_A (.DIODE(net269));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout269_A (.DIODE(net282));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout270_A (.DIODE(net275));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout271_A (.DIODE(net275));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout272_A (.DIODE(net275));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout273_A (.DIODE(net274));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout274_A (.DIODE(net275));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout275_A (.DIODE(net282));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout276_A (.DIODE(net277));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout277_A (.DIODE(net281));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout278_A (.DIODE(net281));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout279_A (.DIODE(net281));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout280_A (.DIODE(net281));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout281_A (.DIODE(net282));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout283_A (.DIODE(net291));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout284_A (.DIODE(net291));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout286_A (.DIODE(net291));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout287_A (.DIODE(net291));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout288_A (.DIODE(net291));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout289_A (.DIODE(net291));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout290_A (.DIODE(net291));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout291_A (.DIODE(net292));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout292_A (.DIODE(_00000_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout293_A (.DIODE(net307));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout295_A (.DIODE(net307));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout296_A (.DIODE(net307));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout298_A (.DIODE(net307));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout299_A (.DIODE(net307));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout300_A (.DIODE(net307));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout301_A (.DIODE(net307));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout302_A (.DIODE(net307));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout303_A (.DIODE(net306));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout304_A (.DIODE(net306));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout305_A (.DIODE(net306));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout306_A (.DIODE(net307));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout307_A (.DIODE(_00000_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout311_A (.DIODE(net333));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout312_A (.DIODE(net313));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout313_A (.DIODE(net333));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout314_A (.DIODE(net320));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout315_A (.DIODE(net320));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout316_A (.DIODE(net320));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout317_A (.DIODE(net320));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout318_A (.DIODE(net319));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout319_A (.DIODE(net320));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout320_A (.DIODE(net333));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout321_A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout322_A (.DIODE(net323));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout323_A (.DIODE(net333));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout326_A (.DIODE(net333));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout329_A (.DIODE(net332));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout330_A (.DIODE(net332));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout331_A (.DIODE(net332));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout332_A (.DIODE(net333));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout333_A (.DIODE(_00000_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout334_A (.DIODE(\tholin_riscv.Bimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout335_A (.DIODE(net336));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout336_A (.DIODE(\tholin_riscv.Jimm[19] ));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout337_A (.DIODE(net341));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout338_A (.DIODE(net341));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout339_A (.DIODE(net341));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout340_A (.DIODE(net341));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout342_A (.DIODE(net343));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout343_A (.DIODE(\tholin_riscv.Jimm[17] ));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout344_A (.DIODE(\tholin_riscv.Jimm[17] ));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout345_A (.DIODE(\tholin_riscv.Jimm[17] ));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout346_A (.DIODE(\tholin_riscv.Jimm[17] ));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout347_A (.DIODE(\tholin_riscv.Jimm[17] ));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout348_A (.DIODE(net350));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout349_A (.DIODE(net350));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout350_A (.DIODE(\tholin_riscv.Jimm[17] ));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout351_A (.DIODE(net359));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout352_A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout353_A (.DIODE(net354));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout354_A (.DIODE(net359));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout355_A (.DIODE(net359));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout356_A (.DIODE(net359));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout357_A (.DIODE(net358));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout358_A (.DIODE(net359));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout359_A (.DIODE(\tholin_riscv.Jimm[16] ));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout360_A (.DIODE(net370));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout361_A (.DIODE(net370));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout362_A (.DIODE(net363));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout363_A (.DIODE(net370));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout364_A (.DIODE(net365));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout365_A (.DIODE(net370));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout366_A (.DIODE(net370));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout367_A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout368_A (.DIODE(net369));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout369_A (.DIODE(net370));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout370_A (.DIODE(\tholin_riscv.Jimm[16] ));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout371_A (.DIODE(\tholin_riscv.io_size[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout372_A (.DIODE(net373));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout373_A (.DIODE(net410));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout377_A (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout378_A (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout379_A (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout381_A (.DIODE(net382));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout382_A (.DIODE(net410));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout383_A (.DIODE(net384));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout384_A (.DIODE(net410));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout385_A (.DIODE(net410));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout386_A (.DIODE(net410));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout387_A (.DIODE(net388));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout388_A (.DIODE(net394));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout389_A (.DIODE(net394));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout390_A (.DIODE(net394));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout391_A (.DIODE(net394));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout393_A (.DIODE(net394));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout394_A (.DIODE(net410));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout395_A (.DIODE(net396));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout396_A (.DIODE(net409));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout397_A (.DIODE(net400));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout398_A (.DIODE(net400));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout399_A (.DIODE(net400));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout400_A (.DIODE(net409));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout401_A (.DIODE(net408));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout402_A (.DIODE(net408));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout404_A (.DIODE(net408));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout405_A (.DIODE(net408));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout406_A (.DIODE(net408));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout407_A (.DIODE(net408));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout408_A (.DIODE(net409));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout409_A (.DIODE(net410));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout411_A (.DIODE(net1798));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout412_A (.DIODE(net413));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout414_A (.DIODE(net415));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout416_A (.DIODE(net417));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout418_A (.DIODE(_02550_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout419_A (.DIODE(net420));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout420_A (.DIODE(_02481_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout421_A (.DIODE(net422));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout423_A (.DIODE(net424));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout424_A (.DIODE(_25874_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout425_A (.DIODE(net426));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout427_A (.DIODE(net428));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout429_A (.DIODE(net430));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout431_A (.DIODE(net432));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout433_A (.DIODE(_25035_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout436_A (.DIODE(net437));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout438_A (.DIODE(net439));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout442_A (.DIODE(net443));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout446_A (.DIODE(net447));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout448_A (.DIODE(net449));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout450_A (.DIODE(net451));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout452_A (.DIODE(_24580_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout453_A (.DIODE(_24580_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout456_A (.DIODE(net457));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout457_A (.DIODE(_24479_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout462_A (.DIODE(net463));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout464_A (.DIODE(net465));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout470_A (.DIODE(net471));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout472_A (.DIODE(net473));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout474_A (.DIODE(net475));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout478_A (.DIODE(net479));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout479_A (.DIODE(_23643_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout480_A (.DIODE(net481));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout482_A (.DIODE(_23624_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout483_A (.DIODE(_23624_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout485_A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout486_A (.DIODE(net487));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout487_A (.DIODE(net496));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout489_A (.DIODE(net496));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout492_A (.DIODE(net496));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout493_A (.DIODE(net494));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout494_A (.DIODE(net495));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout495_A (.DIODE(net496));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout496_A (.DIODE(net524));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout497_A (.DIODE(net499));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout498_A (.DIODE(net499));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout499_A (.DIODE(net524));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout500_A (.DIODE(net502));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout501_A (.DIODE(net502));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout502_A (.DIODE(net524));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout503_A (.DIODE(net504));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout504_A (.DIODE(net524));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout505_A (.DIODE(net509));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout506_A (.DIODE(net509));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout507_A (.DIODE(net509));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout508_A (.DIODE(net509));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout509_A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout511_A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout512_A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout513_A (.DIODE(net514));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout514_A (.DIODE(net524));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout517_A (.DIODE(net522));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout518_A (.DIODE(net522));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout520_A (.DIODE(net522));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout521_A (.DIODE(net522));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout522_A (.DIODE(net523));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout523_A (.DIODE(net524));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout524_A (.DIODE(net22));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout525_A (.DIODE(net526));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout526_A (.DIODE(net22));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout527_A (.DIODE(net22));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout74_A (.DIODE(net75));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout76_A (.DIODE(net77));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout77_A (.DIODE(_13479_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout78_A (.DIODE(net79));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout83_A (.DIODE(_24939_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout84_A (.DIODE(_24939_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout87_A (.DIODE(net88));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout88_A (.DIODE(_24550_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout92_A (.DIODE(net93));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout94_A (.DIODE(_17897_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout95_A (.DIODE(_17897_));
 sky130_as_sc_hs__diode_2 ANTENNA_fanout97_A (.DIODE(net98));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1056_A (.DIODE(\tholin_riscv.instr[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1137_A (.DIODE(\tholin_riscv.Jimm[12] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1143_A (.DIODE(\tholin_riscv.instr[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1144_A (.DIODE(net1597));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1147_A (.DIODE(\tholin_riscv.Bimm[11] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1149_A (.DIODE(\tholin_riscv.Jimm[13] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1162_A (.DIODE(\tholin_riscv.requested_addr[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1169_A (.DIODE(\tholin_riscv.Bimm[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1238_A (.DIODE(\tholin_riscv.Bimm[9] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1239_A (.DIODE(\tholin_riscv.Bimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1240_A (.DIODE(\tholin_riscv.Bimm[6] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1250_A (.DIODE(\tholin_riscv.Bimm[3] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1251_A (.DIODE(\tholin_riscv.Bimm[4] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1252_A (.DIODE(\tholin_riscv.Bimm[3] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1253_A (.DIODE(\tholin_riscv.Bimm[4] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1255_A (.DIODE(\tholin_riscv.Jimm[14] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1257_A (.DIODE(\tholin_riscv.Jimm[14] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold1291_A (.DIODE(\tholin_riscv.Bimm[9] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold491_A (.DIODE(net1798));
 sky130_as_sc_hs__diode_2 ANTENNA_hold627_A (.DIODE(\tholin_riscv.Bimm[2] ));
 sky130_as_sc_hs__diode_2 ANTENNA_hold719_A (.DIODE(\tholin_riscv.Bimm[1] ));
 sky130_as_sc_hs__diode_2 ANTENNA_output29_A (.DIODE(net29));
 sky130_as_sc_hs__diode_2 ANTENNA_output55_A (.DIODE(net55));
 sky130_as_sc_hs__fill_1 FILLER_0_0_1007 ();
 sky130_as_sc_hs__decap_16 FILLER_0_0_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_1025 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_1033 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_1037 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_1045 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_1061 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_1065 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_1085 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_1089 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_1093 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_11 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_110 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_1101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_0_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_0_113 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_1142 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_1146 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_1165 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_1173 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_1177 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_1183 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_1202 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_1214 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_1218 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_1226 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_1230 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_1249 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_1257 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_129 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_137 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_157 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_166 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_169 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_188 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_0_225 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_241 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_269 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_277 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_0_29 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_305 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_309 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_317 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_321 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_324 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_332 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_353 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_361 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_365 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_383 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_391 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_393 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_400 ();
 sky130_as_sc_hs__decap_16 FILLER_0_0_421 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_437 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_445 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_45 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_465 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_473 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_481 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_500 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_513 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_517 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_524 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_53 ();
 sky130_as_sc_hs__decap_16 FILLER_0_0_533 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_549 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_557 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_561 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_578 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_586 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_641 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_663 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_667 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_671 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_691 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_695 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_699 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_701 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_709 ();
 sky130_as_sc_hs__decap_16 FILLER_0_0_729 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_73 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_745 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_753 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_773 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_781 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_789 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_799 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_807 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_810 ();
 sky130_as_sc_hs__decap_16 FILLER_0_0_813 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_829 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_837 ();
 sky130_as_sc_hs__decap_16 FILLER_0_0_841 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_85 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_857 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_865 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_869 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_873 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_890 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_894 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_897 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_0_909 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_916 ();
 sky130_as_sc_hs__decap_16 FILLER_0_0_925 ();
 sky130_as_sc_hs__fill_1 FILLER_0_0_93 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_941 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_949 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_969 ();
 sky130_as_sc_hs__decap_3 FILLER_0_0_977 ();
 sky130_as_sc_hs__fill_8 FILLER_0_0_981 ();
 sky130_as_sc_hs__fill_2 FILLER_0_0_989 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1001 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1017 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1053 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_1069 ();
 sky130_as_sc_hs__fill_8 FILLER_0_100_1077 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1093 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_110 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1125 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_114 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_132 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_136 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_147 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_156 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_168 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_189 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_212 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_218 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_227 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_234 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_248 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_25 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_253 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_260 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_264 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_267 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_271 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_275 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_279 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_283 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_295 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_307 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_309 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_317 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_323 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_332 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_34 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_349 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_370 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_382 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_386 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_403 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_429 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_461 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_487 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_554 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_574 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_585 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_594 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_60 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_625 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_641 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_659 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_66 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_669 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_680 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_75 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_776 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_804 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_808 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_813 ();
 sky130_as_sc_hs__fill_8 FILLER_0_100_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_866 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_888 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_9 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_909 ();
 sky130_as_sc_hs__fill_8 FILLER_0_100_915 ();
 sky130_as_sc_hs__fill_1 FILLER_0_100_923 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_100_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_100_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_100_977 ();
 sky130_as_sc_hs__fill_2 FILLER_0_100_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_101_1003 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_1007 ();
 sky130_as_sc_hs__fill_8 FILLER_0_101_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_1040 ();
 sky130_as_sc_hs__fill_8 FILLER_0_101_1056 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_1084 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_110 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_1100 ();
 sky130_as_sc_hs__decap_4 FILLER_0_101_1116 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_101_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_101_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_1229 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_101_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_101_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_144 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_15 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_167 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_182 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_189 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_193 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_201 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_220 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_225 ();
 sky130_as_sc_hs__decap_4 FILLER_0_101_246 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_262 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_279 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_337 ();
 sky130_as_sc_hs__decap_4 FILLER_0_101_346 ();
 sky130_as_sc_hs__decap_4 FILLER_0_101_38 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_382 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_391 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_405 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_44 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_463 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_484 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_505 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_53 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_549 ();
 sky130_as_sc_hs__decap_4 FILLER_0_101_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_577 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_61 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_663 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_669 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_687 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_711 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_716 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_734 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_749 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_774 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_781 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_804 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_808 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_812 ();
 sky130_as_sc_hs__fill_8 FILLER_0_101_828 ();
 sky130_as_sc_hs__decap_4 FILLER_0_101_836 ();
 sky130_as_sc_hs__decap_4 FILLER_0_101_846 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_850 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_87 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_877 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_889 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_895 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_101_91 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_913 ();
 sky130_as_sc_hs__fill_1 FILLER_0_101_929 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_101_953 ();
 sky130_as_sc_hs__decap_4 FILLER_0_101_969 ();
 sky130_as_sc_hs__decap_3 FILLER_0_101_973 ();
 sky130_as_sc_hs__fill_8 FILLER_0_101_995 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_1013 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_102 ();
 sky130_as_sc_hs__decap_4 FILLER_0_102_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_1033 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_106 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_1060 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_1076 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_102_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_1165 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_102_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_102_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_1261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_137 ();
 sky130_as_sc_hs__decap_4 FILLER_0_102_141 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_145 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_153 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_167 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_176 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_21 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_216 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_233 ();
 sky130_as_sc_hs__decap_4 FILLER_0_102_242 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_248 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_253 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_276 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_287 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_293 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_300 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_34 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_340 ();
 sky130_as_sc_hs__decap_4 FILLER_0_102_358 ();
 sky130_as_sc_hs__decap_4 FILLER_0_102_365 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_369 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_372 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_419 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_448 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_464 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_482 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_486 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_490 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_503 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_512 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_516 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_520 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_55 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_585 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_594 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_616 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_633 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_642 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_699 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_755 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_792 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_80 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_817 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_821 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_837 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_853 ();
 sky130_as_sc_hs__fill_8 FILLER_0_102_859 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_867 ();
 sky130_as_sc_hs__decap_4 FILLER_0_102_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_873 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_879 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_895 ();
 sky130_as_sc_hs__fill_8 FILLER_0_102_911 ();
 sky130_as_sc_hs__decap_4 FILLER_0_102_919 ();
 sky130_as_sc_hs__fill_1 FILLER_0_102_923 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_102_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_102_977 ();
 sky130_as_sc_hs__fill_2 FILLER_0_102_98 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_102_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1009 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1065 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_107 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1121 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1177 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_119 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_103_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_1273 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_130 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_146 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_166 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_183 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_188 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_201 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_22 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_220 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_230 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_249 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_258 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_262 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_281 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_313 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_333 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_342 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_364 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_370 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_377 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_383 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_39 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_425 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_43 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_434 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_476 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_495 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_501 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_505 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_539 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_552 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_561 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_572 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_576 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_586 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_590 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_609 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_67 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_670 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_673 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_700 ();
 sky130_as_sc_hs__decap_3 FILLER_0_103_706 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_71 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_734 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_817 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_825 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_833 ();
 sky130_as_sc_hs__fill_1 FILLER_0_103_868 ();
 sky130_as_sc_hs__fill_8 FILLER_0_103_897 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_905 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_914 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_930 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_94 ();
 sky130_as_sc_hs__decap_4 FILLER_0_103_946 ();
 sky130_as_sc_hs__fill_2 FILLER_0_103_950 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_103_985 ();
 sky130_as_sc_hs__decap_4 FILLER_0_104_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_104_1041 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_106 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_1068 ();
 sky130_as_sc_hs__fill_8 FILLER_0_104_1084 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_104_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_1149 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_115 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_104_1197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_120 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_1237 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_124 ();
 sky130_as_sc_hs__decap_4 FILLER_0_104_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_128 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_137 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_156 ();
 sky130_as_sc_hs__fill_1 FILLER_0_104_185 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_202 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_222 ();
 sky130_as_sc_hs__fill_1 FILLER_0_104_253 ();
 sky130_as_sc_hs__decap_4 FILLER_0_104_274 ();
 sky130_as_sc_hs__fill_1 FILLER_0_104_278 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_29 ();
 sky130_as_sc_hs__fill_1 FILLER_0_104_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_306 ();
 sky130_as_sc_hs__fill_1 FILLER_0_104_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_315 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_320 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_328 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_352 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_381 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_406 ();
 sky130_as_sc_hs__fill_1 FILLER_0_104_41 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_418 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_421 ();
 sky130_as_sc_hs__decap_4 FILLER_0_104_442 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_448 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_452 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_456 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_473 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_512 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_52 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_525 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_538 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_576 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_608 ();
 sky130_as_sc_hs__fill_1 FILLER_0_104_634 ();
 sky130_as_sc_hs__fill_1 FILLER_0_104_643 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_658 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_674 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_693 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_716 ();
 sky130_as_sc_hs__decap_4 FILLER_0_104_74 ();
 sky130_as_sc_hs__fill_1 FILLER_0_104_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_80 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_809 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_817 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_825 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_829 ();
 sky130_as_sc_hs__fill_8 FILLER_0_104_845 ();
 sky130_as_sc_hs__fill_1 FILLER_0_104_85 ();
 sky130_as_sc_hs__decap_4 FILLER_0_104_853 ();
 sky130_as_sc_hs__fill_1 FILLER_0_104_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_104_866 ();
 sky130_as_sc_hs__fill_8 FILLER_0_104_893 ();
 sky130_as_sc_hs__decap_4 FILLER_0_104_901 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_104_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_104_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_104_997 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_1007 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1193 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_120 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_105_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_136 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_153 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_164 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_173 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_187 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_20 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_201 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_211 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_215 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_225 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_242 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_259 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_267 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_274 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_281 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_293 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_337 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_351 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_377 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_405 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_435 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_441 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_445 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_462 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_476 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_484 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_49 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_499 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_514 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_523 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_543 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_569 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_592 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_615 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_625 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_650 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_707 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_719 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_733 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_803 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_823 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_827 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_83 ();
 sky130_as_sc_hs__fill_8 FILLER_0_105_831 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_839 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_841 ();
 sky130_as_sc_hs__fill_8 FILLER_0_105_850 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_858 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_864 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_87 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_878 ();
 sky130_as_sc_hs__fill_8 FILLER_0_105_887 ();
 sky130_as_sc_hs__fill_1 FILLER_0_105_895 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_934 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_95 ();
 sky130_as_sc_hs__fill_2 FILLER_0_105_950 ();
 sky130_as_sc_hs__decap_16 FILLER_0_105_953 ();
 sky130_as_sc_hs__decap_4 FILLER_0_105_969 ();
 sky130_as_sc_hs__decap_3 FILLER_0_105_973 ();
 sky130_as_sc_hs__fill_8 FILLER_0_105_999 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_106_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_1033 ();
 sky130_as_sc_hs__fill_8 FILLER_0_106_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_1068 ();
 sky130_as_sc_hs__fill_8 FILLER_0_106_1084 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_106_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_106_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_1237 ();
 sky130_as_sc_hs__fill_1 FILLER_0_106_1253 ();
 sky130_as_sc_hs__fill_1 FILLER_0_106_1259 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_166 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_175 ();
 sky130_as_sc_hs__decap_4 FILLER_0_106_183 ();
 sky130_as_sc_hs__fill_1 FILLER_0_106_187 ();
 sky130_as_sc_hs__fill_1 FILLER_0_106_190 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_220 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_243 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_26 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_276 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_29 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_319 ();
 sky130_as_sc_hs__decap_4 FILLER_0_106_343 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_359 ();
 sky130_as_sc_hs__fill_1 FILLER_0_106_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_371 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_378 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_39 ();
 sky130_as_sc_hs__decap_4 FILLER_0_106_405 ();
 sky130_as_sc_hs__fill_1 FILLER_0_106_409 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_437 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_46 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_494 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_498 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_529 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_552 ();
 sky130_as_sc_hs__fill_1 FILLER_0_106_579 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_64 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_653 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_657 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_663 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_678 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_706 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_753 ();
 sky130_as_sc_hs__decap_4 FILLER_0_106_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_796 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_800 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_804 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_808 ();
 sky130_as_sc_hs__fill_1 FILLER_0_106_81 ();
 sky130_as_sc_hs__decap_4 FILLER_0_106_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_864 ();
 sky130_as_sc_hs__fill_1 FILLER_0_106_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_885 ();
 sky130_as_sc_hs__fill_8 FILLER_0_106_889 ();
 sky130_as_sc_hs__decap_4 FILLER_0_106_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_9 ();
 sky130_as_sc_hs__fill_2 FILLER_0_106_901 ();
 sky130_as_sc_hs__fill_8 FILLER_0_106_913 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_106_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_106_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_106_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_107_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_1005 ();
 sky130_as_sc_hs__fill_8 FILLER_0_107_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_107_1017 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_1021 ();
 sky130_as_sc_hs__decap_16 FILLER_0_107_1046 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_107_1065 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_108 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_1081 ();
 sky130_as_sc_hs__fill_8 FILLER_0_107_1107 ();
 sky130_as_sc_hs__decap_4 FILLER_0_107_1115 ();
 sky130_as_sc_hs__fill_1 FILLER_0_107_1119 ();
 sky130_as_sc_hs__decap_16 FILLER_0_107_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_107_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_107_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_107_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_107_1177 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_107_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_107_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_107_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_1229 ();
 sky130_as_sc_hs__fill_8 FILLER_0_107_1233 ();
 sky130_as_sc_hs__decap_4 FILLER_0_107_1241 ();
 sky130_as_sc_hs__fill_1 FILLER_0_107_1245 ();
 sky130_as_sc_hs__decap_16 FILLER_0_107_1251 ();
 sky130_as_sc_hs__fill_8 FILLER_0_107_1267 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_1275 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_128 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_137 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_142 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_146 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_150 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_164 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_17 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_191 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_204 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_222 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_229 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_244 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_248 ();
 sky130_as_sc_hs__fill_1 FILLER_0_107_26 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_263 ();
 sky130_as_sc_hs__decap_4 FILLER_0_107_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_292 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_296 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_305 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_313 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_317 ();
 sky130_as_sc_hs__decap_4 FILLER_0_107_32 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_331 ();
 sky130_as_sc_hs__decap_4 FILLER_0_107_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_343 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_347 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_376 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_38 ();
 sky130_as_sc_hs__fill_1 FILLER_0_107_383 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_409 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_430 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_454 ();
 sky130_as_sc_hs__decap_4 FILLER_0_107_469 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_47 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_483 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_500 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_52 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_524 ();
 sky130_as_sc_hs__fill_1 FILLER_0_107_561 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_594 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_598 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_626 ();
 sky130_as_sc_hs__fill_1 FILLER_0_107_641 ();
 sky130_as_sc_hs__fill_1 FILLER_0_107_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_656 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_673 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_683 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_708 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_721 ();
 sky130_as_sc_hs__fill_1 FILLER_0_107_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_771 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_781 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_785 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_79 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_807 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_825 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_833 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_841 ();
 sky130_as_sc_hs__decap_4 FILLER_0_107_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_107_897 ();
 sky130_as_sc_hs__fill_1 FILLER_0_107_903 ();
 sky130_as_sc_hs__fill_8 FILLER_0_107_908 ();
 sky130_as_sc_hs__fill_1 FILLER_0_107_92 ();
 sky130_as_sc_hs__decap_3 FILLER_0_107_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_107_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_107_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_107_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_1004 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_1020 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_1037 ();
 sky130_as_sc_hs__fill_8 FILLER_0_108_1053 ();
 sky130_as_sc_hs__decap_4 FILLER_0_108_1061 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_1065 ();
 sky130_as_sc_hs__decap_4 FILLER_0_108_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_1093 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_11 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_108_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_108_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_108_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_127 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_136 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_147 ();
 sky130_as_sc_hs__decap_4 FILLER_0_108_156 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_183 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_195 ();
 sky130_as_sc_hs__decap_4 FILLER_0_108_202 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_208 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_216 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_223 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_23 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_232 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_236 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_264 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_288 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_29 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_295 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_108_324 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_348 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_373 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_381 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_409 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_418 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_433 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_463 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_483 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_492 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_498 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_502 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_506 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_522 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_533 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_551 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_570 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_610 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_675 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_697 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_70 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_724 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_75 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_785 ();
 sky130_as_sc_hs__fill_1 FILLER_0_108_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_840 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_844 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_848 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_858 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_865 ();
 sky130_as_sc_hs__fill_2 FILLER_0_108_90 ();
 sky130_as_sc_hs__decap_3 FILLER_0_108_907 ();
 sky130_as_sc_hs__decap_4 FILLER_0_108_920 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_940 ();
 sky130_as_sc_hs__decap_16 FILLER_0_108_956 ();
 sky130_as_sc_hs__fill_8 FILLER_0_108_972 ();
 sky130_as_sc_hs__decap_4 FILLER_0_109_1003 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_1007 ();
 sky130_as_sc_hs__fill_8 FILLER_0_109_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_109_1017 ();
 sky130_as_sc_hs__decap_4 FILLER_0_109_1040 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_1044 ();
 sky130_as_sc_hs__decap_4 FILLER_0_109_106 ();
 sky130_as_sc_hs__fill_8 FILLER_0_109_1069 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_1077 ();
 sky130_as_sc_hs__decap_16 FILLER_0_109_1101 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_109_1121 ();
 sky130_as_sc_hs__decap_4 FILLER_0_109_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_109_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_109_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_109_1169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_117 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_109_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_109_1193 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_120 ();
 sky130_as_sc_hs__decap_16 FILLER_0_109_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_109_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_1229 ();
 sky130_as_sc_hs__fill_8 FILLER_0_109_1233 ();
 sky130_as_sc_hs__decap_4 FILLER_0_109_1241 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_1245 ();
 sky130_as_sc_hs__decap_16 FILLER_0_109_1252 ();
 sky130_as_sc_hs__fill_8 FILLER_0_109_1268 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_1276 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_134 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_150 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_164 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_183 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_208 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_21 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_218 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_225 ();
 sky130_as_sc_hs__decap_4 FILLER_0_109_246 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_252 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_266 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_275 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_281 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_319 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_32 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_333 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_364 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_368 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_382 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_401 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_43 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_446 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_481 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_495 ();
 sky130_as_sc_hs__decap_4 FILLER_0_109_50 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_501 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_505 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_534 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_561 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_575 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_584 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_589 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_644 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_649 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_656 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_697 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_701 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_727 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_74 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_741 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_748 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_769 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_790 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_794 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_798 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_802 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_811 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_815 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_82 ();
 sky130_as_sc_hs__decap_3 FILLER_0_109_837 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_857 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_895 ();
 sky130_as_sc_hs__decap_16 FILLER_0_109_935 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_951 ();
 sky130_as_sc_hs__decap_4 FILLER_0_109_953 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_957 ();
 sky130_as_sc_hs__fill_2 FILLER_0_109_974 ();
 sky130_as_sc_hs__fill_8 FILLER_0_109_978 ();
 sky130_as_sc_hs__decap_4 FILLER_0_109_986 ();
 sky130_as_sc_hs__fill_1 FILLER_0_109_990 ();
 sky130_as_sc_hs__fill_8 FILLER_0_109_995 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_10_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_213 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_229 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_245 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_249 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_253 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_269 ();
 sky130_as_sc_hs__fill_1 FILLER_0_10_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_285 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_301 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_305 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_309 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_325 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_341 ();
 sky130_as_sc_hs__fill_1 FILLER_0_10_357 ();
 sky130_as_sc_hs__fill_1 FILLER_0_10_363 ();
 sky130_as_sc_hs__fill_8 FILLER_0_10_370 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_378 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_391 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_416 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_426 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_430 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_10_467 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_484 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_501 ();
 sky130_as_sc_hs__fill_1 FILLER_0_10_538 ();
 sky130_as_sc_hs__fill_8 FILLER_0_10_560 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_568 ();
 sky130_as_sc_hs__fill_1 FILLER_0_10_572 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_589 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_61 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_664 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_680 ();
 sky130_as_sc_hs__fill_1 FILLER_0_10_684 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_687 ();
 sky130_as_sc_hs__fill_1 FILLER_0_10_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_741 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_753 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_757 ();
 sky130_as_sc_hs__fill_1 FILLER_0_10_761 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_764 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_77 ();
 sky130_as_sc_hs__fill_1 FILLER_0_10_778 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_809 ();
 sky130_as_sc_hs__decap_3 FILLER_0_10_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_842 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_10_882 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_888 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_892 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_896 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_912 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_922 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_958 ();
 sky130_as_sc_hs__decap_4 FILLER_0_10_974 ();
 sky130_as_sc_hs__fill_2 FILLER_0_10_978 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_10_997 ();
 sky130_as_sc_hs__fill_8 FILLER_0_110_1023 ();
 sky130_as_sc_hs__decap_4 FILLER_0_110_1031 ();
 sky130_as_sc_hs__fill_1 FILLER_0_110_1035 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_1041 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_106 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_1073 ();
 sky130_as_sc_hs__fill_8 FILLER_0_110_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_1125 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_114 ();
 sky130_as_sc_hs__decap_4 FILLER_0_110_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_1181 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_119 ();
 sky130_as_sc_hs__decap_4 FILLER_0_110_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_110_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_128 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_135 ();
 sky130_as_sc_hs__fill_1 FILLER_0_110_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_152 ();
 sky130_as_sc_hs__decap_4 FILLER_0_110_175 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_186 ();
 sky130_as_sc_hs__fill_1 FILLER_0_110_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_217 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_233 ();
 sky130_as_sc_hs__decap_4 FILLER_0_110_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_269 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_281 ();
 sky130_as_sc_hs__fill_1 FILLER_0_110_29 ();
 sky130_as_sc_hs__fill_1 FILLER_0_110_298 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_304 ();
 sky130_as_sc_hs__decap_4 FILLER_0_110_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_315 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_347 ();
 sky130_as_sc_hs__fill_1 FILLER_0_110_354 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_382 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_402 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_406 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_418 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_110_435 ();
 sky130_as_sc_hs__decap_4 FILLER_0_110_449 ();
 sky130_as_sc_hs__fill_1 FILLER_0_110_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_110_453 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_456 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_460 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_472 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_110_484 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_490 ();
 sky130_as_sc_hs__fill_1 FILLER_0_110_501 ();
 sky130_as_sc_hs__decap_4 FILLER_0_110_51 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_510 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_529 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_549 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_568 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_586 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_589 ();
 sky130_as_sc_hs__decap_4 FILLER_0_110_593 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_627 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_642 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_658 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_71 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_719 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_746 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_753 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_770 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_813 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_817 ();
 sky130_as_sc_hs__fill_1 FILLER_0_110_83 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_85 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_852 ();
 sky130_as_sc_hs__decap_4 FILLER_0_110_860 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_864 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_90 ();
 sky130_as_sc_hs__decap_3 FILLER_0_110_910 ();
 sky130_as_sc_hs__fill_1 FILLER_0_110_918 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_929 ();
 sky130_as_sc_hs__fill_2 FILLER_0_110_94 ();
 sky130_as_sc_hs__decap_16 FILLER_0_110_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_1041 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_1057 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_1063 ();
 sky130_as_sc_hs__decap_4 FILLER_0_111_1065 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_1069 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_108 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_1100 ();
 sky130_as_sc_hs__decap_4 FILLER_0_111_1116 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_111_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_111_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_1229 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_1249 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_111_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_129 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_149 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_155 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_161 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_174 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_194 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_222 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_233 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_237 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_25 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_254 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_278 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_281 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_294 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_111_330 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_337 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_34 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_367 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_387 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_393 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_40 ();
 sky130_as_sc_hs__decap_4 FILLER_0_111_405 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_409 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_420 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_424 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_428 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_432 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_444 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_457 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_46 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_462 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_474 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_485 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_513 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_518 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_534 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_54 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_551 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_577 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_581 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_585 ();
 sky130_as_sc_hs__decap_4 FILLER_0_111_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_595 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_599 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_61 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_611 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_623 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_633 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_673 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_683 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_699 ();
 sky130_as_sc_hs__decap_3 FILLER_0_111_720 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_741 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_790 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_794 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_849 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_857 ();
 sky130_as_sc_hs__decap_4 FILLER_0_111_861 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_874 ();
 sky130_as_sc_hs__fill_1 FILLER_0_111_895 ();
 sky130_as_sc_hs__fill_2 FILLER_0_111_90 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_917 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_957 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_973 ();
 sky130_as_sc_hs__decap_16 FILLER_0_111_989 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_1033 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_1037 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_1041 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_1062 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_1086 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_109 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_1090 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_1145 ();
 sky130_as_sc_hs__fill_8 FILLER_0_112_1149 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_1157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_1166 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_1182 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_1198 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_1202 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_1205 ();
 sky130_as_sc_hs__fill_8 FILLER_0_112_1221 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_1229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_1233 ();
 sky130_as_sc_hs__fill_8 FILLER_0_112_1245 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_139 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_147 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_166 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_192 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_202 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_237 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_248 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_283 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_287 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_327 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_331 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_342 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_355 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_362 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_365 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_369 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_372 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_381 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_387 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_391 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_395 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_40 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_407 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_419 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_429 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_467 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_475 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_487 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_505 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_549 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_557 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_581 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_585 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_608 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_645 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_671 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_698 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_725 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_747 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_755 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_762 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_77 ();
 sky130_as_sc_hs__fill_1 FILLER_0_112_784 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_836 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_856 ();
 sky130_as_sc_hs__fill_8 FILLER_0_112_860 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_869 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_884 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_9 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_906 ();
 sky130_as_sc_hs__fill_2 FILLER_0_112_922 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_957 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_96 ();
 sky130_as_sc_hs__decap_4 FILLER_0_112_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_112_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_112_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_1005 ();
 sky130_as_sc_hs__fill_8 FILLER_0_113_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_1017 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_1056 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_1060 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_1121 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_1177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_119 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_1249 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_1265 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_1274 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_133 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_154 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_179 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_192 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_205 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_220 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_24 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_248 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_252 ();
 sky130_as_sc_hs__fill_1 FILLER_0_113_281 ();
 sky130_as_sc_hs__fill_1 FILLER_0_113_287 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_293 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_297 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_310 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_318 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_322 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_342 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_352 ();
 sky130_as_sc_hs__fill_1 FILLER_0_113_360 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_366 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_374 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_380 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_389 ();
 sky130_as_sc_hs__fill_1 FILLER_0_113_397 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_406 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_411 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_415 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_427 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_441 ();
 sky130_as_sc_hs__fill_1 FILLER_0_113_445 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_457 ();
 sky130_as_sc_hs__fill_1 FILLER_0_113_461 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_464 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_47 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_484 ();
 sky130_as_sc_hs__fill_1 FILLER_0_113_488 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_513 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_526 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_531 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_566 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_57 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_570 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_584 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_614 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_633 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_670 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_682 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_726 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_747 ();
 sky130_as_sc_hs__fill_1 FILLER_0_113_772 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_78 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_801 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_819 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_823 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_827 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_113_862 ();
 sky130_as_sc_hs__decap_3 FILLER_0_113_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_916 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_92 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_932 ();
 sky130_as_sc_hs__decap_4 FILLER_0_113_948 ();
 sky130_as_sc_hs__decap_16 FILLER_0_113_953 ();
 sky130_as_sc_hs__fill_1 FILLER_0_113_96 ();
 sky130_as_sc_hs__fill_1 FILLER_0_113_969 ();
 sky130_as_sc_hs__fill_8 FILLER_0_113_993 ();
 sky130_as_sc_hs__fill_8 FILLER_0_114_1024 ();
 sky130_as_sc_hs__decap_4 FILLER_0_114_1032 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_1041 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_1057 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_1073 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_1109 ();
 sky130_as_sc_hs__decap_4 FILLER_0_114_1125 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_1149 ();
 sky130_as_sc_hs__decap_4 FILLER_0_114_115 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_114_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_114_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_131 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_141 ();
 sky130_as_sc_hs__decap_4 FILLER_0_114_152 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_156 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_159 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_163 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_172 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_185 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_195 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_197 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_210 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_231 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_24 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_249 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_257 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_264 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_270 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_287 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_291 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_297 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_301 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_305 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_309 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_313 ();
 sky130_as_sc_hs__decap_4 FILLER_0_114_329 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_335 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_34 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_378 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_429 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_441 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_474 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_477 ();
 sky130_as_sc_hs__decap_4 FILLER_0_114_488 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_494 ();
 sky130_as_sc_hs__decap_4 FILLER_0_114_506 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_512 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_524 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_528 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_537 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_541 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_564 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_62 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_66 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_678 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_698 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_70 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_708 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_715 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_749 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_797 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_8 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_801 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_805 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_809 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_825 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_851 ();
 sky130_as_sc_hs__fill_2 FILLER_0_114_855 ();
 sky130_as_sc_hs__fill_8 FILLER_0_114_859 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_867 ();
 sky130_as_sc_hs__fill_8 FILLER_0_114_869 ();
 sky130_as_sc_hs__decap_4 FILLER_0_114_877 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_881 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_886 ();
 sky130_as_sc_hs__decap_4 FILLER_0_114_891 ();
 sky130_as_sc_hs__fill_1 FILLER_0_114_895 ();
 sky130_as_sc_hs__fill_8 FILLER_0_114_912 ();
 sky130_as_sc_hs__decap_4 FILLER_0_114_920 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_114_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_114_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_114_981 ();
 sky130_as_sc_hs__fill_8 FILLER_0_114_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_115_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_1025 ();
 sky130_as_sc_hs__decap_4 FILLER_0_115_1041 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_1045 ();
 sky130_as_sc_hs__fill_8 FILLER_0_115_1050 ();
 sky130_as_sc_hs__decap_4 FILLER_0_115_1058 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_1065 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_1099 ();
 sky130_as_sc_hs__decap_4 FILLER_0_115_1115 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_1119 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_115_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_1173 ();
 sky130_as_sc_hs__fill_8 FILLER_0_115_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_1190 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_1206 ();
 sky130_as_sc_hs__fill_8 FILLER_0_115_1222 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_1230 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_115_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_115_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_138 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_146 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_165 ();
 sky130_as_sc_hs__decap_4 FILLER_0_115_169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_180 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_198 ();
 sky130_as_sc_hs__decap_4 FILLER_0_115_205 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_211 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_215 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_248 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_252 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_268 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_281 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_295 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_303 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_315 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_319 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_328 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_332 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_342 ();
 sky130_as_sc_hs__decap_4 FILLER_0_115_353 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_357 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_370 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_413 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_430 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_465 ();
 sky130_as_sc_hs__decap_4 FILLER_0_115_475 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_479 ();
 sky130_as_sc_hs__decap_4 FILLER_0_115_490 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_513 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_549 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_601 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_62 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_637 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_648 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_670 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_677 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_725 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_743 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_76 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_783 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_785 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_803 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_825 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_833 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_849 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_853 ();
 sky130_as_sc_hs__fill_8 FILLER_0_115_874 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_882 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_893 ();
 sky130_as_sc_hs__fill_1 FILLER_0_115_9 ();
 sky130_as_sc_hs__decap_3 FILLER_0_115_90 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_910 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_926 ();
 sky130_as_sc_hs__fill_8 FILLER_0_115_942 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_95 ();
 sky130_as_sc_hs__fill_2 FILLER_0_115_950 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_115_985 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_10 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1000 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1016 ();
 sky130_as_sc_hs__decap_4 FILLER_0_116_1032 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1056 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1072 ();
 sky130_as_sc_hs__decap_4 FILLER_0_116_1088 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_116_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1165 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_116_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1205 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1227 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1243 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_1259 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_133 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_148 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_188 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_195 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_201 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_26 ();
 sky130_as_sc_hs__decap_4 FILLER_0_116_270 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_274 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_277 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_285 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_293 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_297 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_329 ();
 sky130_as_sc_hs__decap_4 FILLER_0_116_337 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_341 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_344 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_348 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_352 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_356 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_373 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_38 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_401 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_419 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_421 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_427 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_440 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_475 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_501 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_510 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_529 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_54 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_584 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_602 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_619 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_623 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_627 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_653 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_657 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_661 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_687 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_691 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_717 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_754 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_768 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_788 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_813 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_83 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_836 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_849 ();
 sky130_as_sc_hs__fill_1 FILLER_0_116_85 ();
 sky130_as_sc_hs__fill_8 FILLER_0_116_853 ();
 sky130_as_sc_hs__decap_4 FILLER_0_116_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_865 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_869 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_91 ();
 sky130_as_sc_hs__decap_4 FILLER_0_116_918 ();
 sky130_as_sc_hs__fill_2 FILLER_0_116_922 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_116_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_116_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_116_977 ();
 sky130_as_sc_hs__decap_4 FILLER_0_117_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_117_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1065 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_108 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1085 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1101 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_117_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1177 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_117_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_117_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_117_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_128 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_140 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_144 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_16 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_185 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_192 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_211 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_223 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_232 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_236 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_240 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_247 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_251 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_255 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_266 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_274 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_281 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_314 ();
 sky130_as_sc_hs__decap_4 FILLER_0_117_320 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_363 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_37 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_372 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_376 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_380 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_410 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_414 ();
 sky130_as_sc_hs__decap_4 FILLER_0_117_426 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_430 ();
 sky130_as_sc_hs__decap_4 FILLER_0_117_44 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_446 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_458 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_463 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_48 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_486 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_499 ();
 sky130_as_sc_hs__decap_4 FILLER_0_117_505 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_509 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_520 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_558 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_574 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_594 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_605 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_614 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_625 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_630 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_634 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_638 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_650 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_654 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_670 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_673 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_682 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_687 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_691 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_710 ();
 sky130_as_sc_hs__decap_4 FILLER_0_117_72 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_727 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_729 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_773 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_785 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_789 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_800 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_83 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_833 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_849 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_858 ();
 sky130_as_sc_hs__decap_4 FILLER_0_117_862 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_866 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_876 ();
 sky130_as_sc_hs__decap_3 FILLER_0_117_893 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_911 ();
 sky130_as_sc_hs__decap_4 FILLER_0_117_92 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_927 ();
 sky130_as_sc_hs__fill_8 FILLER_0_117_943 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_951 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_953 ();
 sky130_as_sc_hs__fill_1 FILLER_0_117_96 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_117_985 ();
 sky130_as_sc_hs__fill_2 FILLER_0_117_99 ();
 sky130_as_sc_hs__decap_4 FILLER_0_118_1013 ();
 sky130_as_sc_hs__decap_3 FILLER_0_118_103 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_1037 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_1053 ();
 sky130_as_sc_hs__fill_8 FILLER_0_118_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_1106 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_111 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_1122 ();
 sky130_as_sc_hs__fill_8 FILLER_0_118_1138 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_1146 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_1165 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_118_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_118_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_1221 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_123 ();
 sky130_as_sc_hs__fill_8 FILLER_0_118_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_118_1245 ();
 sky130_as_sc_hs__decap_4 FILLER_0_118_1254 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_1258 ();
 sky130_as_sc_hs__fill_8 FILLER_0_118_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_1269 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_1275 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_134 ();
 sky130_as_sc_hs__decap_4 FILLER_0_118_151 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_157 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_161 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_175 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_202 ();
 sky130_as_sc_hs__decap_3 FILLER_0_118_229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_242 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_246 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_250 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_258 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_272 ();
 sky130_as_sc_hs__decap_3 FILLER_0_118_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_289 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_293 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_304 ();
 sky130_as_sc_hs__decap_4 FILLER_0_118_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_320 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_328 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_332 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_346 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_352 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_365 ();
 sky130_as_sc_hs__decap_3 FILLER_0_118_371 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_379 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_383 ();
 sky130_as_sc_hs__decap_3 FILLER_0_118_395 ();
 sky130_as_sc_hs__decap_4 FILLER_0_118_406 ();
 sky130_as_sc_hs__decap_3 FILLER_0_118_429 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_453 ();
 sky130_as_sc_hs__decap_3 FILLER_0_118_473 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_500 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_531 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_54 ();
 sky130_as_sc_hs__decap_4 FILLER_0_118_577 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_118_623 ();
 sky130_as_sc_hs__decap_4 FILLER_0_118_63 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_645 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_67 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_674 ();
 sky130_as_sc_hs__decap_3 FILLER_0_118_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_70 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_705 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_717 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_734 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_755 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_762 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_785 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_8 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_821 ();
 sky130_as_sc_hs__decap_3 FILLER_0_118_825 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_883 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_907 ();
 sky130_as_sc_hs__fill_2 FILLER_0_118_91 ();
 sky130_as_sc_hs__fill_1 FILLER_0_118_923 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_118_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_118_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_118_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_119_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_1005 ();
 sky130_as_sc_hs__fill_8 FILLER_0_119_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_119_101 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_1017 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_1047 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_1063 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_119_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_1137 ();
 sky130_as_sc_hs__decap_4 FILLER_0_119_1153 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_1157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_1209 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_121 ();
 sky130_as_sc_hs__decap_4 FILLER_0_119_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_1238 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_1254 ();
 sky130_as_sc_hs__decap_4 FILLER_0_119_1270 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_1274 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_134 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_174 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_180 ();
 sky130_as_sc_hs__decap_4 FILLER_0_119_196 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_200 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_208 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_216 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_225 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_244 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_291 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_297 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_310 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_37 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_370 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_379 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_390 ();
 sky130_as_sc_hs__decap_4 FILLER_0_119_393 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_407 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_432 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_447 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_484 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_498 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_513 ();
 sky130_as_sc_hs__decap_4 FILLER_0_119_538 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_561 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_580 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_636 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_65 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_660 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_670 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_678 ();
 sky130_as_sc_hs__fill_1 FILLER_0_119_727 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_753 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_79 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_828 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_893 ();
 sky130_as_sc_hs__fill_2 FILLER_0_119_902 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_909 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_925 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_93 ();
 sky130_as_sc_hs__fill_8 FILLER_0_119_941 ();
 sky130_as_sc_hs__decap_3 FILLER_0_119_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_119_985 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_11_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_225 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_241 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_277 ();
 sky130_as_sc_hs__fill_8 FILLER_0_11_281 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_289 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_300 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_304 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_312 ();
 sky130_as_sc_hs__fill_8 FILLER_0_11_316 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_324 ();
 sky130_as_sc_hs__fill_1 FILLER_0_11_328 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_331 ();
 sky130_as_sc_hs__fill_1 FILLER_0_11_335 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_35 ();
 sky130_as_sc_hs__fill_1 FILLER_0_11_353 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_356 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_375 ();
 sky130_as_sc_hs__fill_8 FILLER_0_11_379 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_403 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_418 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_445 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_449 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_453 ();
 sky130_as_sc_hs__fill_1 FILLER_0_11_457 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_489 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_500 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_512 ();
 sky130_as_sc_hs__fill_1 FILLER_0_11_537 ();
 sky130_as_sc_hs__fill_1 FILLER_0_11_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_551 ();
 sky130_as_sc_hs__decap_4 FILLER_0_11_555 ();
 sky130_as_sc_hs__fill_1 FILLER_0_11_559 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_11_598 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_613 ();
 sky130_as_sc_hs__fill_1 FILLER_0_11_617 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_623 ();
 sky130_as_sc_hs__fill_1 FILLER_0_11_634 ();
 sky130_as_sc_hs__fill_8 FILLER_0_11_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_696 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_726 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_73 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_733 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_765 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_782 ();
 sky130_as_sc_hs__decap_3 FILLER_0_11_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_814 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_834 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_854 ();
 sky130_as_sc_hs__fill_1 FILLER_0_11_858 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_89 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_927 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_934 ();
 sky130_as_sc_hs__fill_2 FILLER_0_11_948 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_11_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_120_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_120_1033 ();
 sky130_as_sc_hs__decap_3 FILLER_0_120_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_1063 ();
 sky130_as_sc_hs__fill_8 FILLER_0_120_1079 ();
 sky130_as_sc_hs__decap_4 FILLER_0_120_1087 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_1091 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_120_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_120_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_120_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_120_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_1205 ();
 sky130_as_sc_hs__fill_8 FILLER_0_120_1221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_1239 ();
 sky130_as_sc_hs__decap_4 FILLER_0_120_1255 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_1259 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_120_15 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_150 ();
 sky130_as_sc_hs__decap_4 FILLER_0_120_159 ();
 sky130_as_sc_hs__decap_4 FILLER_0_120_175 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_181 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_195 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_20 ();
 sky130_as_sc_hs__decap_4 FILLER_0_120_219 ();
 sky130_as_sc_hs__decap_3 FILLER_0_120_230 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_238 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_24 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_250 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_264 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_268 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_272 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_279 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_283 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_290 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_296 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_120_318 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_326 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_330 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_334 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_338 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_34 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_342 ();
 sky130_as_sc_hs__decap_3 FILLER_0_120_381 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_392 ();
 sky130_as_sc_hs__decap_4 FILLER_0_120_404 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_408 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_419 ();
 sky130_as_sc_hs__decap_3 FILLER_0_120_440 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_455 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_464 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_472 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_48 ();
 sky130_as_sc_hs__decap_3 FILLER_0_120_497 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_516 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_522 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_531 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_533 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_54 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_584 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_608 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_626 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_65 ();
 sky130_as_sc_hs__decap_3 FILLER_0_120_661 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_672 ();
 sky130_as_sc_hs__decap_4 FILLER_0_120_676 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_690 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_720 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_772 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_784 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_8 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_80 ();
 sky130_as_sc_hs__decap_3 FILLER_0_120_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_835 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_847 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_851 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_855 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_859 ();
 sky130_as_sc_hs__fill_1 FILLER_0_120_863 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_876 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_897 ();
 sky130_as_sc_hs__decap_4 FILLER_0_120_918 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_922 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_120_93 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_120_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_120_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_120_997 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_10 ();
 sky130_as_sc_hs__decap_4 FILLER_0_121_1004 ();
 sky130_as_sc_hs__decap_16 FILLER_0_121_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_121_1025 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_1041 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_1062 ();
 sky130_as_sc_hs__decap_4 FILLER_0_121_1065 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_121_1095 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_1099 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_121_1130 ();
 sky130_as_sc_hs__decap_16 FILLER_0_121_1146 ();
 sky130_as_sc_hs__fill_8 FILLER_0_121_1162 ();
 sky130_as_sc_hs__decap_4 FILLER_0_121_1170 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_1174 ();
 sky130_as_sc_hs__decap_16 FILLER_0_121_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_121_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_121_1209 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_122 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_1225 ();
 sky130_as_sc_hs__decap_16 FILLER_0_121_1246 ();
 sky130_as_sc_hs__fill_8 FILLER_0_121_1262 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_127 ();
 sky130_as_sc_hs__decap_4 FILLER_0_121_1270 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_1274 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_131 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_135 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_139 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_121_17 ();
 sky130_as_sc_hs__fill_1 FILLER_0_121_176 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_210 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_235 ();
 sky130_as_sc_hs__fill_1 FILLER_0_121_268 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_274 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_278 ();
 sky130_as_sc_hs__fill_1 FILLER_0_121_28 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_285 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_289 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_303 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_331 ();
 sky130_as_sc_hs__fill_1 FILLER_0_121_342 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_356 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_366 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_417 ();
 sky130_as_sc_hs__decap_4 FILLER_0_121_441 ();
 sky130_as_sc_hs__fill_1 FILLER_0_121_445 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_449 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_475 ();
 sky130_as_sc_hs__decap_4 FILLER_0_121_49 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_494 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_502 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_521 ();
 sky130_as_sc_hs__fill_1 FILLER_0_121_53 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_543 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_558 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_569 ();
 sky130_as_sc_hs__fill_1 FILLER_0_121_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_574 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_597 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_617 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_68 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_689 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_693 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_701 ();
 sky130_as_sc_hs__fill_1 FILLER_0_121_705 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_724 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_733 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_741 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_759 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_76 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_763 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_797 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_80 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_801 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_805 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_809 ();
 sky130_as_sc_hs__fill_1 FILLER_0_121_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_84 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_854 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_858 ();
 sky130_as_sc_hs__fill_1 FILLER_0_121_862 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_868 ();
 sky130_as_sc_hs__decap_3 FILLER_0_121_876 ();
 sky130_as_sc_hs__fill_2 FILLER_0_121_88 ();
 sky130_as_sc_hs__decap_16 FILLER_0_121_927 ();
 sky130_as_sc_hs__fill_8 FILLER_0_121_943 ();
 sky130_as_sc_hs__fill_1 FILLER_0_121_951 ();
 sky130_as_sc_hs__decap_16 FILLER_0_121_972 ();
 sky130_as_sc_hs__decap_16 FILLER_0_121_988 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_1013 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_1034 ();
 sky130_as_sc_hs__decap_16 FILLER_0_122_1041 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_1057 ();
 sky130_as_sc_hs__decap_16 FILLER_0_122_1063 ();
 sky130_as_sc_hs__fill_8 FILLER_0_122_1079 ();
 sky130_as_sc_hs__decap_4 FILLER_0_122_1087 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_1091 ();
 sky130_as_sc_hs__decap_16 FILLER_0_122_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_122_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_122_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_122_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_1145 ();
 sky130_as_sc_hs__fill_8 FILLER_0_122_1154 ();
 sky130_as_sc_hs__decap_4 FILLER_0_122_1162 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_1166 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_119 ();
 sky130_as_sc_hs__fill_8 FILLER_0_122_1195 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_12 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_1203 ();
 sky130_as_sc_hs__decap_16 FILLER_0_122_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_122_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_122_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_122_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_1257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_122_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_122_1271 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_1275 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_139 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_157 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_161 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_165 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_183 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_202 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_247 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_251 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_253 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_257 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_26 ();
 sky130_as_sc_hs__decap_4 FILLER_0_122_293 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_297 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_304 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_309 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_316 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_322 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_34 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_349 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_363 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_365 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_371 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_376 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_38 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_380 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_384 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_409 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_419 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_42 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_430 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_467 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_473 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_51 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_533 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_563 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_581 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_586 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_589 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_616 ();
 sky130_as_sc_hs__decap_4 FILLER_0_122_633 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_639 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_651 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_676 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_72 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_723 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_734 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_753 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_789 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_818 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_822 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_826 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_846 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_866 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_893 ();
 sky130_as_sc_hs__decap_4 FILLER_0_122_918 ();
 sky130_as_sc_hs__fill_2 FILLER_0_122_922 ();
 sky130_as_sc_hs__decap_16 FILLER_0_122_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_122_941 ();
 sky130_as_sc_hs__fill_1 FILLER_0_122_957 ();
 sky130_as_sc_hs__decap_3 FILLER_0_122_977 ();
 sky130_as_sc_hs__decap_4 FILLER_0_122_98 ();
 sky130_as_sc_hs__decap_16 FILLER_0_122_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_122_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_1003 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_1007 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_1025 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_1041 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_1045 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_1097 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_111 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_1249 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_125 ();
 sky130_as_sc_hs__fill_8 FILLER_0_123_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_138 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_14 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_164 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_184 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_190 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_202 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_213 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_22 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_231 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_249 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_255 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_276 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_291 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_304 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_308 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_334 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_337 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_344 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_349 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_353 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_357 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_361 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_38 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_384 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_398 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_431 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_444 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_454 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_460 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_469 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_488 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_503 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_510 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_517 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_52 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_541 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_553 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_557 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_561 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_584 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_588 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_591 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_595 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_599 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_617 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_656 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_668 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_683 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_746 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_750 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_773 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_78 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_798 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_825 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_829 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_833 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_841 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_123_857 ();
 sky130_as_sc_hs__fill_1 FILLER_0_123_876 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_924 ();
 sky130_as_sc_hs__fill_8 FILLER_0_123_940 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_948 ();
 sky130_as_sc_hs__fill_8 FILLER_0_123_953 ();
 sky130_as_sc_hs__decap_4 FILLER_0_123_961 ();
 sky130_as_sc_hs__decap_3 FILLER_0_123_965 ();
 sky130_as_sc_hs__decap_16 FILLER_0_123_987 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_124_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_1033 ();
 sky130_as_sc_hs__fill_8 FILLER_0_124_1037 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_1045 ();
 sky130_as_sc_hs__decap_4 FILLER_0_124_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_124_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_1149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_115 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_1165 ();
 sky130_as_sc_hs__decap_4 FILLER_0_124_1181 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_1185 ();
 sky130_as_sc_hs__fill_8 FILLER_0_124_1191 ();
 sky130_as_sc_hs__decap_4 FILLER_0_124_1199 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_1203 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_1210 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_122 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_1226 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_1242 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_1258 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_124_129 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_146 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_154 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_17 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_197 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_210 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_221 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_231 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_235 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_247 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_251 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_257 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_268 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_279 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_284 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_314 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_325 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_330 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_36 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_363 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_369 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_373 ();
 sky130_as_sc_hs__decap_4 FILLER_0_124_390 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_394 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_416 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_429 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_452 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_468 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_494 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_510 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_533 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_549 ();
 sky130_as_sc_hs__decap_4 FILLER_0_124_569 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_573 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_584 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_594 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_614 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_618 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_635 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_653 ();
 sky130_as_sc_hs__decap_4 FILLER_0_124_657 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_661 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_665 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_669 ();
 sky130_as_sc_hs__decap_4 FILLER_0_124_673 ();
 sky130_as_sc_hs__decap_4 FILLER_0_124_679 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_685 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_694 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_698 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_705 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_713 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_717 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_738 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_754 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_797 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_809 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_813 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_817 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_859 ();
 sky130_as_sc_hs__fill_2 FILLER_0_124_863 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_867 ();
 sky130_as_sc_hs__fill_1 FILLER_0_124_877 ();
 sky130_as_sc_hs__fill_8 FILLER_0_124_887 ();
 sky130_as_sc_hs__decap_4 FILLER_0_124_899 ();
 sky130_as_sc_hs__fill_8 FILLER_0_124_916 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_124_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_124_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_124_997 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_10 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_1002 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_1006 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1041 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1209 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_122 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_1249 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_1265 ();
 sky130_as_sc_hs__fill_1 FILLER_0_125_1269 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_1275 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_134 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_138 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_162 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_179 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_192 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_233 ();
 sky130_as_sc_hs__fill_1 FILLER_0_125_241 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_277 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_281 ();
 sky130_as_sc_hs__fill_1 FILLER_0_125_285 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_288 ();
 sky130_as_sc_hs__fill_1 FILLER_0_125_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_292 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_301 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_306 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_315 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_320 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_328 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_332 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_388 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_398 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_40 ();
 sky130_as_sc_hs__fill_1 FILLER_0_125_402 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_405 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_430 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_454 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_461 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_476 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_490 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_496 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_500 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_510 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_53 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_534 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_561 ();
 sky130_as_sc_hs__fill_1 FILLER_0_125_572 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_617 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_647 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_669 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_713 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_717 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_721 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_729 ();
 sky130_as_sc_hs__fill_1 FILLER_0_125_783 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_828 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_836 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_864 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_868 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_876 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_880 ();
 sky130_as_sc_hs__fill_8 FILLER_0_125_884 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_892 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_929 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_93 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_125_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_125_953 ();
 sky130_as_sc_hs__decap_4 FILLER_0_125_969 ();
 sky130_as_sc_hs__fill_1 FILLER_0_125_973 ();
 sky130_as_sc_hs__fill_2 FILLER_0_125_990 ();
 sky130_as_sc_hs__fill_8 FILLER_0_125_994 ();
 sky130_as_sc_hs__decap_4 FILLER_0_126_1013 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_1037 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_1042 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_1066 ();
 sky130_as_sc_hs__fill_8 FILLER_0_126_1082 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_1090 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_1109 ();
 sky130_as_sc_hs__decap_4 FILLER_0_126_112 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_126_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_126_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_126_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_138 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_146 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_150 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_159 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_173 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_181 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_188 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_197 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_20 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_208 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_212 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_249 ();
 sky130_as_sc_hs__decap_4 FILLER_0_126_253 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_257 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_26 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_260 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_264 ();
 sky130_as_sc_hs__decap_4 FILLER_0_126_273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_280 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_284 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_307 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_317 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_322 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_350 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_360 ();
 sky130_as_sc_hs__decap_4 FILLER_0_126_365 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_369 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_372 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_389 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_417 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_429 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_438 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_44 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_468 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_472 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_489 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_521 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_554 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_56 ();
 sky130_as_sc_hs__decap_4 FILLER_0_126_565 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_571 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_584 ();
 sky130_as_sc_hs__decap_4 FILLER_0_126_629 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_635 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_65 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_653 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_658 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_686 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_709 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_740 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_765 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_78 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_790 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_794 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_798 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_817 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_825 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_859 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_863 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_867 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_873 ();
 sky130_as_sc_hs__fill_2 FILLER_0_126_877 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_881 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_897 ();
 sky130_as_sc_hs__fill_8 FILLER_0_126_913 ();
 sky130_as_sc_hs__decap_3 FILLER_0_126_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_126_941 ();
 sky130_as_sc_hs__decap_4 FILLER_0_126_957 ();
 sky130_as_sc_hs__fill_8 FILLER_0_126_981 ();
 sky130_as_sc_hs__fill_1 FILLER_0_126_989 ();
 sky130_as_sc_hs__decap_4 FILLER_0_127_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_1009 ();
 sky130_as_sc_hs__fill_8 FILLER_0_127_1025 ();
 sky130_as_sc_hs__decap_4 FILLER_0_127_1033 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_1037 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_1084 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_1100 ();
 sky130_as_sc_hs__decap_4 FILLER_0_127_1116 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_127_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_1209 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_122 ();
 sky130_as_sc_hs__decap_4 FILLER_0_127_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_127_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_127_1273 ();
 sky130_as_sc_hs__decap_4 FILLER_0_127_130 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_134 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_142 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_17 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_183 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_192 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_200 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_214 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_220 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_233 ();
 sky130_as_sc_hs__decap_4 FILLER_0_127_240 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_244 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_252 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_276 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_306 ();
 sky130_as_sc_hs__decap_4 FILLER_0_127_330 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_337 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_34 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_371 ();
 sky130_as_sc_hs__decap_4 FILLER_0_127_381 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_385 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_388 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_447 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_449 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_476 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_492 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_496 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_500 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_505 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_52 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_526 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_561 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_579 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_583 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_638 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_642 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_648 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_652 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_671 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_683 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_71 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_756 ();
 sky130_as_sc_hs__decap_3 FILLER_0_127_760 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_79 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_796 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_800 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_809 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_819 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_823 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_833 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_855 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_859 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_863 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_867 ();
 sky130_as_sc_hs__fill_8 FILLER_0_127_887 ();
 sky130_as_sc_hs__fill_1 FILLER_0_127_895 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_897 ();
 sky130_as_sc_hs__fill_8 FILLER_0_127_913 ();
 sky130_as_sc_hs__decap_4 FILLER_0_127_921 ();
 sky130_as_sc_hs__fill_2 FILLER_0_127_93 ();
 sky130_as_sc_hs__fill_8 FILLER_0_127_944 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_127_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_128_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_128_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_1037 ();
 sky130_as_sc_hs__decap_3 FILLER_0_128_104 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_128_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_128_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_1093 ();
 sky130_as_sc_hs__decap_4 FILLER_0_128_1109 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_1113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_1120 ();
 sky130_as_sc_hs__fill_8 FILLER_0_128_1136 ();
 sky130_as_sc_hs__decap_4 FILLER_0_128_1144 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_1165 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_128_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_128_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_128_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_128_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_129 ();
 sky130_as_sc_hs__decap_3 FILLER_0_128_135 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_128_147 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_170 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_174 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_178 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_194 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_197 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_218 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_244 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_251 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_26 ();
 sky130_as_sc_hs__decap_3 FILLER_0_128_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_128_301 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_305 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_317 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_343 ();
 sky130_as_sc_hs__decap_3 FILLER_0_128_361 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_378 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_39 ();
 sky130_as_sc_hs__decap_3 FILLER_0_128_392 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_397 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_419 ();
 sky130_as_sc_hs__decap_4 FILLER_0_128_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_425 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_43 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_455 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_472 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_498 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_504 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_549 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_574 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_128_593 ();
 sky130_as_sc_hs__decap_4 FILLER_0_128_598 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_602 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_62 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_640 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_680 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_724 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_728 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_751 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_755 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_78 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_781 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_806 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_813 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_856 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_860 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_864 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_128_873 ();
 sky130_as_sc_hs__fill_8 FILLER_0_128_877 ();
 sky130_as_sc_hs__fill_1 FILLER_0_128_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_128_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_128_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_128_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_129_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_129_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_1025 ();
 sky130_as_sc_hs__decap_4 FILLER_0_129_1041 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_105 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_1065 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_108 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_1097 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_1113 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_1119 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_1149 ();
 sky130_as_sc_hs__fill_8 FILLER_0_129_1165 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_129_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_1229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_129_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_129_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_140 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_154 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_158 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_16 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_165 ();
 sky130_as_sc_hs__decap_4 FILLER_0_129_174 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_178 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_20 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_211 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_235 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_249 ();
 sky130_as_sc_hs__decap_4 FILLER_0_129_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_264 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_268 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_29 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_294 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_323 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_328 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_332 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_341 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_361 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_38 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_409 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_415 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_426 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_438 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_457 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_474 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_483 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_50 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_517 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_537 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_580 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_641 ();
 sky130_as_sc_hs__decap_4 FILLER_0_129_645 ();
 sky130_as_sc_hs__decap_4 FILLER_0_129_651 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_655 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_658 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_666 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_670 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_697 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_727 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_754 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_758 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_76 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_762 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_766 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_783 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_83 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_835 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_861 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_865 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_869 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_873 ();
 sky130_as_sc_hs__fill_1 FILLER_0_129_895 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_913 ();
 sky130_as_sc_hs__fill_2 FILLER_0_129_92 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_129_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_129_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_129_985 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1037 ();
 sky130_as_sc_hs__fill_1 FILLER_0_12_105 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1069 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_108 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1109 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_112 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1165 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1205 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_122 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_1257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_126 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_12_130 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_133 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_138 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_12_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_213 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_229 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_245 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_249 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_253 ();
 sky130_as_sc_hs__fill_8 FILLER_0_12_269 ();
 sky130_as_sc_hs__fill_1 FILLER_0_12_27 ();
 sky130_as_sc_hs__fill_1 FILLER_0_12_277 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_12_307 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_322 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_333 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_337 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_341 ();
 sky130_as_sc_hs__fill_1 FILLER_0_12_345 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_350 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_389 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_416 ();
 sky130_as_sc_hs__fill_1 FILLER_0_12_440 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_45 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_465 ();
 sky130_as_sc_hs__fill_1 FILLER_0_12_469 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_494 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_529 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_547 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_554 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_561 ();
 sky130_as_sc_hs__fill_1 FILLER_0_12_565 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_574 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_586 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_598 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_602 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_632 ();
 sky130_as_sc_hs__fill_1 FILLER_0_12_656 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_665 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_669 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_694 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_701 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_739 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_743 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_77 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_846 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_858 ();
 sky130_as_sc_hs__fill_1 FILLER_0_12_862 ();
 sky130_as_sc_hs__fill_1 FILLER_0_12_894 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_914 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_918 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_922 ();
 sky130_as_sc_hs__fill_2 FILLER_0_12_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_12_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_12_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_12_997 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_1013 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_102 ();
 sky130_as_sc_hs__decap_4 FILLER_0_130_1029 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_1033 ();
 sky130_as_sc_hs__fill_8 FILLER_0_130_1053 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_1061 ();
 sky130_as_sc_hs__decap_4 FILLER_0_130_1067 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_1071 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_1097 ();
 sky130_as_sc_hs__fill_8 FILLER_0_130_1113 ();
 sky130_as_sc_hs__decap_4 FILLER_0_130_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_1125 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_1147 ();
 sky130_as_sc_hs__decap_3 FILLER_0_130_1164 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_1187 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_1203 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_1237 ();
 sky130_as_sc_hs__decap_3 FILLER_0_130_124 ();
 sky130_as_sc_hs__decap_4 FILLER_0_130_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_130_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_132 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_136 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_145 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_152 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_158 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_172 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_181 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_130_193 ();
 sky130_as_sc_hs__decap_3 FILLER_0_130_197 ();
 sky130_as_sc_hs__decap_4 FILLER_0_130_215 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_219 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_227 ();
 sky130_as_sc_hs__decap_3 FILLER_0_130_25 ();
 sky130_as_sc_hs__decap_4 FILLER_0_130_253 ();
 sky130_as_sc_hs__decap_4 FILLER_0_130_264 ();
 sky130_as_sc_hs__decap_4 FILLER_0_130_278 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_29 ();
 sky130_as_sc_hs__decap_4 FILLER_0_130_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_314 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_352 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_416 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_421 ();
 sky130_as_sc_hs__decap_3 FILLER_0_130_440 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_445 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_465 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_475 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_490 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_50 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_523 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_533 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_548 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_565 ();
 sky130_as_sc_hs__decap_4 FILLER_0_130_569 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_573 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_576 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_584 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_589 ();
 sky130_as_sc_hs__decap_4 FILLER_0_130_609 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_619 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_623 ();
 sky130_as_sc_hs__decap_3 FILLER_0_130_627 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_632 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_636 ();
 sky130_as_sc_hs__decap_3 FILLER_0_130_64 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_640 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_664 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_668 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_672 ();
 sky130_as_sc_hs__decap_3 FILLER_0_130_676 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_681 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_688 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_692 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_696 ();
 sky130_as_sc_hs__decap_3 FILLER_0_130_717 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_755 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_792 ();
 sky130_as_sc_hs__fill_1 FILLER_0_130_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_864 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_130_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_130_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_941 ();
 sky130_as_sc_hs__fill_2 FILLER_0_130_95 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_130_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_130_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_130_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_131_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_1009 ();
 sky130_as_sc_hs__fill_8 FILLER_0_131_1025 ();
 sky130_as_sc_hs__fill_1 FILLER_0_131_1033 ();
 sky130_as_sc_hs__decap_4 FILLER_0_131_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_131_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_1121 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_131_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_1173 ();
 sky130_as_sc_hs__fill_1 FILLER_0_131_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_131_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_1229 ();
 sky130_as_sc_hs__fill_8 FILLER_0_131_1233 ();
 sky130_as_sc_hs__decap_4 FILLER_0_131_1241 ();
 sky130_as_sc_hs__fill_1 FILLER_0_131_1245 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_1254 ();
 sky130_as_sc_hs__decap_4 FILLER_0_131_1270 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_1274 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_13 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_131_177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_183 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_200 ();
 sky130_as_sc_hs__decap_4 FILLER_0_131_216 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_220 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_225 ();
 sky130_as_sc_hs__fill_1 FILLER_0_131_237 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_25 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_270 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_281 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_302 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_313 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_328 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_332 ();
 sky130_as_sc_hs__decap_4 FILLER_0_131_337 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_34 ();
 sky130_as_sc_hs__fill_1 FILLER_0_131_341 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_344 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_374 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_416 ();
 sky130_as_sc_hs__decap_4 FILLER_0_131_42 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_472 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_48 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_482 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_52 ();
 sky130_as_sc_hs__fill_1 FILLER_0_131_559 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_561 ();
 sky130_as_sc_hs__fill_1 FILLER_0_131_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_587 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_614 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_625 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_63 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_646 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_653 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_67 ();
 sky130_as_sc_hs__fill_1 FILLER_0_131_671 ();
 sky130_as_sc_hs__fill_1 FILLER_0_131_708 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_71 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_80 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_813 ();
 sky130_as_sc_hs__decap_4 FILLER_0_131_84 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_860 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_864 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_880 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_131_90 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_131_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_131_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_131_985 ();
 sky130_as_sc_hs__fill_8 FILLER_0_132_1002 ();
 sky130_as_sc_hs__decap_4 FILLER_0_132_1010 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_1014 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_1034 ();
 sky130_as_sc_hs__fill_8 FILLER_0_132_1041 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_1049 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_106 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_1070 ();
 sky130_as_sc_hs__decap_16 FILLER_0_132_1097 ();
 sky130_as_sc_hs__decap_16 FILLER_0_132_1113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_132_1129 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_132_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_132_1165 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_132_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_132_1197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_12 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_132_1205 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_132_1221 ();
 sky130_as_sc_hs__fill_8 FILLER_0_132_1237 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_1245 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_125 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_1259 ();
 sky130_as_sc_hs__decap_16 FILLER_0_132_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_129 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_133 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_151 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_155 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_16 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_132_184 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_188 ();
 sky130_as_sc_hs__decap_4 FILLER_0_132_202 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_206 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_224 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_235 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_240 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_248 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_25 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_279 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_283 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_287 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_291 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_309 ();
 sky130_as_sc_hs__decap_4 FILLER_0_132_320 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_324 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_346 ();
 sky130_as_sc_hs__decap_4 FILLER_0_132_36 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_365 ();
 sky130_as_sc_hs__decap_4 FILLER_0_132_393 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_397 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_400 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_434 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_462 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_492 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_496 ();
 sky130_as_sc_hs__decap_4 FILLER_0_132_505 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_509 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_512 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_516 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_520 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_524 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_528 ();
 sky130_as_sc_hs__decap_4 FILLER_0_132_533 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_537 ();
 sky130_as_sc_hs__decap_4 FILLER_0_132_561 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_565 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_587 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_594 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_631 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_638 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_667 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_67 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_694 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_698 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_701 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_723 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_753 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_762 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_766 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_770 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_78 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_784 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_788 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_792 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_796 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_8 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_800 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_809 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_818 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_822 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_826 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_83 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_830 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_834 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_842 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_846 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_850 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_854 ();
 sky130_as_sc_hs__fill_8 FILLER_0_132_858 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_866 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_869 ();
 sky130_as_sc_hs__fill_8 FILLER_0_132_889 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_897 ();
 sky130_as_sc_hs__fill_1 FILLER_0_132_90 ();
 sky130_as_sc_hs__decap_4 FILLER_0_132_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_132_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_132_944 ();
 sky130_as_sc_hs__decap_16 FILLER_0_132_960 ();
 sky130_as_sc_hs__decap_4 FILLER_0_132_976 ();
 sky130_as_sc_hs__fill_2 FILLER_0_132_981 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_1025 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_1045 ();
 sky130_as_sc_hs__fill_8 FILLER_0_133_1049 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_1065 ();
 sky130_as_sc_hs__fill_8 FILLER_0_133_1081 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_1089 ();
 sky130_as_sc_hs__fill_1 FILLER_0_133_1093 ();
 sky130_as_sc_hs__fill_8 FILLER_0_133_1112 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_1254 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_1270 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_1274 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_135 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_148 ();
 sky130_as_sc_hs__fill_1 FILLER_0_133_152 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_133_200 ();
 sky130_as_sc_hs__fill_1 FILLER_0_133_211 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_217 ();
 sky130_as_sc_hs__fill_1 FILLER_0_133_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_246 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_269 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_30 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_300 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_312 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_331 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_337 ();
 sky130_as_sc_hs__fill_1 FILLER_0_133_341 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_362 ();
 sky130_as_sc_hs__fill_1 FILLER_0_133_366 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_369 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_38 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_403 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_42 ();
 sky130_as_sc_hs__fill_1 FILLER_0_133_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_440 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_444 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_449 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_489 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_498 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_505 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_511 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_544 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_553 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_557 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_599 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_603 ();
 sky130_as_sc_hs__fill_1 FILLER_0_133_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_62 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_638 ();
 sky130_as_sc_hs__fill_1 FILLER_0_133_66 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_673 ();
 sky130_as_sc_hs__fill_1 FILLER_0_133_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_707 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_754 ();
 sky130_as_sc_hs__fill_1 FILLER_0_133_758 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_767 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_778 ();
 sky130_as_sc_hs__fill_1 FILLER_0_133_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_805 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_822 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_826 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_833 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_860 ();
 sky130_as_sc_hs__fill_2 FILLER_0_133_864 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_868 ();
 sky130_as_sc_hs__fill_8 FILLER_0_133_884 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_892 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_133_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_133_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_133_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_1013 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_102 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_134_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_1037 ();
 sky130_as_sc_hs__fill_8 FILLER_0_134_1053 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_1061 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_1071 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_1087 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_1091 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_1093 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_1097 ();
 sky130_as_sc_hs__decap_3 FILLER_0_134_11 ();
 sky130_as_sc_hs__decap_3 FILLER_0_134_111 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_1121 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_134_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_1165 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_1181 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_1185 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_119 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_1192 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_1196 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_1203 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_1215 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_1231 ();
 sky130_as_sc_hs__fill_8 FILLER_0_134_1247 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_1255 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_1259 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_130 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_134 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_154 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_170 ();
 sky130_as_sc_hs__fill_8 FILLER_0_134_186 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_194 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_21 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_226 ();
 sky130_as_sc_hs__decap_3 FILLER_0_134_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_264 ();
 sky130_as_sc_hs__decap_3 FILLER_0_134_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_314 ();
 sky130_as_sc_hs__decap_3 FILLER_0_134_323 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_345 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_360 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_365 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_374 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_378 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_397 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_421 ();
 sky130_as_sc_hs__decap_3 FILLER_0_134_44 ();
 sky130_as_sc_hs__decap_3 FILLER_0_134_446 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_451 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_474 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_134_483 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_512 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_52 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_559 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_56 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_563 ();
 sky130_as_sc_hs__decap_3 FILLER_0_134_567 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_583 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_587 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_60 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_64 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_642 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_688 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_692 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_696 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_70 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_746 ();
 sky130_as_sc_hs__fill_1 FILLER_0_134_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_873 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_905 ();
 sky130_as_sc_hs__decap_3 FILLER_0_134_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_94 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_134_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_134_977 ();
 sky130_as_sc_hs__fill_2 FILLER_0_134_98 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_134_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_135_1005 ();
 sky130_as_sc_hs__fill_8 FILLER_0_135_1009 ();
 sky130_as_sc_hs__decap_3 FILLER_0_135_1017 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_106 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_1097 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_110 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_135_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_135_1173 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_1177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_12 ();
 sky130_as_sc_hs__fill_8 FILLER_0_135_1218 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_1226 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_1230 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_135_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_1273 ();
 sky130_as_sc_hs__fill_8 FILLER_0_135_129 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_137 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_146 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_152 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_16 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_163 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_167 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_185 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_20 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_201 ();
 sky130_as_sc_hs__decap_3 FILLER_0_135_205 ();
 sky130_as_sc_hs__fill_8 FILLER_0_135_213 ();
 sky130_as_sc_hs__decap_3 FILLER_0_135_221 ();
 sky130_as_sc_hs__fill_8 FILLER_0_135_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_233 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_237 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_276 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_281 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_285 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_288 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_292 ();
 sky130_as_sc_hs__decap_3 FILLER_0_135_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_135_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_337 ();
 sky130_as_sc_hs__decap_3 FILLER_0_135_371 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_382 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_404 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_41 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_411 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_415 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_423 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_440 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_444 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_449 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_453 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_456 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_460 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_464 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_468 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_472 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_495 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_518 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_52 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_524 ();
 sky130_as_sc_hs__decap_3 FILLER_0_135_557 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_583 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_612 ();
 sky130_as_sc_hs__decap_3 FILLER_0_135_622 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_627 ();
 sky130_as_sc_hs__decap_3 FILLER_0_135_639 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_65 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_655 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_69 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_702 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_706 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_716 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_720 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_724 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_734 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_76 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_775 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_779 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_783 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_8 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_80 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_820 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_824 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_839 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_84 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_859 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_863 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_867 ();
 sky130_as_sc_hs__fill_2 FILLER_0_135_871 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_875 ();
 sky130_as_sc_hs__decap_4 FILLER_0_135_891 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_895 ();
 sky130_as_sc_hs__decap_3 FILLER_0_135_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_90 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_919 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_935 ();
 sky130_as_sc_hs__fill_1 FILLER_0_135_951 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_135_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_136_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_1041 ();
 sky130_as_sc_hs__fill_8 FILLER_0_136_1080 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_1088 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_1093 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_1109 ();
 sky130_as_sc_hs__fill_8 FILLER_0_136_1133 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_136_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_1197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_12 ();
 sky130_as_sc_hs__decap_3 FILLER_0_136_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_1214 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_1230 ();
 sky130_as_sc_hs__fill_8 FILLER_0_136_1246 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_1254 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_136_137 ();
 sky130_as_sc_hs__fill_8 FILLER_0_136_141 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_16 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_163 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_179 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_195 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_20 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_213 ();
 sky130_as_sc_hs__fill_8 FILLER_0_136_229 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_237 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_24 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_241 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_248 ();
 sky130_as_sc_hs__decap_3 FILLER_0_136_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_262 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_29 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_298 ();
 sky130_as_sc_hs__decap_3 FILLER_0_136_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_304 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_323 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_33 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_36 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_362 ();
 sky130_as_sc_hs__decap_3 FILLER_0_136_365 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_381 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_40 ();
 sky130_as_sc_hs__decap_3 FILLER_0_136_417 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_429 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_470 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_485 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_489 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_508 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_528 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_541 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_567 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_587 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_589 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_593 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_596 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_600 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_645 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_657 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_66 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_666 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_686 ();
 sky130_as_sc_hs__decap_3 FILLER_0_136_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_70 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_705 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_709 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_74 ();
 sky130_as_sc_hs__decap_3 FILLER_0_136_753 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_8 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_80 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_817 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_839 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_136_865 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_873 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_877 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_881 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_897 ();
 sky130_as_sc_hs__fill_8 FILLER_0_136_913 ();
 sky130_as_sc_hs__decap_3 FILLER_0_136_921 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_925 ();
 sky130_as_sc_hs__fill_1 FILLER_0_136_929 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_946 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_950 ();
 sky130_as_sc_hs__fill_8 FILLER_0_136_966 ();
 sky130_as_sc_hs__decap_4 FILLER_0_136_974 ();
 sky130_as_sc_hs__fill_2 FILLER_0_136_978 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_136_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_1065 ();
 sky130_as_sc_hs__fill_8 FILLER_0_137_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_1089 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_109 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_1115 ();
 sky130_as_sc_hs__fill_1 FILLER_0_137_1119 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_113 ();
 sky130_as_sc_hs__fill_8 FILLER_0_137_1163 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_1171 ();
 sky130_as_sc_hs__fill_1 FILLER_0_137_1175 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_1229 ();
 sky130_as_sc_hs__fill_8 FILLER_0_137_1233 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_1241 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_1245 ();
 sky130_as_sc_hs__fill_8 FILLER_0_137_1269 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_129 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_13 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_145 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_166 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_17 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_21 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_241 ();
 sky130_as_sc_hs__fill_1 FILLER_0_137_25 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_28 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_290 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_294 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_137_335 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_337 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_34 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_39 ();
 sky130_as_sc_hs__fill_1 FILLER_0_137_391 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_43 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_430 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_445 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_47 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_472 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_481 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_485 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_494 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_500 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_505 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_51 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_511 ();
 sky130_as_sc_hs__fill_1 FILLER_0_137_543 ();
 sky130_as_sc_hs__fill_1 FILLER_0_137_55 ();
 sky130_as_sc_hs__fill_1 FILLER_0_137_561 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_588 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_61 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_611 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_617 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_65 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_669 ();
 sky130_as_sc_hs__fill_1 FILLER_0_137_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_682 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_694 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_720 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_724 ();
 sky130_as_sc_hs__fill_1 FILLER_0_137_729 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_751 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_762 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_797 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_833 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_861 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_865 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_873 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_877 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_137_9 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_137_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_137_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_969 ();
 sky130_as_sc_hs__fill_8 FILLER_0_137_97 ();
 sky130_as_sc_hs__decap_16 FILLER_0_137_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_1033 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_1062 ();
 sky130_as_sc_hs__fill_8 FILLER_0_138_1078 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_1086 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_1090 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_1093 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_11 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_1145 ();
 sky130_as_sc_hs__fill_8 FILLER_0_138_1149 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_1157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_1164 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_1180 ();
 sky130_as_sc_hs__fill_8 FILLER_0_138_1196 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_15 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_172 ();
 sky130_as_sc_hs__fill_8 FILLER_0_138_188 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_20 ();
 sky130_as_sc_hs__fill_8 FILLER_0_138_213 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_24 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_248 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_273 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_29 ();
 sky130_as_sc_hs__fill_8 FILLER_0_138_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_304 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_309 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_328 ();
 sky130_as_sc_hs__fill_1 FILLER_0_138_33 ();
 sky130_as_sc_hs__fill_1 FILLER_0_138_332 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_335 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_339 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_343 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_347 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_36 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_361 ();
 sky130_as_sc_hs__fill_1 FILLER_0_138_365 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_401 ();
 sky130_as_sc_hs__fill_1 FILLER_0_138_405 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_41 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_416 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_435 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_138_456 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_470 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_49 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_501 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_525 ();
 sky130_as_sc_hs__fill_1 FILLER_0_138_546 ();
 sky130_as_sc_hs__fill_1 FILLER_0_138_555 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_584 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_589 ();
 sky130_as_sc_hs__fill_1 FILLER_0_138_600 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_609 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_621 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_626 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_630 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_639 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_645 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_65 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_726 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_730 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_734 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_738 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_742 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_746 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_754 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_765 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_783 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_787 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_791 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_795 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_817 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_138_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_865 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_138_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_138_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_138_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_1002 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_1006 ();
 sky130_as_sc_hs__fill_1 FILLER_0_139_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_1033 ();
 sky130_as_sc_hs__fill_8 FILLER_0_139_1049 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_139_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_185 ();
 sky130_as_sc_hs__fill_8 FILLER_0_139_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_257 ();
 sky130_as_sc_hs__fill_1 FILLER_0_139_279 ();
 sky130_as_sc_hs__fill_8 FILLER_0_139_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_326 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_332 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_337 ();
 sky130_as_sc_hs__fill_1 FILLER_0_139_341 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_344 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_348 ();
 sky130_as_sc_hs__fill_1 FILLER_0_139_37 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_371 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_387 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_40 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_428 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_454 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_501 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_510 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_535 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_553 ();
 sky130_as_sc_hs__fill_1 FILLER_0_139_557 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_569 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_574 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_605 ();
 sky130_as_sc_hs__fill_1 FILLER_0_139_625 ();
 sky130_as_sc_hs__fill_1 FILLER_0_139_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_667 ();
 sky130_as_sc_hs__fill_1 FILLER_0_139_671 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_689 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_710 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_721 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_725 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_761 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_779 ();
 sky130_as_sc_hs__fill_1 FILLER_0_139_783 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_820 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_824 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_828 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_836 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_859 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_863 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_867 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_871 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_875 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_89 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_891 ();
 sky130_as_sc_hs__fill_1 FILLER_0_139_895 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_139_949 ();
 sky130_as_sc_hs__fill_8 FILLER_0_139_953 ();
 sky130_as_sc_hs__decap_4 FILLER_0_139_961 ();
 sky130_as_sc_hs__fill_2 FILLER_0_139_965 ();
 sky130_as_sc_hs__decap_16 FILLER_0_139_986 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_1002 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_1006 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1025 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_103 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1065 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_108 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1121 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1177 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1233 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_124 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_13_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_128 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_132 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_136 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_140 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_144 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_148 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_152 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_225 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_241 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_257 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_292 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_370 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_386 ();
 sky130_as_sc_hs__fill_1 FILLER_0_13_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_399 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_434 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_449 ();
 sky130_as_sc_hs__fill_1 FILLER_0_13_465 ();
 sky130_as_sc_hs__fill_1 FILLER_0_13_471 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_490 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_502 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_51 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_510 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_533 ();
 sky130_as_sc_hs__fill_1 FILLER_0_13_543 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_549 ();
 sky130_as_sc_hs__fill_1 FILLER_0_13_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_558 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_588 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_603 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_13_666 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_700 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_708 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_729 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_733 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_748 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_752 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_756 ();
 sky130_as_sc_hs__fill_1 FILLER_0_13_771 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_79 ();
 sky130_as_sc_hs__fill_1 FILLER_0_13_805 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_83 ();
 sky130_as_sc_hs__fill_1 FILLER_0_13_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_849 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_870 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_88 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_910 ();
 sky130_as_sc_hs__decap_4 FILLER_0_13_93 ();
 sky130_as_sc_hs__decap_3 FILLER_0_13_935 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_958 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_962 ();
 sky130_as_sc_hs__decap_16 FILLER_0_13_978 ();
 sky130_as_sc_hs__fill_2 FILLER_0_13_99 ();
 sky130_as_sc_hs__fill_8 FILLER_0_13_994 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_1004 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_1020 ();
 sky130_as_sc_hs__decap_4 FILLER_0_140_1037 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_1041 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_1066 ();
 sky130_as_sc_hs__fill_8 FILLER_0_140_1082 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_1090 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_140_1141 ();
 sky130_as_sc_hs__fill_1 FILLER_0_140_1145 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_117 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_1176 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_1188 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_140_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_140_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_140_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_140_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_140_213 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_221 ();
 sky130_as_sc_hs__fill_1 FILLER_0_140_243 ();
 sky130_as_sc_hs__fill_1 FILLER_0_140_258 ();
 sky130_as_sc_hs__fill_1 FILLER_0_140_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_283 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_325 ();
 sky130_as_sc_hs__decap_4 FILLER_0_140_353 ();
 sky130_as_sc_hs__fill_1 FILLER_0_140_357 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_384 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_407 ();
 sky130_as_sc_hs__fill_1 FILLER_0_140_419 ();
 sky130_as_sc_hs__fill_1 FILLER_0_140_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_140_438 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_458 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_468 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_472 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_522 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_557 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_580 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_610 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_622 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_630 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_634 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_664 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_697 ();
 sky130_as_sc_hs__fill_1 FILLER_0_140_706 ();
 sky130_as_sc_hs__fill_1 FILLER_0_140_755 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_757 ();
 sky130_as_sc_hs__decap_4 FILLER_0_140_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_789 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_793 ();
 sky130_as_sc_hs__fill_1 FILLER_0_140_801 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_837 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_852 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_856 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_860 ();
 sky130_as_sc_hs__fill_2 FILLER_0_140_864 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_140_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_140_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_977 ();
 sky130_as_sc_hs__decap_3 FILLER_0_140_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_140_988 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_1002 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_1006 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_1009 ();
 sky130_as_sc_hs__fill_8 FILLER_0_141_1025 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_1033 ();
 sky130_as_sc_hs__fill_8 FILLER_0_141_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_1049 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_105 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_1053 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_141_1061 ();
 sky130_as_sc_hs__fill_8 FILLER_0_141_1065 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_1073 ();
 sky130_as_sc_hs__decap_3 FILLER_0_141_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_1094 ();
 sky130_as_sc_hs__fill_8 FILLER_0_141_1110 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_1118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_141_1173 ();
 sky130_as_sc_hs__decap_3 FILLER_0_141_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_1196 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_1212 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_1228 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_141_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_141_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_141_221 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_231 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_235 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_243 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_260 ();
 sky130_as_sc_hs__fill_1 FILLER_0_141_264 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_299 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_141_303 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_306 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_310 ();
 sky130_as_sc_hs__decap_3 FILLER_0_141_314 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_35 ();
 sky130_as_sc_hs__fill_1 FILLER_0_141_363 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_388 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_393 ();
 sky130_as_sc_hs__fill_1 FILLER_0_141_397 ();
 sky130_as_sc_hs__decap_3 FILLER_0_141_439 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_444 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_470 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_493 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_500 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_141_524 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_542 ();
 sky130_as_sc_hs__fill_1 FILLER_0_141_55 ();
 sky130_as_sc_hs__decap_3 FILLER_0_141_557 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_569 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_573 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_612 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_141_678 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_684 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_688 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_692 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_696 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_700 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_707 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_714 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_718 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_722 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_726 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_73 ();
 sky130_as_sc_hs__decap_3 FILLER_0_141_733 ();
 sky130_as_sc_hs__decap_3 FILLER_0_141_744 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_795 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_799 ();
 sky130_as_sc_hs__fill_1 FILLER_0_141_803 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_814 ();
 sky130_as_sc_hs__decap_3 FILLER_0_141_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_846 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_850 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_854 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_858 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_862 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_878 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_89 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_894 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_141_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_141_953 ();
 sky130_as_sc_hs__fill_8 FILLER_0_141_969 ();
 sky130_as_sc_hs__decap_4 FILLER_0_141_977 ();
 sky130_as_sc_hs__fill_1 FILLER_0_141_981 ();
 sky130_as_sc_hs__fill_2 FILLER_0_141_998 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_101 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_1014 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_1037 ();
 sky130_as_sc_hs__fill_1 FILLER_0_142_1055 ();
 sky130_as_sc_hs__fill_8 FILLER_0_142_1079 ();
 sky130_as_sc_hs__decap_4 FILLER_0_142_1087 ();
 sky130_as_sc_hs__fill_1 FILLER_0_142_1091 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_1097 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_1101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_1117 ();
 sky130_as_sc_hs__fill_8 FILLER_0_142_1133 ();
 sky130_as_sc_hs__decap_4 FILLER_0_142_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_1145 ();
 sky130_as_sc_hs__fill_8 FILLER_0_142_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_117 ();
 sky130_as_sc_hs__decap_4 FILLER_0_142_1175 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_1179 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_1187 ();
 sky130_as_sc_hs__fill_1 FILLER_0_142_1203 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_142_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_1257 ();
 sky130_as_sc_hs__fill_8 FILLER_0_142_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_142_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_142_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_142_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_142_213 ();
 sky130_as_sc_hs__decap_4 FILLER_0_142_221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_244 ();
 sky130_as_sc_hs__decap_4 FILLER_0_142_266 ();
 sky130_as_sc_hs__fill_1 FILLER_0_142_27 ();
 sky130_as_sc_hs__fill_1 FILLER_0_142_270 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_289 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_142_307 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_313 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_317 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_321 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_325 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_330 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_334 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_338 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_342 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_354 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_361 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_370 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_392 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_397 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_434 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_457 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_471 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_481 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_485 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_489 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_512 ();
 sky130_as_sc_hs__fill_1 FILLER_0_142_544 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_566 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_570 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_574 ();
 sky130_as_sc_hs__fill_1 FILLER_0_142_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_603 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_625 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_629 ();
 sky130_as_sc_hs__decap_4 FILLER_0_142_634 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_640 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_669 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_677 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_689 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_709 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_713 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_726 ();
 sky130_as_sc_hs__decap_4 FILLER_0_142_77 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_783 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_805 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_809 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_818 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_822 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_826 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_830 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_834 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_842 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_846 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_850 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_854 ();
 sky130_as_sc_hs__fill_8 FILLER_0_142_858 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_866 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_142_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_142_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_142_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_142_977 ();
 sky130_as_sc_hs__fill_8 FILLER_0_142_981 ();
 sky130_as_sc_hs__decap_4 FILLER_0_142_989 ();
 sky130_as_sc_hs__fill_2 FILLER_0_142_993 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_1005 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_1015 ();
 sky130_as_sc_hs__fill_8 FILLER_0_143_1031 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_1039 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_105 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_1061 ();
 sky130_as_sc_hs__fill_8 FILLER_0_143_1065 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_1073 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_109 ();
 sky130_as_sc_hs__fill_8 FILLER_0_143_1112 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_143_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_217 ();
 sky130_as_sc_hs__fill_1 FILLER_0_143_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_246 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_143_277 ();
 sky130_as_sc_hs__fill_1 FILLER_0_143_289 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_344 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_364 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_404 ();
 sky130_as_sc_hs__fill_1 FILLER_0_143_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_440 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_444 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_449 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_459 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_465 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_488 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_499 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_51 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_519 ();
 sky130_as_sc_hs__fill_1 FILLER_0_143_523 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_545 ();
 sky130_as_sc_hs__fill_1 FILLER_0_143_55 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_569 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_143_610 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_622 ();
 sky130_as_sc_hs__fill_8 FILLER_0_143_626 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_634 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_638 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_642 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_646 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_670 ();
 sky130_as_sc_hs__fill_1 FILLER_0_143_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_698 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_702 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_724 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_73 ();
 sky130_as_sc_hs__fill_1 FILLER_0_143_745 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_846 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_850 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_854 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_858 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_862 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_866 ();
 sky130_as_sc_hs__fill_8 FILLER_0_143_882 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_89 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_890 ();
 sky130_as_sc_hs__fill_2 FILLER_0_143_894 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_143_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_143_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_143_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_1037 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_1053 ();
 sky130_as_sc_hs__fill_1 FILLER_0_144_1057 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_1062 ();
 sky130_as_sc_hs__fill_8 FILLER_0_144_1078 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_1086 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_1090 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_1093 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_1100 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_1104 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_1129 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_1149 ();
 sky130_as_sc_hs__fill_8 FILLER_0_144_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_117 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_1173 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_1184 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_1200 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_1257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_1261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_1265 ();
 sky130_as_sc_hs__fill_1 FILLER_0_144_1276 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_144_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_144_213 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_221 ();
 sky130_as_sc_hs__fill_1 FILLER_0_144_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_228 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_232 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_236 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_240 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_248 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_266 ();
 sky130_as_sc_hs__fill_1 FILLER_0_144_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_270 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_282 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_287 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_291 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_295 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_299 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_322 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_349 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_362 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_365 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_386 ();
 sky130_as_sc_hs__fill_1 FILLER_0_144_390 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_404 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_416 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_421 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_432 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_45 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_469 ();
 sky130_as_sc_hs__fill_1 FILLER_0_144_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_510 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_525 ();
 sky130_as_sc_hs__fill_1 FILLER_0_144_529 ();
 sky130_as_sc_hs__fill_1 FILLER_0_144_552 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_574 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_578 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_582 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_589 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_61 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_628 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_636 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_640 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_664 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_676 ();
 sky130_as_sc_hs__fill_1 FILLER_0_144_680 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_709 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_713 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_757 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_790 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_794 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_798 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_802 ();
 sky130_as_sc_hs__fill_1 FILLER_0_144_806 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_813 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_865 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_144_873 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_877 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_893 ();
 sky130_as_sc_hs__fill_8 FILLER_0_144_909 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_144_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_944 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_960 ();
 sky130_as_sc_hs__decap_4 FILLER_0_144_976 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_144_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_145_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_145_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_1009 ();
 sky130_as_sc_hs__fill_1 FILLER_0_145_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_1045 ();
 sky130_as_sc_hs__decap_4 FILLER_0_145_105 ();
 sky130_as_sc_hs__decap_3 FILLER_0_145_1061 ();
 sky130_as_sc_hs__decap_3 FILLER_0_145_1088 ();
 sky130_as_sc_hs__decap_3 FILLER_0_145_109 ();
 sky130_as_sc_hs__decap_4 FILLER_0_145_1096 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_1100 ();
 sky130_as_sc_hs__decap_4 FILLER_0_145_1106 ();
 sky130_as_sc_hs__fill_1 FILLER_0_145_1110 ();
 sky130_as_sc_hs__decap_4 FILLER_0_145_1116 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_1126 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_1142 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_1158 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_1174 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_145_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_145_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_1233 ();
 sky130_as_sc_hs__fill_8 FILLER_0_145_1249 ();
 sky130_as_sc_hs__decap_4 FILLER_0_145_1257 ();
 sky130_as_sc_hs__decap_3 FILLER_0_145_1274 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_145_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_145_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_145_217 ();
 sky130_as_sc_hs__fill_1 FILLER_0_145_221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_145_225 ();
 sky130_as_sc_hs__fill_1 FILLER_0_145_247 ();
 sky130_as_sc_hs__decap_4 FILLER_0_145_266 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_145_304 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_313 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_361 ();
 sky130_as_sc_hs__fill_1 FILLER_0_145_391 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_393 ();
 sky130_as_sc_hs__decap_4 FILLER_0_145_405 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_411 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_415 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_419 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_423 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_446 ();
 sky130_as_sc_hs__fill_1 FILLER_0_145_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_466 ();
 sky130_as_sc_hs__fill_1 FILLER_0_145_487 ();
 sky130_as_sc_hs__fill_1 FILLER_0_145_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_145_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_530 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_534 ();
 sky130_as_sc_hs__fill_1 FILLER_0_145_55 ();
 sky130_as_sc_hs__decap_3 FILLER_0_145_557 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_571 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_575 ();
 sky130_as_sc_hs__decap_3 FILLER_0_145_579 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_606 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_610 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_614 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_649 ();
 sky130_as_sc_hs__fill_1 FILLER_0_145_661 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_681 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_685 ();
 sky130_as_sc_hs__fill_1 FILLER_0_145_727 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_753 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_761 ();
 sky130_as_sc_hs__fill_1 FILLER_0_145_773 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_797 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_801 ();
 sky130_as_sc_hs__decap_3 FILLER_0_145_816 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_861 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_865 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_145_873 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_877 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_145_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_145_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_145_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_145_985 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_1005 ();
 sky130_as_sc_hs__fill_1 FILLER_0_146_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_101 ();
 sky130_as_sc_hs__decap_3 FILLER_0_146_1033 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_1037 ();
 sky130_as_sc_hs__fill_1 FILLER_0_146_1041 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_1046 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_1062 ();
 sky130_as_sc_hs__fill_8 FILLER_0_146_1078 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_1086 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_1090 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_1132 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_146_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_146_1257 ();
 sky130_as_sc_hs__fill_8 FILLER_0_146_1261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_146_1274 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_146_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_146_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_146_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_146_213 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_221 ();
 sky130_as_sc_hs__fill_1 FILLER_0_146_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_265 ();
 sky130_as_sc_hs__fill_1 FILLER_0_146_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_277 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_289 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_295 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_299 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_325 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_331 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_348 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_362 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_400 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_404 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_416 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_440 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_146_450 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_472 ();
 sky130_as_sc_hs__decap_3 FILLER_0_146_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_525 ();
 sky130_as_sc_hs__decap_3 FILLER_0_146_529 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_533 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_537 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_543 ();
 sky130_as_sc_hs__decap_3 FILLER_0_146_566 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_571 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_601 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_605 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_626 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_630 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_642 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_653 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_695 ();
 sky130_as_sc_hs__fill_1 FILLER_0_146_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_733 ();
 sky130_as_sc_hs__fill_1 FILLER_0_146_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_763 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_77 ();
 sky130_as_sc_hs__decap_3 FILLER_0_146_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_825 ();
 sky130_as_sc_hs__fill_1 FILLER_0_146_829 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_854 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_858 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_862 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_866 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_146_873 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_877 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_893 ();
 sky130_as_sc_hs__fill_8 FILLER_0_146_909 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_146_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_146_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_146_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_146_981 ();
 sky130_as_sc_hs__fill_8 FILLER_0_146_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_147_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_1009 ();
 sky130_as_sc_hs__fill_8 FILLER_0_147_1025 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_1033 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_1037 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_105 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_147_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_147_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_1126 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_113 ();
 sky130_as_sc_hs__fill_8 FILLER_0_147_1142 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_1150 ();
 sky130_as_sc_hs__decap_3 FILLER_0_147_1154 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_147_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_1249 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_1265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_1275 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_147_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_147_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_233 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_237 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_241 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_245 ();
 sky130_as_sc_hs__decap_3 FILLER_0_147_257 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_278 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_281 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_299 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_313 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_353 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_363 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_390 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_398 ();
 sky130_as_sc_hs__fill_1 FILLER_0_147_402 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_405 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_409 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_413 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_436 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_484 ();
 sky130_as_sc_hs__fill_1 FILLER_0_147_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_51 ();
 sky130_as_sc_hs__decap_3 FILLER_0_147_527 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_532 ();
 sky130_as_sc_hs__fill_1 FILLER_0_147_546 ();
 sky130_as_sc_hs__fill_1 FILLER_0_147_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_552 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_556 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_147_584 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_609 ();
 sky130_as_sc_hs__fill_1 FILLER_0_147_613 ();
 sky130_as_sc_hs__decap_3 FILLER_0_147_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_656 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_660 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_664 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_668 ();
 sky130_as_sc_hs__fill_1 FILLER_0_147_681 ();
 sky130_as_sc_hs__decap_3 FILLER_0_147_725 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_747 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_793 ();
 sky130_as_sc_hs__fill_1 FILLER_0_147_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_854 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_858 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_862 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_866 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_870 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_874 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_878 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_882 ();
 sky130_as_sc_hs__fill_8 FILLER_0_147_886 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_89 ();
 sky130_as_sc_hs__fill_2 FILLER_0_147_894 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_147_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_147_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_147_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_1004 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_1020 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_1037 ();
 sky130_as_sc_hs__decap_4 FILLER_0_148_1053 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_1057 ();
 sky130_as_sc_hs__fill_8 FILLER_0_148_1082 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_1090 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_148_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_1149 ();
 sky130_as_sc_hs__fill_1 FILLER_0_148_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_117 ();
 sky130_as_sc_hs__fill_1 FILLER_0_148_1171 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_1177 ();
 sky130_as_sc_hs__fill_8 FILLER_0_148_1193 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_148_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_1257 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_1274 ();
 sky130_as_sc_hs__decap_4 FILLER_0_148_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_148_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_148_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_148_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_247 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_253 ();
 sky130_as_sc_hs__fill_1 FILLER_0_148_27 ();
 sky130_as_sc_hs__fill_1 FILLER_0_148_276 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_29 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_290 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_148_317 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_342 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_384 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_407 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_416 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_450 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_482 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_492 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_560 ();
 sky130_as_sc_hs__fill_1 FILLER_0_148_582 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_605 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_610 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_614 ();
 sky130_as_sc_hs__decap_4 FILLER_0_148_634 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_640 ();
 sky130_as_sc_hs__fill_1 FILLER_0_148_674 ();
 sky130_as_sc_hs__fill_1 FILLER_0_148_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_714 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_754 ();
 sky130_as_sc_hs__decap_4 FILLER_0_148_77 ();
 sky130_as_sc_hs__fill_1 FILLER_0_148_781 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_809 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_865 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_148_873 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_877 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_893 ();
 sky130_as_sc_hs__fill_8 FILLER_0_148_909 ();
 sky130_as_sc_hs__decap_4 FILLER_0_148_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_148_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_148_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_148_977 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_1032 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_1048 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_105 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_1137 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_1172 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_1190 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_1206 ();
 sky130_as_sc_hs__fill_8 FILLER_0_149_1222 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_1230 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_1249 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_333 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_35 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_353 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_359 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_363 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_367 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_371 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_375 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_379 ();
 sky130_as_sc_hs__fill_1 FILLER_0_149_391 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_393 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_414 ();
 sky130_as_sc_hs__fill_1 FILLER_0_149_438 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_444 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_462 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_484 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_51 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_526 ();
 sky130_as_sc_hs__fill_1 FILLER_0_149_530 ();
 sky130_as_sc_hs__fill_1 FILLER_0_149_546 ();
 sky130_as_sc_hs__fill_1 FILLER_0_149_55 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_555 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_149_646 ();
 sky130_as_sc_hs__fill_1 FILLER_0_149_655 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_673 ();
 sky130_as_sc_hs__fill_1 FILLER_0_149_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_724 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_73 ();
 sky130_as_sc_hs__fill_1 FILLER_0_149_801 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_834 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_861 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_865 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_873 ();
 sky130_as_sc_hs__fill_2 FILLER_0_149_877 ();
 sky130_as_sc_hs__fill_8 FILLER_0_149_881 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_149_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_149_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_149_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1013 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_102 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1053 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_106 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1093 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_110 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1125 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_114 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1165 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1205 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_122 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_1257 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_126 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_130 ();
 sky130_as_sc_hs__fill_1 FILLER_0_14_134 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_137 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_145 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_153 ();
 sky130_as_sc_hs__fill_8 FILLER_0_14_157 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_165 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_171 ();
 sky130_as_sc_hs__fill_8 FILLER_0_14_176 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_186 ();
 sky130_as_sc_hs__fill_8 FILLER_0_14_19 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_190 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_194 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_213 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_229 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_245 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_249 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_253 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_269 ();
 sky130_as_sc_hs__fill_1 FILLER_0_14_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_316 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_330 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_338 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_365 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_397 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_421 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_463 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_472 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_482 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_510 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_556 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_572 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_597 ();
 sky130_as_sc_hs__fill_8 FILLER_0_14_61 ();
 sky130_as_sc_hs__fill_1 FILLER_0_14_620 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_634 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_642 ();
 sky130_as_sc_hs__fill_1 FILLER_0_14_672 ();
 sky130_as_sc_hs__fill_1 FILLER_0_14_69 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_711 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_72 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_76 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_80 ();
 sky130_as_sc_hs__fill_1 FILLER_0_14_811 ();
 sky130_as_sc_hs__fill_1 FILLER_0_14_832 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_854 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_858 ();
 sky130_as_sc_hs__decap_4 FILLER_0_14_862 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_89 ();
 sky130_as_sc_hs__fill_1 FILLER_0_14_892 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_921 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_925 ();
 sky130_as_sc_hs__fill_1 FILLER_0_14_929 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_93 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_953 ();
 sky130_as_sc_hs__fill_8 FILLER_0_14_969 ();
 sky130_as_sc_hs__decap_3 FILLER_0_14_977 ();
 sky130_as_sc_hs__fill_2 FILLER_0_14_98 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_14_997 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_150_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_150_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_1060 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_1076 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_1132 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_1149 ();
 sky130_as_sc_hs__decap_4 FILLER_0_150_1165 ();
 sky130_as_sc_hs__fill_1 FILLER_0_150_1169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_117 ();
 sky130_as_sc_hs__fill_8 FILLER_0_150_1175 ();
 sky130_as_sc_hs__decap_4 FILLER_0_150_1183 ();
 sky130_as_sc_hs__fill_1 FILLER_0_150_1187 ();
 sky130_as_sc_hs__fill_8 FILLER_0_150_1193 ();
 sky130_as_sc_hs__decap_3 FILLER_0_150_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_150_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_150_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_150_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_150_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_150_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_150_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_150_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_197 ();
 sky130_as_sc_hs__decap_4 FILLER_0_150_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_238 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_245 ();
 sky130_as_sc_hs__decap_4 FILLER_0_150_261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_150_265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_268 ();
 sky130_as_sc_hs__fill_1 FILLER_0_150_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_272 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_280 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_150_336 ();
 sky130_as_sc_hs__fill_1 FILLER_0_150_340 ();
 sky130_as_sc_hs__decap_3 FILLER_0_150_351 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_369 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_418 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_150_442 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_467 ();
 sky130_as_sc_hs__fill_1 FILLER_0_150_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_150_510 ();
 sky130_as_sc_hs__fill_1 FILLER_0_150_554 ();
 sky130_as_sc_hs__decap_3 FILLER_0_150_560 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_565 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_629 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_671 ();
 sky130_as_sc_hs__decap_3 FILLER_0_150_697 ();
 sky130_as_sc_hs__decap_3 FILLER_0_150_722 ();
 sky130_as_sc_hs__fill_1 FILLER_0_150_744 ();
 sky130_as_sc_hs__decap_4 FILLER_0_150_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_773 ();
 sky130_as_sc_hs__decap_3 FILLER_0_150_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_818 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_854 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_858 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_862 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_866 ();
 sky130_as_sc_hs__fill_2 FILLER_0_150_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_873 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_905 ();
 sky130_as_sc_hs__decap_3 FILLER_0_150_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_150_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_150_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_150_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_1004 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_1009 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_1013 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_1038 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_105 ();
 sky130_as_sc_hs__fill_8 FILLER_0_151_1054 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_151_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_151_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_151_1173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_1202 ();
 sky130_as_sc_hs__fill_8 FILLER_0_151_1218 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_1226 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_1230 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_151_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_151_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_151_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_249 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_278 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_281 ();
 sky130_as_sc_hs__fill_1 FILLER_0_151_285 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_288 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_292 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_296 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_304 ();
 sky130_as_sc_hs__fill_1 FILLER_0_151_327 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_35 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_355 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_380 ();
 sky130_as_sc_hs__fill_1 FILLER_0_151_414 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_420 ();
 sky130_as_sc_hs__fill_1 FILLER_0_151_424 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_427 ();
 sky130_as_sc_hs__fill_1 FILLER_0_151_447 ();
 sky130_as_sc_hs__fill_1 FILLER_0_151_462 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_500 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_151_55 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_603 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_607 ();
 sky130_as_sc_hs__decap_3 FILLER_0_151_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_151_644 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_664 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_668 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_724 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_754 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_820 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_849 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_861 ();
 sky130_as_sc_hs__fill_2 FILLER_0_151_865 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_869 ();
 sky130_as_sc_hs__fill_8 FILLER_0_151_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_151_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_151_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_151_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_151_953 ();
 sky130_as_sc_hs__fill_8 FILLER_0_151_969 ();
 sky130_as_sc_hs__fill_8 FILLER_0_151_996 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1013 ();
 sky130_as_sc_hs__fill_1 FILLER_0_152_1029 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_1032 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_152_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_152_213 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_221 ();
 sky130_as_sc_hs__fill_1 FILLER_0_152_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_228 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_232 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_269 ();
 sky130_as_sc_hs__fill_1 FILLER_0_152_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_283 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_29 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_292 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_303 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_318 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_340 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_354 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_384 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_418 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_430 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_152_458 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_467 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_496 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_549 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_571 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_581 ();
 sky130_as_sc_hs__fill_1 FILLER_0_152_585 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_61 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_626 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_677 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_752 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_765 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_769 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_77 ();
 sky130_as_sc_hs__fill_1 FILLER_0_152_773 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_795 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_152_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_865 ();
 sky130_as_sc_hs__decap_3 FILLER_0_152_869 ();
 sky130_as_sc_hs__fill_8 FILLER_0_152_891 ();
 sky130_as_sc_hs__fill_1 FILLER_0_152_899 ();
 sky130_as_sc_hs__decap_4 FILLER_0_152_919 ();
 sky130_as_sc_hs__fill_1 FILLER_0_152_923 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_152_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_153_1005 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_1009 ();
 sky130_as_sc_hs__fill_1 FILLER_0_153_1013 ();
 sky130_as_sc_hs__decap_3 FILLER_0_153_1030 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_105 ();
 sky130_as_sc_hs__fill_8 FILLER_0_153_1056 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_1088 ();
 sky130_as_sc_hs__decap_3 FILLER_0_153_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_1104 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_113 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_1156 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_1172 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_1177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_1203 ();
 sky130_as_sc_hs__fill_8 FILLER_0_153_1219 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_1227 ();
 sky130_as_sc_hs__fill_1 FILLER_0_153_1231 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_153_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_153_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_153_221 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_153_229 ();
 sky130_as_sc_hs__fill_1 FILLER_0_153_261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_153_270 ();
 sky130_as_sc_hs__fill_1 FILLER_0_153_279 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_153_304 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_326 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_35 ();
 sky130_as_sc_hs__decap_3 FILLER_0_153_350 ();
 sky130_as_sc_hs__decap_3 FILLER_0_153_372 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_380 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_418 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_441 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_449 ();
 sky130_as_sc_hs__decap_3 FILLER_0_153_485 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_521 ();
 sky130_as_sc_hs__fill_1 FILLER_0_153_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_579 ();
 sky130_as_sc_hs__decap_3 FILLER_0_153_613 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_652 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_681 ();
 sky130_as_sc_hs__fill_1 FILLER_0_153_685 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_715 ();
 sky130_as_sc_hs__decap_3 FILLER_0_153_725 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_73 ();
 sky130_as_sc_hs__fill_1 FILLER_0_153_771 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_809 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_817 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_828 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_832 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_836 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_849 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_153_861 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_865 ();
 sky130_as_sc_hs__fill_8 FILLER_0_153_881 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_153_893 ();
 sky130_as_sc_hs__decap_4 FILLER_0_153_897 ();
 sky130_as_sc_hs__fill_1 FILLER_0_153_901 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_920 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_936 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_153_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_1012 ();
 sky130_as_sc_hs__fill_8 FILLER_0_154_1028 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_154_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_154_1089 ();
 sky130_as_sc_hs__fill_8 FILLER_0_154_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_1119 ();
 sky130_as_sc_hs__fill_1 FILLER_0_154_1135 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_1146 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_1168 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_117 ();
 sky130_as_sc_hs__decap_4 FILLER_0_154_1184 ();
 sky130_as_sc_hs__decap_3 FILLER_0_154_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_1210 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_1226 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_1242 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_1258 ();
 sky130_as_sc_hs__decap_4 FILLER_0_154_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_1265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_1275 ();
 sky130_as_sc_hs__decap_4 FILLER_0_154_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_154_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_154_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_154_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_154_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_154_213 ();
 sky130_as_sc_hs__decap_4 FILLER_0_154_221 ();
 sky130_as_sc_hs__fill_1 FILLER_0_154_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_250 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_253 ();
 sky130_as_sc_hs__fill_1 FILLER_0_154_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_154_303 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_392 ();
 sky130_as_sc_hs__fill_1 FILLER_0_154_413 ();
 sky130_as_sc_hs__fill_1 FILLER_0_154_419 ();
 sky130_as_sc_hs__decap_3 FILLER_0_154_429 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_434 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_154_470 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_154_529 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_544 ();
 sky130_as_sc_hs__decap_3 FILLER_0_154_556 ();
 sky130_as_sc_hs__fill_1 FILLER_0_154_608 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_650 ();
 sky130_as_sc_hs__fill_1 FILLER_0_154_668 ();
 sky130_as_sc_hs__decap_3 FILLER_0_154_688 ();
 sky130_as_sc_hs__fill_1 FILLER_0_154_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_701 ();
 sky130_as_sc_hs__fill_1 FILLER_0_154_757 ();
 sky130_as_sc_hs__decap_4 FILLER_0_154_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_792 ();
 sky130_as_sc_hs__decap_3 FILLER_0_154_809 ();
 sky130_as_sc_hs__decap_3 FILLER_0_154_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_154_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_857 ();
 sky130_as_sc_hs__decap_4 FILLER_0_154_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_154_865 ();
 sky130_as_sc_hs__decap_4 FILLER_0_154_869 ();
 sky130_as_sc_hs__fill_1 FILLER_0_154_873 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_887 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_903 ();
 sky130_as_sc_hs__decap_4 FILLER_0_154_919 ();
 sky130_as_sc_hs__fill_1 FILLER_0_154_923 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_154_941 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_957 ();
 sky130_as_sc_hs__fill_2 FILLER_0_154_978 ();
 sky130_as_sc_hs__fill_8 FILLER_0_154_985 ();
 sky130_as_sc_hs__fill_1 FILLER_0_155_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_1033 ();
 sky130_as_sc_hs__fill_8 FILLER_0_155_1049 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_1061 ();
 sky130_as_sc_hs__fill_8 FILLER_0_155_1065 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_1073 ();
 sky130_as_sc_hs__fill_1 FILLER_0_155_1077 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_113 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_1152 ();
 sky130_as_sc_hs__fill_8 FILLER_0_155_1168 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_155_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_225 ();
 sky130_as_sc_hs__fill_1 FILLER_0_155_247 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_25 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_259 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_263 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_276 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_286 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_297 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_302 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_306 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_310 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_318 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_322 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_345 ();
 sky130_as_sc_hs__fill_1 FILLER_0_155_349 ();
 sky130_as_sc_hs__fill_1 FILLER_0_155_371 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_390 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_401 ();
 sky130_as_sc_hs__fill_1 FILLER_0_155_405 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_408 ();
 sky130_as_sc_hs__fill_8 FILLER_0_155_41 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_425 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_438 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_444 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_454 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_458 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_462 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_49 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_53 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_537 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_556 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_577 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_595 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_604 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_608 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_612 ();
 sky130_as_sc_hs__fill_1 FILLER_0_155_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_626 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_641 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_646 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_665 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_673 ();
 sky130_as_sc_hs__fill_1 FILLER_0_155_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_726 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_742 ();
 sky130_as_sc_hs__decap_3 FILLER_0_155_763 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_805 ();
 sky130_as_sc_hs__fill_1 FILLER_0_155_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_851 ();
 sky130_as_sc_hs__fill_2 FILLER_0_155_855 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_859 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_875 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_89 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_891 ();
 sky130_as_sc_hs__fill_1 FILLER_0_155_895 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_9 ();
 sky130_as_sc_hs__decap_16 FILLER_0_155_913 ();
 sky130_as_sc_hs__decap_4 FILLER_0_155_929 ();
 sky130_as_sc_hs__fill_8 FILLER_0_155_996 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_1004 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_1020 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_1064 ();
 sky130_as_sc_hs__fill_8 FILLER_0_156_1080 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_1088 ();
 sky130_as_sc_hs__fill_1 FILLER_0_156_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_1098 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_1114 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_1118 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_1126 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_1134 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_1154 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_117 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_1170 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_1174 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_1182 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_1198 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_1202 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_189 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_213 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_229 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_23 ();
 sky130_as_sc_hs__fill_1 FILLER_0_156_253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_267 ();
 sky130_as_sc_hs__fill_1 FILLER_0_156_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_289 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_29 ();
 sky130_as_sc_hs__fill_1 FILLER_0_156_307 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_318 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_322 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_353 ();
 sky130_as_sc_hs__fill_1 FILLER_0_156_357 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_360 ();
 sky130_as_sc_hs__fill_1 FILLER_0_156_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_408 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_440 ();
 sky130_as_sc_hs__fill_1 FILLER_0_156_444 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_447 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_451 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_455 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_469 ();
 sky130_as_sc_hs__fill_1 FILLER_0_156_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_481 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_501 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_513 ();
 sky130_as_sc_hs__fill_1 FILLER_0_156_531 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_533 ();
 sky130_as_sc_hs__fill_1 FILLER_0_156_551 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_576 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_586 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_605 ();
 sky130_as_sc_hs__fill_1 FILLER_0_156_609 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_612 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_624 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_642 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_649 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_685 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_697 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_749 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_753 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_77 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_156_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_842 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_854 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_858 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_862 ();
 sky130_as_sc_hs__fill_2 FILLER_0_156_866 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_156_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_156_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_156_975 ();
 sky130_as_sc_hs__fill_1 FILLER_0_156_979 ();
 sky130_as_sc_hs__decap_3 FILLER_0_157_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_1016 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_1032 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_1048 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_105 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_1065 ();
 sky130_as_sc_hs__fill_8 FILLER_0_157_1081 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_1089 ();
 sky130_as_sc_hs__decap_3 FILLER_0_157_109 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_1116 ();
 sky130_as_sc_hs__fill_8 FILLER_0_157_1121 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_1129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_157_1133 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_1141 ();
 sky130_as_sc_hs__fill_8 FILLER_0_157_1157 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_1165 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_1169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_157_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_157_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_157_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_157_221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_225 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_241 ();
 sky130_as_sc_hs__fill_1 FILLER_0_157_245 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_248 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_252 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_264 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_268 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_272 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_276 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_305 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_313 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_35 ();
 sky130_as_sc_hs__decap_3 FILLER_0_157_371 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_390 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_438 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_444 ();
 sky130_as_sc_hs__decap_3 FILLER_0_157_473 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_157_524 ();
 sky130_as_sc_hs__fill_1 FILLER_0_157_55 ();
 sky130_as_sc_hs__decap_3 FILLER_0_157_557 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_157_588 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_610 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_157_621 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_640 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_668 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_692 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_720 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_724 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_73 ();
 sky130_as_sc_hs__decap_3 FILLER_0_157_753 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_795 ();
 sky130_as_sc_hs__decap_3 FILLER_0_157_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_861 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_865 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_873 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_157_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_157_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_919 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_935 ();
 sky130_as_sc_hs__fill_1 FILLER_0_157_951 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_157_969 ();
 sky130_as_sc_hs__decap_4 FILLER_0_157_985 ();
 sky130_as_sc_hs__fill_8 FILLER_0_158_1000 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_1008 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_101 ();
 sky130_as_sc_hs__fill_1 FILLER_0_158_1035 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_1037 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_1041 ();
 sky130_as_sc_hs__fill_8 FILLER_0_158_1082 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_1090 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_1257 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_1266 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_158_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_158_213 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_247 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_253 ();
 sky130_as_sc_hs__fill_1 FILLER_0_158_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_280 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_284 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_293 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_297 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_158_301 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_304 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_318 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_322 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_326 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_330 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_334 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_356 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_410 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_416 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_434 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_439 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_158_470 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_158_496 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_516 ();
 sky130_as_sc_hs__fill_1 FILLER_0_158_541 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_564 ();
 sky130_as_sc_hs__fill_1 FILLER_0_158_568 ();
 sky130_as_sc_hs__fill_1 FILLER_0_158_576 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_582 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_602 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_606 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_610 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_661 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_665 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_674 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_678 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_713 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_717 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_727 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_731 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_735 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_767 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_77 ();
 sky130_as_sc_hs__fill_1 FILLER_0_158_771 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_791 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_803 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_807 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_158_811 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_848 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_852 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_856 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_860 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_864 ();
 sky130_as_sc_hs__fill_8 FILLER_0_158_869 ();
 sky130_as_sc_hs__decap_4 FILLER_0_158_877 ();
 sky130_as_sc_hs__fill_2 FILLER_0_158_881 ();
 sky130_as_sc_hs__decap_3 FILLER_0_158_921 ();
 sky130_as_sc_hs__fill_8 FILLER_0_158_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_158_956 ();
 sky130_as_sc_hs__fill_8 FILLER_0_158_972 ();
 sky130_as_sc_hs__decap_4 FILLER_0_159_105 ();
 sky130_as_sc_hs__fill_8 FILLER_0_159_1051 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_1059 ();
 sky130_as_sc_hs__fill_8 FILLER_0_159_1065 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_1073 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_1079 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_1095 ();
 sky130_as_sc_hs__fill_8 FILLER_0_159_1111 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_1119 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_1137 ();
 sky130_as_sc_hs__fill_8 FILLER_0_159_1145 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_1153 ();
 sky130_as_sc_hs__fill_8 FILLER_0_159_1161 ();
 sky130_as_sc_hs__decap_4 FILLER_0_159_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_159_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_159_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_159_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_159_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_159_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_221 ();
 sky130_as_sc_hs__decap_4 FILLER_0_159_225 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_229 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_249 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_277 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_294 ();
 sky130_as_sc_hs__decap_4 FILLER_0_159_299 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_305 ();
 sky130_as_sc_hs__decap_4 FILLER_0_159_309 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_313 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_316 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_320 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_328 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_332 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_341 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_345 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_393 ();
 sky130_as_sc_hs__decap_4 FILLER_0_159_405 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_409 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_431 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_445 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_478 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_159_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_539 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_556 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_569 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_615 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_628 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_632 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_644 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_648 ();
 sky130_as_sc_hs__decap_4 FILLER_0_159_653 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_659 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_663 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_715 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_725 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_745 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_749 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_774 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_778 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_785 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_821 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_832 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_838 ();
 sky130_as_sc_hs__fill_1 FILLER_0_159_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_850 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_854 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_858 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_862 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_878 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_89 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_894 ();
 sky130_as_sc_hs__decap_3 FILLER_0_159_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_904 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_920 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_936 ();
 sky130_as_sc_hs__fill_8 FILLER_0_159_953 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_961 ();
 sky130_as_sc_hs__fill_2 FILLER_0_159_986 ();
 sky130_as_sc_hs__decap_16 FILLER_0_159_992 ();
 sky130_as_sc_hs__decap_4 FILLER_0_15_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1025 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_103 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_15_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1065 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_107 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1097 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_111 ();
 sky130_as_sc_hs__decap_4 FILLER_0_15_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_15_1169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_117 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_15_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_15_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_15_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_136 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_140 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_144 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_148 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_152 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_156 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_160 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_164 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_15_177 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_181 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_184 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_188 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_192 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_208 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_225 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_241 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_15_273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_285 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_309 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_315 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_321 ();
 sky130_as_sc_hs__fill_8 FILLER_0_15_35 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_372 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_393 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_415 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_423 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_43 ();
 sky130_as_sc_hs__decap_4 FILLER_0_15_431 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_437 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_446 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_453 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_47 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_475 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_492 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_501 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_513 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_517 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_521 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_532 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_536 ();
 sky130_as_sc_hs__decap_4 FILLER_0_15_548 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_55 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_552 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_561 ();
 sky130_as_sc_hs__decap_4 FILLER_0_15_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_573 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_581 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_589 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_599 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_614 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_64 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_669 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_678 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_68 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_711 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_72 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_723 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_727 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_735 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_745 ();
 sky130_as_sc_hs__decap_4 FILLER_0_15_77 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_770 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_781 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_805 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_809 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_820 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_824 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_828 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_832 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_84 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_857 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_861 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_88 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_894 ();
 sky130_as_sc_hs__fill_1 FILLER_0_15_909 ();
 sky130_as_sc_hs__decap_4 FILLER_0_15_92 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_929 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_941 ();
 sky130_as_sc_hs__fill_2 FILLER_0_15_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_969 ();
 sky130_as_sc_hs__decap_3 FILLER_0_15_98 ();
 sky130_as_sc_hs__decap_16 FILLER_0_15_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_101 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_1019 ();
 sky130_as_sc_hs__fill_8 FILLER_0_160_1025 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_1033 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_1041 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_1057 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_1073 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_1114 ();
 sky130_as_sc_hs__decap_4 FILLER_0_160_1130 ();
 sky130_as_sc_hs__fill_1 FILLER_0_160_1139 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_1170 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_1186 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_1202 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_1221 ();
 sky130_as_sc_hs__fill_8 FILLER_0_160_1237 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_1245 ();
 sky130_as_sc_hs__fill_8 FILLER_0_160_1252 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_160_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_160_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_160_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_160_213 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_226 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_230 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_234 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_238 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_242 ();
 sky130_as_sc_hs__fill_1 FILLER_0_160_251 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_258 ();
 sky130_as_sc_hs__fill_1 FILLER_0_160_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_306 ();
 sky130_as_sc_hs__decap_4 FILLER_0_160_309 ();
 sky130_as_sc_hs__decap_4 FILLER_0_160_334 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_340 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_344 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_348 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_352 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_360 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_389 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_418 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_461 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_489 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_493 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_497 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_514 ();
 sky130_as_sc_hs__decap_4 FILLER_0_160_526 ();
 sky130_as_sc_hs__fill_1 FILLER_0_160_546 ();
 sky130_as_sc_hs__fill_1 FILLER_0_160_555 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_575 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_585 ();
 sky130_as_sc_hs__fill_1 FILLER_0_160_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_598 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_61 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_628 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_640 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_649 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_675 ();
 sky130_as_sc_hs__fill_1 FILLER_0_160_679 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_698 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_701 ();
 sky130_as_sc_hs__fill_1 FILLER_0_160_717 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_726 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_742 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_746 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_754 ();
 sky130_as_sc_hs__fill_1 FILLER_0_160_757 ();
 sky130_as_sc_hs__decap_4 FILLER_0_160_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_785 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_813 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_857 ();
 sky130_as_sc_hs__decap_4 FILLER_0_160_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_865 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_869 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_160_906 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_922 ();
 sky130_as_sc_hs__decap_4 FILLER_0_160_944 ();
 sky130_as_sc_hs__fill_2 FILLER_0_160_948 ();
 sky130_as_sc_hs__fill_8 FILLER_0_160_969 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_977 ();
 sky130_as_sc_hs__fill_8 FILLER_0_160_981 ();
 sky130_as_sc_hs__decap_4 FILLER_0_160_989 ();
 sky130_as_sc_hs__decap_3 FILLER_0_160_993 ();
 sky130_as_sc_hs__fill_1 FILLER_0_161_1007 ();
 sky130_as_sc_hs__fill_8 FILLER_0_161_1009 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_1017 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_105 ();
 sky130_as_sc_hs__fill_8 FILLER_0_161_1054 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_113 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_1137 ();
 sky130_as_sc_hs__fill_1 FILLER_0_161_1141 ();
 sky130_as_sc_hs__fill_8 FILLER_0_161_1147 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_1155 ();
 sky130_as_sc_hs__fill_8 FILLER_0_161_1162 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_1170 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_1174 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_1229 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_1233 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_1237 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_1260 ();
 sky130_as_sc_hs__fill_1 FILLER_0_161_1276 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_217 ();
 sky130_as_sc_hs__fill_1 FILLER_0_161_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_229 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_289 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_313 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_319 ();
 sky130_as_sc_hs__fill_1 FILLER_0_161_342 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_362 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_366 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_370 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_374 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_378 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_393 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_403 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_409 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_413 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_438 ();
 sky130_as_sc_hs__fill_1 FILLER_0_161_460 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_513 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_536 ();
 sky130_as_sc_hs__fill_1 FILLER_0_161_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_556 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_561 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_566 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_594 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_613 ();
 sky130_as_sc_hs__fill_1 FILLER_0_161_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_642 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_646 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_656 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_660 ();
 sky130_as_sc_hs__fill_1 FILLER_0_161_678 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_722 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_726 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_777 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_781 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_818 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_822 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_833 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_161_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_853 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_869 ();
 sky130_as_sc_hs__fill_8 FILLER_0_161_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_161_953 ();
 sky130_as_sc_hs__decap_4 FILLER_0_161_969 ();
 sky130_as_sc_hs__decap_3 FILLER_0_161_973 ();
 sky130_as_sc_hs__fill_8 FILLER_0_161_999 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_1001 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_1017 ();
 sky130_as_sc_hs__decap_3 FILLER_0_162_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_1064 ();
 sky130_as_sc_hs__fill_8 FILLER_0_162_1080 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_1088 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_1109 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_1125 ();
 sky130_as_sc_hs__fill_8 FILLER_0_162_1134 ();
 sky130_as_sc_hs__fill_1 FILLER_0_162_1147 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_1154 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_1170 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_1186 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_1202 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_162_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_162_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_162_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_162_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_197 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_217 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_229 ();
 sky130_as_sc_hs__decap_3 FILLER_0_162_266 ();
 sky130_as_sc_hs__fill_1 FILLER_0_162_27 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_285 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_162_307 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_328 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_338 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_371 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_407 ();
 sky130_as_sc_hs__fill_1 FILLER_0_162_414 ();
 sky130_as_sc_hs__fill_1 FILLER_0_162_421 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_459 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_469 ();
 sky130_as_sc_hs__fill_1 FILLER_0_162_473 ();
 sky130_as_sc_hs__fill_1 FILLER_0_162_493 ();
 sky130_as_sc_hs__decap_3 FILLER_0_162_510 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_544 ();
 sky130_as_sc_hs__fill_1 FILLER_0_162_587 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_597 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_601 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_607 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_61 ();
 sky130_as_sc_hs__fill_1 FILLER_0_162_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_634 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_638 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_642 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_664 ();
 sky130_as_sc_hs__fill_1 FILLER_0_162_668 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_679 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_683 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_687 ();
 sky130_as_sc_hs__decap_3 FILLER_0_162_691 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_696 ();
 sky130_as_sc_hs__decap_3 FILLER_0_162_706 ();
 sky130_as_sc_hs__decap_3 FILLER_0_162_722 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_746 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_765 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_769 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_77 ();
 sky130_as_sc_hs__decap_3 FILLER_0_162_773 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_794 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_798 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_802 ();
 sky130_as_sc_hs__decap_3 FILLER_0_162_809 ();
 sky130_as_sc_hs__decap_3 FILLER_0_162_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_162_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_843 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_847 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_85 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_863 ();
 sky130_as_sc_hs__fill_1 FILLER_0_162_867 ();
 sky130_as_sc_hs__fill_8 FILLER_0_162_869 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_877 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_881 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_906 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_922 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_162_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_162_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_162_977 ();
 sky130_as_sc_hs__fill_2 FILLER_0_162_997 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_1036 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_105 ();
 sky130_as_sc_hs__fill_8 FILLER_0_163_1052 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_1060 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_163_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_163_1117 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_1125 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_1159 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_1175 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_163_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_163_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_163_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_19 ();
 sky130_as_sc_hs__fill_8 FILLER_0_163_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_209 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_216 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_220 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_245 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_270 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_315 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_319 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_323 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_332 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_345 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_35 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_372 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_409 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_449 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_466 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_470 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_163_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_513 ();
 sky130_as_sc_hs__decap_3 FILLER_0_163_519 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_524 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_528 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_532 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_536 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_55 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_554 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_590 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_602 ();
 sky130_as_sc_hs__decap_3 FILLER_0_163_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_628 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_648 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_689 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_695 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_73 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_746 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_754 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_758 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_762 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_815 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_819 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_823 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_827 ();
 sky130_as_sc_hs__fill_8 FILLER_0_163_831 ();
 sky130_as_sc_hs__fill_1 FILLER_0_163_839 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_841 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_857 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_873 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_163_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_163_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_163_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_163_949 ();
 sky130_as_sc_hs__fill_8 FILLER_0_163_953 ();
 sky130_as_sc_hs__fill_2 FILLER_0_163_961 ();
 sky130_as_sc_hs__decap_3 FILLER_0_163_986 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_1004 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_1020 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_1037 ();
 sky130_as_sc_hs__decap_3 FILLER_0_164_1041 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_1063 ();
 sky130_as_sc_hs__fill_8 FILLER_0_164_1079 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_1087 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_1091 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_1109 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_1125 ();
 sky130_as_sc_hs__fill_8 FILLER_0_164_1134 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_1142 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_1146 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_164_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_164_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_164_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_164_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_164_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_197 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_213 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_217 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_220 ();
 sky130_as_sc_hs__decap_3 FILLER_0_164_243 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_251 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_269 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_27 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_281 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_285 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_288 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_292 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_296 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_304 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_309 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_313 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_316 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_320 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_329 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_343 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_347 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_350 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_362 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_365 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_369 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_372 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_376 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_380 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_384 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_388 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_410 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_416 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_421 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_494 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_517 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_526 ();
 sky130_as_sc_hs__decap_3 FILLER_0_164_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_555 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_581 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_585 ();
 sky130_as_sc_hs__decap_3 FILLER_0_164_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_602 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_61 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_614 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_631 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_635 ();
 sky130_as_sc_hs__decap_3 FILLER_0_164_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_654 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_698 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_701 ();
 sky130_as_sc_hs__decap_3 FILLER_0_164_705 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_727 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_733 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_754 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_789 ();
 sky130_as_sc_hs__decap_3 FILLER_0_164_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_164_843 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_847 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_85 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_863 ();
 sky130_as_sc_hs__fill_1 FILLER_0_164_867 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_164_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_164_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_164_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_164_977 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_1005 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_1009 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_105 ();
 sky130_as_sc_hs__fill_8 FILLER_0_165_1054 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_1062 ();
 sky130_as_sc_hs__fill_8 FILLER_0_165_1065 ();
 sky130_as_sc_hs__fill_1 FILLER_0_165_1073 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_1117 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_1133 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_1149 ();
 sky130_as_sc_hs__fill_8 FILLER_0_165_1165 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_165_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_201 ();
 sky130_as_sc_hs__fill_1 FILLER_0_165_217 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_220 ();
 sky130_as_sc_hs__fill_1 FILLER_0_165_257 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_266 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_277 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_165_305 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_325 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_345 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_364 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_403 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_407 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_411 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_415 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_419 ();
 sky130_as_sc_hs__fill_1 FILLER_0_165_442 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_461 ();
 sky130_as_sc_hs__fill_1 FILLER_0_165_492 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_498 ();
 sky130_as_sc_hs__fill_1 FILLER_0_165_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_527 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_531 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_539 ();
 sky130_as_sc_hs__fill_1 FILLER_0_165_543 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_546 ();
 sky130_as_sc_hs__fill_1 FILLER_0_165_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_550 ();
 sky130_as_sc_hs__fill_1 FILLER_0_165_559 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_572 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_603 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_625 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_630 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_648 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_660 ();
 sky130_as_sc_hs__fill_1 FILLER_0_165_671 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_689 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_726 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_745 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_765 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_785 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_797 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_816 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_820 ();
 sky130_as_sc_hs__fill_1 FILLER_0_165_824 ();
 sky130_as_sc_hs__fill_2 FILLER_0_165_833 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_837 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_865 ();
 sky130_as_sc_hs__fill_8 FILLER_0_165_881 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_165_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_165_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_165_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_101 ();
 sky130_as_sc_hs__fill_8 FILLER_0_166_1020 ();
 sky130_as_sc_hs__decap_4 FILLER_0_166_1028 ();
 sky130_as_sc_hs__decap_4 FILLER_0_166_1037 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_1041 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_1048 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_1064 ();
 sky130_as_sc_hs__fill_8 FILLER_0_166_1080 ();
 sky130_as_sc_hs__decap_4 FILLER_0_166_1088 ();
 sky130_as_sc_hs__fill_8 FILLER_0_166_1093 ();
 sky130_as_sc_hs__fill_1 FILLER_0_166_1124 ();
 sky130_as_sc_hs__fill_8 FILLER_0_166_1138 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_1146 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_1184 ();
 sky130_as_sc_hs__decap_4 FILLER_0_166_1200 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_166_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_166_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_166_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_166_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_166_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_223 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_227 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_231 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_235 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_243 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_266 ();
 sky130_as_sc_hs__fill_1 FILLER_0_166_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_289 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_304 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_328 ();
 sky130_as_sc_hs__fill_1 FILLER_0_166_346 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_355 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_362 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_416 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_442 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_45 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_467 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_472 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_481 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_490 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_513 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_529 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_541 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_561 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_579 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_584 ();
 sky130_as_sc_hs__fill_1 FILLER_0_166_597 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_61 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_611 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_633 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_650 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_660 ();
 sky130_as_sc_hs__fill_1 FILLER_0_166_679 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_688 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_713 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_717 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_721 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_745 ();
 sky130_as_sc_hs__fill_1 FILLER_0_166_755 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_761 ();
 sky130_as_sc_hs__fill_1 FILLER_0_166_765 ();
 sky130_as_sc_hs__decap_4 FILLER_0_166_77 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_796 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_807 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_166_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_166_853 ();
 sky130_as_sc_hs__fill_8 FILLER_0_166_857 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_865 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_166_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_166_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_166_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_166_981 ();
 sky130_as_sc_hs__decap_4 FILLER_0_166_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_167_1002 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_1006 ();
 sky130_as_sc_hs__fill_8 FILLER_0_167_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_167_1017 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_1021 ();
 sky130_as_sc_hs__fill_1 FILLER_0_167_1042 ();
 sky130_as_sc_hs__decap_4 FILLER_0_167_105 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_1069 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_167_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_1101 ();
 sky130_as_sc_hs__decap_3 FILLER_0_167_1117 ();
 sky130_as_sc_hs__decap_4 FILLER_0_167_1121 ();
 sky130_as_sc_hs__decap_3 FILLER_0_167_1125 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_1133 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_1149 ();
 sky130_as_sc_hs__fill_8 FILLER_0_167_1165 ();
 sky130_as_sc_hs__decap_3 FILLER_0_167_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_167_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_167_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_167_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_167_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_167_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_167_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_19 ();
 sky130_as_sc_hs__fill_8 FILLER_0_167_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_167_209 ();
 sky130_as_sc_hs__fill_1 FILLER_0_167_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_216 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_220 ();
 sky130_as_sc_hs__fill_1 FILLER_0_167_225 ();
 sky130_as_sc_hs__fill_1 FILLER_0_167_245 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_267 ();
 sky130_as_sc_hs__decap_3 FILLER_0_167_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_323 ();
 sky130_as_sc_hs__fill_1 FILLER_0_167_335 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_342 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_35 ();
 sky130_as_sc_hs__decap_4 FILLER_0_167_373 ();
 sky130_as_sc_hs__decap_3 FILLER_0_167_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_413 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_417 ();
 sky130_as_sc_hs__fill_1 FILLER_0_167_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_465 ();
 sky130_as_sc_hs__decap_3 FILLER_0_167_499 ();
 sky130_as_sc_hs__decap_4 FILLER_0_167_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_532 ();
 sky130_as_sc_hs__fill_1 FILLER_0_167_55 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_585 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_594 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_612 ();
 sky130_as_sc_hs__fill_1 FILLER_0_167_633 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_642 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_646 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_706 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_710 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_714 ();
 sky130_as_sc_hs__decap_4 FILLER_0_167_718 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_724 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_741 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_745 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_779 ();
 sky130_as_sc_hs__fill_1 FILLER_0_167_783 ();
 sky130_as_sc_hs__decap_3 FILLER_0_167_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_809 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_813 ();
 sky130_as_sc_hs__fill_1 FILLER_0_167_839 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_865 ();
 sky130_as_sc_hs__fill_8 FILLER_0_167_881 ();
 sky130_as_sc_hs__decap_4 FILLER_0_167_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_167_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_167_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_167_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_167_953 ();
 sky130_as_sc_hs__fill_8 FILLER_0_167_969 ();
 sky130_as_sc_hs__fill_2 FILLER_0_167_977 ();
 sky130_as_sc_hs__fill_1 FILLER_0_168_1001 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_101 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_1025 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_1029 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_1057 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_1073 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_1145 ();
 sky130_as_sc_hs__fill_8 FILLER_0_168_1149 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_1157 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_1161 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_1183 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_1199 ();
 sky130_as_sc_hs__fill_1 FILLER_0_168_1203 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_1257 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_1272 ();
 sky130_as_sc_hs__fill_1 FILLER_0_168_1276 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_168_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_168_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_221 ();
 sky130_as_sc_hs__fill_1 FILLER_0_168_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_306 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_333 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_361 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_370 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_374 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_378 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_398 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_448 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_45 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_495 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_517 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_529 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_538 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_542 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_547 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_586 ();
 sky130_as_sc_hs__fill_1 FILLER_0_168_589 ();
 sky130_as_sc_hs__fill_1 FILLER_0_168_595 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_61 ();
 sky130_as_sc_hs__fill_1 FILLER_0_168_612 ();
 sky130_as_sc_hs__fill_1 FILLER_0_168_632 ();
 sky130_as_sc_hs__fill_1 FILLER_0_168_643 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_653 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_657 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_663 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_667 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_671 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_675 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_679 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_683 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_694 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_698 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_705 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_713 ();
 sky130_as_sc_hs__fill_8 FILLER_0_168_717 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_725 ();
 sky130_as_sc_hs__fill_1 FILLER_0_168_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_754 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_800 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_804 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_808 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_168_821 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_830 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_842 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_846 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_85 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_862 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_866 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_168_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_925 ();
 sky130_as_sc_hs__fill_8 FILLER_0_168_941 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_949 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_974 ();
 sky130_as_sc_hs__fill_2 FILLER_0_168_978 ();
 sky130_as_sc_hs__decap_16 FILLER_0_168_981 ();
 sky130_as_sc_hs__decap_4 FILLER_0_168_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_169_1005 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_1034 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_1038 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_105 ();
 sky130_as_sc_hs__fill_1 FILLER_0_169_1063 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_169_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_169_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_169_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_169_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_1249 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_1265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_1269 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_1275 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_169_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_217 ();
 sky130_as_sc_hs__fill_1 FILLER_0_169_221 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_231 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_235 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_243 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_260 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_264 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_268 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_272 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_276 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_300 ();
 sky130_as_sc_hs__fill_1 FILLER_0_169_304 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_326 ();
 sky130_as_sc_hs__fill_1 FILLER_0_169_335 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_406 ();
 sky130_as_sc_hs__fill_1 FILLER_0_169_428 ();
 sky130_as_sc_hs__decap_3 FILLER_0_169_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_460 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_483 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_498 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_527 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_548 ();
 sky130_as_sc_hs__fill_1 FILLER_0_169_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_552 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_556 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_566 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_570 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_574 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_591 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_683 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_687 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_708 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_712 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_73 ();
 sky130_as_sc_hs__fill_8 FILLER_0_169_733 ();
 sky130_as_sc_hs__fill_1 FILLER_0_169_741 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_744 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_793 ();
 sky130_as_sc_hs__decap_3 FILLER_0_169_797 ();
 sky130_as_sc_hs__fill_1 FILLER_0_169_808 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_817 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_821 ();
 sky130_as_sc_hs__fill_1 FILLER_0_169_825 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_834 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_169_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_853 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_869 ();
 sky130_as_sc_hs__fill_8 FILLER_0_169_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_169_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_169_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_169_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_169_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_1029 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_103 ();
 sky130_as_sc_hs__decap_3 FILLER_0_16_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1069 ();
 sky130_as_sc_hs__decap_3 FILLER_0_16_107 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_16_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1093 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_11 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1109 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_112 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_16_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_116 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_16_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_16_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_15 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_151 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_155 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_159 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_163 ();
 sky130_as_sc_hs__fill_1 FILLER_0_16_167 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_170 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_174 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_178 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_182 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_186 ();
 sky130_as_sc_hs__fill_8 FILLER_0_16_19 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_190 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_194 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_203 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_219 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_235 ();
 sky130_as_sc_hs__fill_1 FILLER_0_16_251 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_253 ();
 sky130_as_sc_hs__fill_8 FILLER_0_16_269 ();
 sky130_as_sc_hs__fill_1 FILLER_0_16_27 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_277 ();
 sky130_as_sc_hs__fill_1 FILLER_0_16_281 ();
 sky130_as_sc_hs__fill_8 FILLER_0_16_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_306 ();
 sky130_as_sc_hs__fill_1 FILLER_0_16_333 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_357 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_384 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_388 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_39 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_392 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_418 ();
 sky130_as_sc_hs__fill_1 FILLER_0_16_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_43 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_438 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_448 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_452 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_464 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_47 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_474 ();
 sky130_as_sc_hs__decap_3 FILLER_0_16_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_488 ();
 sky130_as_sc_hs__decap_3 FILLER_0_16_495 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_500 ();
 sky130_as_sc_hs__fill_1 FILLER_0_16_504 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_51 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_510 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_516 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_520 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_537 ();
 sky130_as_sc_hs__fill_8 FILLER_0_16_541 ();
 sky130_as_sc_hs__decap_3 FILLER_0_16_549 ();
 sky130_as_sc_hs__fill_1 FILLER_0_16_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_560 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_569 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_578 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_58 ();
 sky130_as_sc_hs__fill_1 FILLER_0_16_582 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_611 ();
 sky130_as_sc_hs__fill_1 FILLER_0_16_62 ();
 sky130_as_sc_hs__fill_8 FILLER_0_16_632 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_640 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_65 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_686 ();
 sky130_as_sc_hs__decap_3 FILLER_0_16_69 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_7 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_709 ();
 sky130_as_sc_hs__decap_3 FILLER_0_16_734 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_74 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_757 ();
 sky130_as_sc_hs__fill_1 FILLER_0_16_772 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_78 ();
 sky130_as_sc_hs__fill_1 FILLER_0_16_797 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_82 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_846 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_85 ();
 sky130_as_sc_hs__decap_3 FILLER_0_16_850 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_866 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_873 ();
 sky130_as_sc_hs__decap_3 FILLER_0_16_889 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_89 ();
 sky130_as_sc_hs__fill_1 FILLER_0_16_923 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_942 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_946 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_95 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_950 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_954 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_958 ();
 sky130_as_sc_hs__decap_4 FILLER_0_16_974 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_978 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_981 ();
 sky130_as_sc_hs__fill_2 FILLER_0_16_99 ();
 sky130_as_sc_hs__decap_16 FILLER_0_16_997 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_1014 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_1030 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_1034 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_1149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_1185 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_1257 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_1271 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_1275 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_170_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_213 ();
 sky130_as_sc_hs__fill_1 FILLER_0_170_229 ();
 sky130_as_sc_hs__fill_1 FILLER_0_170_251 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_253 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_263 ();
 sky130_as_sc_hs__fill_1 FILLER_0_170_267 ();
 sky130_as_sc_hs__fill_1 FILLER_0_170_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_302 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_314 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_347 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_352 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_384 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_394 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_417 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_434 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_439 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_467 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_474 ();
 sky130_as_sc_hs__fill_1 FILLER_0_170_485 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_502 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_507 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_519 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_529 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_548 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_557 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_561 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_565 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_589 ();
 sky130_as_sc_hs__fill_1 FILLER_0_170_593 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_620 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_624 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_628 ();
 sky130_as_sc_hs__fill_1 FILLER_0_170_643 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_674 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_689 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_693 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_697 ();
 sky130_as_sc_hs__fill_1 FILLER_0_170_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_712 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_716 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_747 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_751 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_761 ();
 sky130_as_sc_hs__fill_1 FILLER_0_170_765 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_77 ();
 sky130_as_sc_hs__fill_1 FILLER_0_170_776 ();
 sky130_as_sc_hs__fill_1 FILLER_0_170_796 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_810 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_85 ();
 sky130_as_sc_hs__fill_8 FILLER_0_170_853 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_865 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_170_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_170_921 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_948 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_966 ();
 sky130_as_sc_hs__fill_8 FILLER_0_170_970 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_978 ();
 sky130_as_sc_hs__fill_8 FILLER_0_170_981 ();
 sky130_as_sc_hs__decap_4 FILLER_0_170_989 ();
 sky130_as_sc_hs__fill_2 FILLER_0_170_993 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_1005 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_1015 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_1031 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_1047 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_105 ();
 sky130_as_sc_hs__fill_1 FILLER_0_171_1063 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_113 ();
 sky130_as_sc_hs__fill_8 FILLER_0_171_1137 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_1157 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_1233 ();
 sky130_as_sc_hs__fill_8 FILLER_0_171_1249 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_1257 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_1272 ();
 sky130_as_sc_hs__fill_1 FILLER_0_171_1276 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_221 ();
 sky130_as_sc_hs__fill_8 FILLER_0_171_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_252 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_275 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_285 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_324 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_333 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_357 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_361 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_374 ();
 sky130_as_sc_hs__fill_1 FILLER_0_171_391 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_397 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_401 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_405 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_409 ();
 sky130_as_sc_hs__fill_1 FILLER_0_171_421 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_441 ();
 sky130_as_sc_hs__fill_1 FILLER_0_171_445 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_468 ();
 sky130_as_sc_hs__fill_1 FILLER_0_171_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_171_55 ();
 sky130_as_sc_hs__fill_1 FILLER_0_171_559 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_561 ();
 sky130_as_sc_hs__fill_1 FILLER_0_171_565 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_568 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_57 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_604 ();
 sky130_as_sc_hs__fill_1 FILLER_0_171_608 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_622 ();
 sky130_as_sc_hs__fill_1 FILLER_0_171_644 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_655 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_659 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_663 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_667 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_683 ();
 sky130_as_sc_hs__fill_1 FILLER_0_171_704 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_713 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_717 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_721 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_754 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_775 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_779 ();
 sky130_as_sc_hs__fill_1 FILLER_0_171_783 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_815 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_819 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_823 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_834 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_171_848 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_852 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_868 ();
 sky130_as_sc_hs__fill_8 FILLER_0_171_884 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_89 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_892 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_171_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_171_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_171_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_101 ();
 sky130_as_sc_hs__decap_4 FILLER_0_172_1013 ();
 sky130_as_sc_hs__fill_8 FILLER_0_172_1064 ();
 sky130_as_sc_hs__decap_4 FILLER_0_172_1072 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_1097 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_1113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_1129 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_172_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_172_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_172_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_137 ();
 sky130_as_sc_hs__fill_8 FILLER_0_172_14 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_172_189 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_213 ();
 sky130_as_sc_hs__decap_4 FILLER_0_172_22 ();
 sky130_as_sc_hs__fill_1 FILLER_0_172_229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_232 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_236 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_240 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_248 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_26 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_266 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_289 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_29 ();
 sky130_as_sc_hs__decap_4 FILLER_0_172_297 ();
 sky130_as_sc_hs__fill_1 FILLER_0_172_301 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_304 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_326 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_352 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_365 ();
 sky130_as_sc_hs__fill_1 FILLER_0_172_383 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_405 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_415 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_429 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_444 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_448 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_452 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_456 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_460 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_474 ();
 sky130_as_sc_hs__fill_1 FILLER_0_172_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_488 ();
 sky130_as_sc_hs__fill_1 FILLER_0_172_503 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_512 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_533 ();
 sky130_as_sc_hs__decap_4 FILLER_0_172_575 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_581 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_602 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_634 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_638 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_642 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_674 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_684 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_688 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_692 ();
 sky130_as_sc_hs__fill_1 FILLER_0_172_701 ();
 sky130_as_sc_hs__fill_1 FILLER_0_172_742 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_751 ();
 sky130_as_sc_hs__fill_1 FILLER_0_172_755 ();
 sky130_as_sc_hs__decap_4 FILLER_0_172_77 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_781 ();
 sky130_as_sc_hs__fill_1 FILLER_0_172_803 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_834 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_85 ();
 sky130_as_sc_hs__fill_8 FILLER_0_172_854 ();
 sky130_as_sc_hs__decap_4 FILLER_0_172_862 ();
 sky130_as_sc_hs__fill_2 FILLER_0_172_866 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_172_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_172_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_172_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_172_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_1028 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_1044 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_1060 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_1065 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_109 ();
 sky130_as_sc_hs__fill_8 FILLER_0_173_1106 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_1114 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_1118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_1177 ();
 sky130_as_sc_hs__fill_1 FILLER_0_173_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_1202 ();
 sky130_as_sc_hs__fill_8 FILLER_0_173_1218 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_1226 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_1230 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_173_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_221 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_250 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_266 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_272 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_276 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_287 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_291 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_314 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_330 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_345 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_388 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_422 ();
 sky130_as_sc_hs__fill_1 FILLER_0_173_447 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_454 ();
 sky130_as_sc_hs__fill_1 FILLER_0_173_458 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_461 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_484 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_505 ();
 sky130_as_sc_hs__fill_1 FILLER_0_173_509 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_512 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_534 ();
 sky130_as_sc_hs__fill_1 FILLER_0_173_538 ();
 sky130_as_sc_hs__fill_1 FILLER_0_173_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_57 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_584 ();
 sky130_as_sc_hs__fill_1 FILLER_0_173_588 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_599 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_609 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_614 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_636 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_659 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_697 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_73 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_773 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_797 ();
 sky130_as_sc_hs__fill_2 FILLER_0_173_812 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_865 ();
 sky130_as_sc_hs__fill_8 FILLER_0_173_881 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_173_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_173_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_173_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_101 ();
 sky130_as_sc_hs__decap_4 FILLER_0_174_1013 ();
 sky130_as_sc_hs__fill_1 FILLER_0_174_1017 ();
 sky130_as_sc_hs__fill_8 FILLER_0_174_1022 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_1030 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_1057 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_1073 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_174_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_174_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_174_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_174_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_174_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_174_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_229 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_266 ();
 sky130_as_sc_hs__fill_1 FILLER_0_174_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_288 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_29 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_295 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_304 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_319 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_328 ();
 sky130_as_sc_hs__decap_4 FILLER_0_174_348 ();
 sky130_as_sc_hs__fill_1 FILLER_0_174_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_390 ();
 sky130_as_sc_hs__decap_4 FILLER_0_174_402 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_416 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_440 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_463 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_467 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_496 ();
 sky130_as_sc_hs__fill_1 FILLER_0_174_506 ();
 sky130_as_sc_hs__fill_1 FILLER_0_174_541 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_552 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_569 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_61 ();
 sky130_as_sc_hs__fill_1 FILLER_0_174_624 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_638 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_642 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_661 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_671 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_698 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_713 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_753 ();
 sky130_as_sc_hs__decap_4 FILLER_0_174_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_789 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_793 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_813 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_817 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_843 ();
 sky130_as_sc_hs__fill_2 FILLER_0_174_847 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_85 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_851 ();
 sky130_as_sc_hs__fill_1 FILLER_0_174_867 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_174_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_174_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_174_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_174_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_175_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_1047 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_105 ();
 sky130_as_sc_hs__fill_1 FILLER_0_175_1063 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_175_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_175_1117 ();
 sky130_as_sc_hs__fill_1 FILLER_0_175_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_1141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_1157 ();
 sky130_as_sc_hs__decap_3 FILLER_0_175_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_175_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_175_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_175_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_217 ();
 sky130_as_sc_hs__fill_1 FILLER_0_175_221 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_231 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_235 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_243 ();
 sky130_as_sc_hs__decap_3 FILLER_0_175_252 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_268 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_272 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_276 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_305 ();
 sky130_as_sc_hs__fill_1 FILLER_0_175_309 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_35 ();
 sky130_as_sc_hs__fill_1 FILLER_0_175_350 ();
 sky130_as_sc_hs__decap_3 FILLER_0_175_389 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_420 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_424 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_428 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_432 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_436 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_440 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_444 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_455 ();
 sky130_as_sc_hs__fill_1 FILLER_0_175_483 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_497 ();
 sky130_as_sc_hs__fill_1 FILLER_0_175_501 ();
 sky130_as_sc_hs__fill_1 FILLER_0_175_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_525 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_535 ();
 sky130_as_sc_hs__fill_1 FILLER_0_175_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_57 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_576 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_614 ();
 sky130_as_sc_hs__decap_3 FILLER_0_175_617 ();
 sky130_as_sc_hs__decap_3 FILLER_0_175_641 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_668 ();
 sky130_as_sc_hs__fill_1 FILLER_0_175_683 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_689 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_693 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_719 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_723 ();
 sky130_as_sc_hs__fill_1 FILLER_0_175_727 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_755 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_759 ();
 sky130_as_sc_hs__decap_3 FILLER_0_175_763 ();
 sky130_as_sc_hs__fill_1 FILLER_0_175_774 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_780 ();
 sky130_as_sc_hs__fill_1 FILLER_0_175_785 ();
 sky130_as_sc_hs__decap_3 FILLER_0_175_794 ();
 sky130_as_sc_hs__fill_2 FILLER_0_175_852 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_856 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_872 ();
 sky130_as_sc_hs__fill_8 FILLER_0_175_888 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_89 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_175_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_175_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_175_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_176_1033 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_1037 ();
 sky130_as_sc_hs__fill_1 FILLER_0_176_1064 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_1088 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_176_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_176_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_176_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_176_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_176_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_176_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_197 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_217 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_258 ();
 sky130_as_sc_hs__fill_1 FILLER_0_176_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_309 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_358 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_418 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_426 ();
 sky130_as_sc_hs__fill_1 FILLER_0_176_430 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_433 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_474 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_500 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_520 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_528 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_539 ();
 sky130_as_sc_hs__decap_3 FILLER_0_176_562 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_581 ();
 sky130_as_sc_hs__fill_1 FILLER_0_176_585 ();
 sky130_as_sc_hs__fill_1 FILLER_0_176_589 ();
 sky130_as_sc_hs__fill_1 FILLER_0_176_595 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_61 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_612 ();
 sky130_as_sc_hs__fill_1 FILLER_0_176_616 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_635 ();
 sky130_as_sc_hs__decap_3 FILLER_0_176_639 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_677 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_719 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_723 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_727 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_731 ();
 sky130_as_sc_hs__decap_3 FILLER_0_176_757 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_77 ();
 sky130_as_sc_hs__fill_1 FILLER_0_176_779 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_803 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_807 ();
 sky130_as_sc_hs__decap_3 FILLER_0_176_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_176_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_176_830 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_85 ();
 sky130_as_sc_hs__fill_8 FILLER_0_176_856 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_864 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_176_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_176_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_176_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_176_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_177_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_177_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_177_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_177_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_177_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_177_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_177_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_177_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_201 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_217 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_220 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_245 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_263 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_281 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_299 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_305 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_313 ();
 sky130_as_sc_hs__decap_3 FILLER_0_177_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_35 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_375 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_420 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_440 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_446 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_473 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_513 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_527 ();
 sky130_as_sc_hs__decap_3 FILLER_0_177_539 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_549 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_55 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_553 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_556 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_576 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_584 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_601 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_607 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_611 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_615 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_621 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_634 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_638 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_642 ();
 sky130_as_sc_hs__decap_3 FILLER_0_177_646 ();
 sky130_as_sc_hs__decap_3 FILLER_0_177_651 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_656 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_660 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_681 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_714 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_718 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_721 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_725 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_73 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_751 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_776 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_797 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_801 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_805 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_809 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_819 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_823 ();
 sky130_as_sc_hs__fill_2 FILLER_0_177_835 ();
 sky130_as_sc_hs__fill_1 FILLER_0_177_839 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_865 ();
 sky130_as_sc_hs__fill_8 FILLER_0_177_881 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_177_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_177_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_177_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_177_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_178_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_1037 ();
 sky130_as_sc_hs__fill_8 FILLER_0_178_1053 ();
 sky130_as_sc_hs__decap_4 FILLER_0_178_1061 ();
 sky130_as_sc_hs__fill_1 FILLER_0_178_1065 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_178_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_178_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_178_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_178_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_178_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_178_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_197 ();
 sky130_as_sc_hs__decap_4 FILLER_0_178_213 ();
 sky130_as_sc_hs__fill_1 FILLER_0_178_217 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_220 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_224 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_228 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_232 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_236 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_240 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_264 ();
 sky130_as_sc_hs__fill_1 FILLER_0_178_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_292 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_178_307 ();
 sky130_as_sc_hs__decap_4 FILLER_0_178_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_315 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_319 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_350 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_361 ();
 sky130_as_sc_hs__fill_1 FILLER_0_178_365 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_392 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_397 ();
 sky130_as_sc_hs__fill_1 FILLER_0_178_419 ();
 sky130_as_sc_hs__fill_1 FILLER_0_178_421 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_45 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_457 ();
 sky130_as_sc_hs__fill_1 FILLER_0_178_496 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_508 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_529 ();
 sky130_as_sc_hs__fill_1 FILLER_0_178_541 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_566 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_589 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_612 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_637 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_680 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_690 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_694 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_698 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_705 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_709 ();
 sky130_as_sc_hs__fill_1 FILLER_0_178_713 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_752 ();
 sky130_as_sc_hs__decap_4 FILLER_0_178_77 ();
 sky130_as_sc_hs__fill_1 FILLER_0_178_773 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_178_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_819 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_823 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_834 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_838 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_842 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_85 ();
 sky130_as_sc_hs__fill_8 FILLER_0_178_858 ();
 sky130_as_sc_hs__fill_2 FILLER_0_178_866 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_178_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_178_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_178_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_178_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_179_1005 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_1009 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_1013 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_1038 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_105 ();
 sky130_as_sc_hs__fill_8 FILLER_0_179_1054 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_1084 ();
 sky130_as_sc_hs__decap_3 FILLER_0_179_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_1100 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_1116 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_179_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_179_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_179_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_179_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_217 ();
 sky130_as_sc_hs__fill_1 FILLER_0_179_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_254 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_272 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_304 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_308 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_312 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_316 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_320 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_328 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_332 ();
 sky130_as_sc_hs__decap_3 FILLER_0_179_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_35 ();
 sky130_as_sc_hs__fill_1 FILLER_0_179_353 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_359 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_385 ();
 sky130_as_sc_hs__fill_1 FILLER_0_179_389 ();
 sky130_as_sc_hs__decap_3 FILLER_0_179_412 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_434 ();
 sky130_as_sc_hs__fill_1 FILLER_0_179_438 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_446 ();
 sky130_as_sc_hs__decap_3 FILLER_0_179_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_460 ();
 sky130_as_sc_hs__decap_3 FILLER_0_179_483 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_491 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_500 ();
 sky130_as_sc_hs__fill_1 FILLER_0_179_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_179_530 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_539 ();
 sky130_as_sc_hs__fill_1 FILLER_0_179_55 ();
 sky130_as_sc_hs__fill_1 FILLER_0_179_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_570 ();
 sky130_as_sc_hs__fill_1 FILLER_0_179_591 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_608 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_612 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_649 ();
 sky130_as_sc_hs__decap_3 FILLER_0_179_669 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_689 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_726 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_752 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_756 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_789 ();
 sky130_as_sc_hs__decap_3 FILLER_0_179_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_815 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_833 ();
 sky130_as_sc_hs__decap_3 FILLER_0_179_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_846 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_850 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_866 ();
 sky130_as_sc_hs__fill_8 FILLER_0_179_882 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_89 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_890 ();
 sky130_as_sc_hs__fill_2 FILLER_0_179_894 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_179_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_179_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_179_985 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1009 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1081 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1097 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_11 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1121 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_1169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_117 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1193 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_120 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_1249 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_125 ();
 sky130_as_sc_hs__fill_8 FILLER_0_17_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_14 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_150 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_156 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_167 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_173 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_176 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_18 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_181 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_185 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_193 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_202 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_206 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_210 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_214 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_218 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_22 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_223 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_225 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_241 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_257 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_26 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_30 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_335 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_34 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_372 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_376 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_38 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_391 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_417 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_42 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_424 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_432 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_436 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_445 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_48 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_483 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_502 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_52 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_532 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_541 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_550 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_561 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_588 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_607 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_65 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_652 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_68 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_691 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_709 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_74 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_753 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_783 ();
 sky130_as_sc_hs__decap_4 FILLER_0_17_79 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_794 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_800 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_807 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_817 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_851 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_89 ();
 sky130_as_sc_hs__fill_1 FILLER_0_17_895 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_905 ();
 sky130_as_sc_hs__decap_3 FILLER_0_17_909 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_93 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_932 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_936 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_940 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_944 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_948 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_969 ();
 sky130_as_sc_hs__fill_2 FILLER_0_17_97 ();
 sky130_as_sc_hs__decap_16 FILLER_0_17_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_1053 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_1069 ();
 sky130_as_sc_hs__fill_1 FILLER_0_180_1073 ();
 sky130_as_sc_hs__fill_8 FILLER_0_180_1078 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_1086 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_1090 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_180_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_180_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_223 ();
 sky130_as_sc_hs__fill_1 FILLER_0_180_246 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_266 ();
 sky130_as_sc_hs__fill_1 FILLER_0_180_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_304 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_328 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_334 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_343 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_348 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_360 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_371 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_402 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_417 ();
 sky130_as_sc_hs__fill_1 FILLER_0_180_440 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_180_457 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_466 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_472 ();
 sky130_as_sc_hs__fill_1 FILLER_0_180_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_499 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_517 ();
 sky130_as_sc_hs__fill_1 FILLER_0_180_541 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_582 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_586 ();
 sky130_as_sc_hs__fill_1 FILLER_0_180_597 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_603 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_607 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_629 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_641 ();
 sky130_as_sc_hs__fill_1 FILLER_0_180_680 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_697 ();
 sky130_as_sc_hs__fill_1 FILLER_0_180_717 ();
 sky130_as_sc_hs__fill_1 FILLER_0_180_742 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_77 ();
 sky130_as_sc_hs__fill_1 FILLER_0_180_783 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_808 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_81 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_180_848 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_85 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_852 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_180_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_180_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_180_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_1009 ();
 sky130_as_sc_hs__fill_8 FILLER_0_181_1025 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_1033 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_1037 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_1059 ();
 sky130_as_sc_hs__fill_1 FILLER_0_181_1063 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_181_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_217 ();
 sky130_as_sc_hs__fill_1 FILLER_0_181_221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_230 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_234 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_238 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_265 ();
 sky130_as_sc_hs__fill_1 FILLER_0_181_269 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_272 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_276 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_290 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_331 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_388 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_404 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_419 ();
 sky130_as_sc_hs__fill_1 FILLER_0_181_441 ();
 sky130_as_sc_hs__fill_1 FILLER_0_181_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_449 ();
 sky130_as_sc_hs__fill_1 FILLER_0_181_464 ();
 sky130_as_sc_hs__fill_1 FILLER_0_181_503 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_524 ();
 sky130_as_sc_hs__fill_1 FILLER_0_181_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_574 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_597 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_608 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_612 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_630 ();
 sky130_as_sc_hs__fill_1 FILLER_0_181_634 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_643 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_647 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_651 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_655 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_664 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_668 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_673 ();
 sky130_as_sc_hs__fill_1 FILLER_0_181_677 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_686 ();
 sky130_as_sc_hs__fill_1 FILLER_0_181_722 ();
 sky130_as_sc_hs__fill_1 FILLER_0_181_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_814 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_181_845 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_865 ();
 sky130_as_sc_hs__fill_8 FILLER_0_181_881 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_181_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_181_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_181_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_101 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_1013 ();
 sky130_as_sc_hs__fill_1 FILLER_0_182_1037 ();
 sky130_as_sc_hs__fill_8 FILLER_0_182_1042 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_1050 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_1054 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_1060 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_1076 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_182_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_197 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_213 ();
 sky130_as_sc_hs__fill_1 FILLER_0_182_217 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_239 ();
 sky130_as_sc_hs__fill_1 FILLER_0_182_251 ();
 sky130_as_sc_hs__fill_1 FILLER_0_182_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_296 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_353 ();
 sky130_as_sc_hs__fill_1 FILLER_0_182_370 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_409 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_432 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_436 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_45 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_461 ();
 sky130_as_sc_hs__fill_1 FILLER_0_182_465 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_468 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_472 ();
 sky130_as_sc_hs__fill_1 FILLER_0_182_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_502 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_544 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_577 ();
 sky130_as_sc_hs__fill_1 FILLER_0_182_581 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_584 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_589 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_629 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_641 ();
 sky130_as_sc_hs__fill_1 FILLER_0_182_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_654 ();
 sky130_as_sc_hs__fill_1 FILLER_0_182_658 ();
 sky130_as_sc_hs__fill_1 FILLER_0_182_678 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_757 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_761 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_772 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_182_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_833 ();
 sky130_as_sc_hs__fill_2 FILLER_0_182_837 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_841 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_85 ();
 sky130_as_sc_hs__fill_8 FILLER_0_182_857 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_865 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_182_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_182_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_182_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_183_1005 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_1029 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_1045 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_105 ();
 sky130_as_sc_hs__decap_3 FILLER_0_183_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_183_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_183_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_183_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_183_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_183_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_183_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_217 ();
 sky130_as_sc_hs__fill_1 FILLER_0_183_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_272 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_276 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_316 ();
 sky130_as_sc_hs__decap_3 FILLER_0_183_333 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_343 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_35 ();
 sky130_as_sc_hs__fill_1 FILLER_0_183_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_434 ();
 sky130_as_sc_hs__fill_1 FILLER_0_183_449 ();
 sky130_as_sc_hs__fill_1 FILLER_0_183_458 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_467 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_502 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_511 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_534 ();
 sky130_as_sc_hs__fill_1 FILLER_0_183_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_183_576 ();
 sky130_as_sc_hs__fill_1 FILLER_0_183_598 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_612 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_627 ();
 sky130_as_sc_hs__decap_3 FILLER_0_183_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_664 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_668 ();
 sky130_as_sc_hs__fill_1 FILLER_0_183_692 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_712 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_716 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_720 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_724 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_754 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_758 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_762 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_772 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_776 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_812 ();
 sky130_as_sc_hs__fill_2 FILLER_0_183_833 ();
 sky130_as_sc_hs__decap_3 FILLER_0_183_837 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_841 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_857 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_873 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_183_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_183_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_183_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_183_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1016 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_1032 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_184_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_197 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_213 ();
 sky130_as_sc_hs__fill_1 FILLER_0_184_217 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_220 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_224 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_228 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_232 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_236 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_250 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_184_265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_268 ();
 sky130_as_sc_hs__fill_1 FILLER_0_184_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_272 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_280 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_284 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_288 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_184_320 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_329 ();
 sky130_as_sc_hs__fill_1 FILLER_0_184_333 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_344 ();
 sky130_as_sc_hs__fill_1 FILLER_0_184_363 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_373 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_388 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_397 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_401 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_405 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_417 ();
 sky130_as_sc_hs__fill_1 FILLER_0_184_421 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_45 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_457 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_496 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_516 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_520 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_544 ();
 sky130_as_sc_hs__fill_1 FILLER_0_184_566 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_584 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_603 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_625 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_629 ();
 sky130_as_sc_hs__fill_1 FILLER_0_184_633 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_636 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_640 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_645 ();
 sky130_as_sc_hs__fill_1 FILLER_0_184_655 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_664 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_668 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_674 ();
 sky130_as_sc_hs__fill_1 FILLER_0_184_678 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_698 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_705 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_733 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_757 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_786 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_790 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_807 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_184_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_184_840 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_844 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_85 ();
 sky130_as_sc_hs__fill_8 FILLER_0_184_860 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_184_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_184_925 ();
 sky130_as_sc_hs__fill_8 FILLER_0_184_941 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_949 ();
 sky130_as_sc_hs__fill_8 FILLER_0_184_972 ();
 sky130_as_sc_hs__fill_8 FILLER_0_184_981 ();
 sky130_as_sc_hs__decap_4 FILLER_0_184_989 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_185_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_201 ();
 sky130_as_sc_hs__fill_1 FILLER_0_185_217 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_220 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_244 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_256 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_277 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_290 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_294 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_185_314 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_331 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_35 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_356 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_367 ();
 sky130_as_sc_hs__fill_1 FILLER_0_185_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_407 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_417 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_423 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_446 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_457 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_461 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_465 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_474 ();
 sky130_as_sc_hs__fill_1 FILLER_0_185_478 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_481 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_485 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_489 ();
 sky130_as_sc_hs__fill_1 FILLER_0_185_503 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_51 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_510 ();
 sky130_as_sc_hs__fill_1 FILLER_0_185_514 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_549 ();
 sky130_as_sc_hs__fill_1 FILLER_0_185_55 ();
 sky130_as_sc_hs__fill_1 FILLER_0_185_553 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_556 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_576 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_580 ();
 sky130_as_sc_hs__fill_1 FILLER_0_185_584 ();
 sky130_as_sc_hs__fill_1 FILLER_0_185_604 ();
 sky130_as_sc_hs__fill_1 FILLER_0_185_610 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_630 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_634 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_638 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_642 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_647 ();
 sky130_as_sc_hs__fill_1 FILLER_0_185_651 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_670 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_673 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_695 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_717 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_73 ();
 sky130_as_sc_hs__fill_1 FILLER_0_185_742 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_772 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_776 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_804 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_808 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_812 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_816 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_820 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_834 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_185_845 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_865 ();
 sky130_as_sc_hs__fill_8 FILLER_0_185_881 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_185_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_185_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_185_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_186_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_186_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_186_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_186_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_1109 ();
 sky130_as_sc_hs__decap_4 FILLER_0_186_1144 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_186_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_186_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_186_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_186_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_186_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_186_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_186_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_186_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_186_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_186_213 ();
 sky130_as_sc_hs__fill_1 FILLER_0_186_221 ();
 sky130_as_sc_hs__fill_1 FILLER_0_186_241 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_250 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_258 ();
 sky130_as_sc_hs__fill_1 FILLER_0_186_27 ();
 sky130_as_sc_hs__decap_4 FILLER_0_186_283 ();
 sky130_as_sc_hs__fill_1 FILLER_0_186_287 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_290 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_186_307 ();
 sky130_as_sc_hs__decap_3 FILLER_0_186_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_326 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_330 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_334 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_338 ();
 sky130_as_sc_hs__fill_1 FILLER_0_186_363 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_418 ();
 sky130_as_sc_hs__decap_3 FILLER_0_186_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_430 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_434 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_438 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_442 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_186_451 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_525 ();
 sky130_as_sc_hs__fill_1 FILLER_0_186_533 ();
 sky130_as_sc_hs__fill_1 FILLER_0_186_539 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_559 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_563 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_586 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_589 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_654 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_658 ();
 sky130_as_sc_hs__fill_1 FILLER_0_186_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_751 ();
 sky130_as_sc_hs__fill_1 FILLER_0_186_755 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_757 ();
 sky130_as_sc_hs__decap_4 FILLER_0_186_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_771 ();
 sky130_as_sc_hs__decap_3 FILLER_0_186_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_810 ();
 sky130_as_sc_hs__decap_3 FILLER_0_186_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_843 ();
 sky130_as_sc_hs__fill_2 FILLER_0_186_847 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_85 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_851 ();
 sky130_as_sc_hs__fill_1 FILLER_0_186_867 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_186_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_186_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_186_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_186_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_186_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_187_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_217 ();
 sky130_as_sc_hs__fill_1 FILLER_0_187_221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_276 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_313 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_334 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_35 ();
 sky130_as_sc_hs__fill_1 FILLER_0_187_356 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_373 ();
 sky130_as_sc_hs__fill_1 FILLER_0_187_377 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_385 ();
 sky130_as_sc_hs__fill_1 FILLER_0_187_389 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_393 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_403 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_414 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_418 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_446 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_470 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_493 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_187_524 ();
 sky130_as_sc_hs__fill_1 FILLER_0_187_546 ();
 sky130_as_sc_hs__fill_1 FILLER_0_187_55 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_569 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_580 ();
 sky130_as_sc_hs__fill_1 FILLER_0_187_601 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_610 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_614 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_621 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_625 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_636 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_662 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_666 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_682 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_686 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_703 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_707 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_711 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_718 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_722 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_726 ();
 sky130_as_sc_hs__fill_1 FILLER_0_187_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_743 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_789 ();
 sky130_as_sc_hs__fill_1 FILLER_0_187_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_802 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_806 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_846 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_850 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_854 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_870 ();
 sky130_as_sc_hs__fill_8 FILLER_0_187_886 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_89 ();
 sky130_as_sc_hs__fill_2 FILLER_0_187_894 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_187_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_187_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_187_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_188_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_188_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_188_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_188_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_188_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_188_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_188_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_188_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_188_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_188_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_188_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_188_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_188_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_188_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_188_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_188_213 ();
 sky130_as_sc_hs__fill_1 FILLER_0_188_27 ();
 sky130_as_sc_hs__decap_4 FILLER_0_188_282 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_288 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_188_305 ();
 sky130_as_sc_hs__decap_4 FILLER_0_188_341 ();
 sky130_as_sc_hs__fill_1 FILLER_0_188_352 ();
 sky130_as_sc_hs__fill_1 FILLER_0_188_363 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_384 ();
 sky130_as_sc_hs__decap_3 FILLER_0_188_394 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_399 ();
 sky130_as_sc_hs__fill_1 FILLER_0_188_419 ();
 sky130_as_sc_hs__fill_1 FILLER_0_188_440 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_45 ();
 sky130_as_sc_hs__decap_4 FILLER_0_188_454 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_460 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_464 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_485 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_489 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_512 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_549 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_559 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_584 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_597 ();
 sky130_as_sc_hs__decap_3 FILLER_0_188_609 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_61 ();
 sky130_as_sc_hs__fill_1 FILLER_0_188_622 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_642 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_698 ();
 sky130_as_sc_hs__fill_1 FILLER_0_188_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_715 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_725 ();
 sky130_as_sc_hs__fill_1 FILLER_0_188_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_754 ();
 sky130_as_sc_hs__decap_4 FILLER_0_188_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_781 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_798 ();
 sky130_as_sc_hs__decap_3 FILLER_0_188_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_817 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_821 ();
 sky130_as_sc_hs__fill_1 FILLER_0_188_825 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_842 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_846 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_850 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_854 ();
 sky130_as_sc_hs__fill_8 FILLER_0_188_858 ();
 sky130_as_sc_hs__fill_2 FILLER_0_188_866 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_188_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_188_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_188_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_188_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_188_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_113 ();
 sky130_as_sc_hs__fill_8 FILLER_0_189_1137 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_1145 ();
 sky130_as_sc_hs__fill_8 FILLER_0_189_1166 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_1174 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_189_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_221 ();
 sky130_as_sc_hs__fill_1 FILLER_0_189_244 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_264 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_268 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_272 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_276 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_300 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_333 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_341 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_35 ();
 sky130_as_sc_hs__fill_1 FILLER_0_189_363 ();
 sky130_as_sc_hs__fill_1 FILLER_0_189_383 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_406 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_410 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_414 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_426 ();
 sky130_as_sc_hs__fill_1 FILLER_0_189_430 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_446 ();
 sky130_as_sc_hs__fill_1 FILLER_0_189_457 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_490 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_495 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_51 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_547 ();
 sky130_as_sc_hs__fill_1 FILLER_0_189_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_558 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_189_579 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_588 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_613 ();
 sky130_as_sc_hs__fill_1 FILLER_0_189_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_189_671 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_684 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_688 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_692 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_726 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_73 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_737 ();
 sky130_as_sc_hs__fill_1 FILLER_0_189_756 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_778 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_812 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_816 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_820 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_830 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_189_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_853 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_869 ();
 sky130_as_sc_hs__fill_8 FILLER_0_189_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_189_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_189_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_189_985 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_10 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_1029 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_103 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1069 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_107 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1205 ();
 sky130_as_sc_hs__fill_1 FILLER_0_18_121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_127 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_133 ();
 sky130_as_sc_hs__fill_1 FILLER_0_18_137 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_14 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_147 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_151 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_184 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_20 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_207 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_211 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_215 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_219 ();
 sky130_as_sc_hs__fill_1 FILLER_0_18_223 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_226 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_230 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_234 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_238 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_24 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_242 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_247 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_253 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_306 ();
 sky130_as_sc_hs__fill_1 FILLER_0_18_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_315 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_33 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_346 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_361 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_365 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_369 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_37 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_41 ();
 sky130_as_sc_hs__fill_1 FILLER_0_18_414 ();
 sky130_as_sc_hs__fill_1 FILLER_0_18_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_430 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_455 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_46 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_496 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_50 ();
 sky130_as_sc_hs__fill_1 FILLER_0_18_513 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_54 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_568 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_58 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_599 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_612 ();
 sky130_as_sc_hs__fill_1 FILLER_0_18_616 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_63 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_630 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_655 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_67 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_676 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_697 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_71 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_711 ();
 sky130_as_sc_hs__fill_1 FILLER_0_18_728 ();
 sky130_as_sc_hs__fill_1 FILLER_0_18_746 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_76 ();
 sky130_as_sc_hs__fill_1 FILLER_0_18_777 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_80 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_809 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_823 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_827 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_831 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_835 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_847 ();
 sky130_as_sc_hs__decap_4 FILLER_0_18_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_851 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_865 ();
 sky130_as_sc_hs__fill_1 FILLER_0_18_874 ();
 sky130_as_sc_hs__fill_1 FILLER_0_18_884 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_91 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_914 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_922 ();
 sky130_as_sc_hs__decap_3 FILLER_0_18_943 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_95 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_958 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_962 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_978 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_981 ();
 sky130_as_sc_hs__fill_2 FILLER_0_18_99 ();
 sky130_as_sc_hs__decap_16 FILLER_0_18_997 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_190_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_190_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_190_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_190_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_190_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_190_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_190_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_190_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_213 ();
 sky130_as_sc_hs__fill_8 FILLER_0_190_229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_248 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_257 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_190_27 ();
 sky130_as_sc_hs__decap_4 FILLER_0_190_278 ();
 sky130_as_sc_hs__fill_1 FILLER_0_190_282 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_285 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_318 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_346 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_365 ();
 sky130_as_sc_hs__fill_1 FILLER_0_190_384 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_417 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_437 ();
 sky130_as_sc_hs__decap_4 FILLER_0_190_447 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_453 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_492 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_513 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_528 ();
 sky130_as_sc_hs__fill_1 FILLER_0_190_533 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_577 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_597 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_61 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_631 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_685 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_695 ();
 sky130_as_sc_hs__fill_1 FILLER_0_190_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_705 ();
 sky130_as_sc_hs__fill_1 FILLER_0_190_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_734 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_752 ();
 sky130_as_sc_hs__decap_4 FILLER_0_190_77 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_776 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_803 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_807 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_190_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_190_826 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_85 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_852 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_190_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_190_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_190_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_190_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_113 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_1158 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_1174 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_191_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_221 ();
 sky130_as_sc_hs__fill_8 FILLER_0_191_225 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_233 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_237 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_277 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_318 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_328 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_332 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_379 ();
 sky130_as_sc_hs__fill_1 FILLER_0_191_391 ();
 sky130_as_sc_hs__fill_1 FILLER_0_191_409 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_420 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_435 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_440 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_444 ();
 sky130_as_sc_hs__fill_1 FILLER_0_191_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_474 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_489 ();
 sky130_as_sc_hs__fill_1 FILLER_0_191_493 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_191_539 ();
 sky130_as_sc_hs__fill_1 FILLER_0_191_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_556 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_587 ();
 sky130_as_sc_hs__fill_1 FILLER_0_191_597 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_614 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_629 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_637 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_666 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_726 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_793 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_797 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_824 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_828 ();
 sky130_as_sc_hs__fill_2 FILLER_0_191_836 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_841 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_857 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_873 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_191_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_191_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_191_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_192_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_193 ();
 sky130_as_sc_hs__fill_8 FILLER_0_192_197 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_205 ();
 sky130_as_sc_hs__fill_1 FILLER_0_192_209 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_248 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_192_265 ();
 sky130_as_sc_hs__fill_1 FILLER_0_192_27 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_305 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_335 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_342 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_348 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_352 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_360 ();
 sky130_as_sc_hs__fill_1 FILLER_0_192_384 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_401 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_411 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_416 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_428 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_192_467 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_482 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_487 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_499 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_527 ();
 sky130_as_sc_hs__fill_1 FILLER_0_192_544 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_569 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_589 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_61 ();
 sky130_as_sc_hs__fill_1 FILLER_0_192_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_696 ();
 sky130_as_sc_hs__fill_1 FILLER_0_192_744 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_765 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_77 ();
 sky130_as_sc_hs__fill_1 FILLER_0_192_787 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_807 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_192_811 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_192_835 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_839 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_85 ();
 sky130_as_sc_hs__fill_8 FILLER_0_192_855 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_863 ();
 sky130_as_sc_hs__fill_1 FILLER_0_192_867 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_192_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_192_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_192_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_193_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_221 ();
 sky130_as_sc_hs__fill_8 FILLER_0_193_225 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_233 ();
 sky130_as_sc_hs__fill_1 FILLER_0_193_237 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_245 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_260 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_264 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_277 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_193_335 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_353 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_357 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_361 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_369 ();
 sky130_as_sc_hs__fill_1 FILLER_0_193_391 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_398 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_437 ();
 sky130_as_sc_hs__fill_1 FILLER_0_193_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_476 ();
 sky130_as_sc_hs__fill_1 FILLER_0_193_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_193_55 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_554 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_604 ();
 sky130_as_sc_hs__fill_1 FILLER_0_193_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_636 ();
 sky130_as_sc_hs__fill_1 FILLER_0_193_673 ();
 sky130_as_sc_hs__fill_1 FILLER_0_193_682 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_706 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_710 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_714 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_718 ();
 sky130_as_sc_hs__fill_1 FILLER_0_193_722 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_73 ();
 sky130_as_sc_hs__fill_1 FILLER_0_193_756 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_781 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_797 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_818 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_822 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_826 ();
 sky130_as_sc_hs__fill_8 FILLER_0_193_830 ();
 sky130_as_sc_hs__fill_2 FILLER_0_193_838 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_841 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_857 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_873 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_193_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_193_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_193_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_194_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_193 ();
 sky130_as_sc_hs__fill_8 FILLER_0_194_197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_205 ();
 sky130_as_sc_hs__fill_1 FILLER_0_194_251 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_258 ();
 sky130_as_sc_hs__fill_1 FILLER_0_194_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_280 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_306 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_319 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_323 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_354 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_360 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_371 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_394 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_416 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_434 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_440 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_444 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_448 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_45 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_465 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_491 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_510 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_562 ();
 sky130_as_sc_hs__fill_1 FILLER_0_194_608 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_61 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_622 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_666 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_693 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_705 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_730 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_77 ();
 sky130_as_sc_hs__fill_1 FILLER_0_194_780 ();
 sky130_as_sc_hs__fill_1 FILLER_0_194_786 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_194_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_813 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_834 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_85 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_850 ();
 sky130_as_sc_hs__fill_2 FILLER_0_194_866 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_194_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_194_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_194_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_1177 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_1216 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_195_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_244 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_254 ();
 sky130_as_sc_hs__fill_1 FILLER_0_195_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_290 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_294 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_298 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_302 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_306 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_310 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_316 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_320 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_329 ();
 sky130_as_sc_hs__fill_1 FILLER_0_195_333 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_345 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_35 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_353 ();
 sky130_as_sc_hs__fill_1 FILLER_0_195_357 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_364 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_368 ();
 sky130_as_sc_hs__fill_1 FILLER_0_195_406 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_434 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_440 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_444 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_473 ();
 sky130_as_sc_hs__fill_1 FILLER_0_195_491 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_500 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_505 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_509 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_51 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_521 ();
 sky130_as_sc_hs__fill_1 FILLER_0_195_525 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_533 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_538 ();
 sky130_as_sc_hs__fill_1 FILLER_0_195_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_566 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_570 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_574 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_578 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_582 ();
 sky130_as_sc_hs__fill_1 FILLER_0_195_586 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_612 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_646 ();
 sky130_as_sc_hs__fill_1 FILLER_0_195_661 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_666 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_678 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_682 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_686 ();
 sky130_as_sc_hs__fill_1 FILLER_0_195_690 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_696 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_752 ();
 sky130_as_sc_hs__fill_1 FILLER_0_195_773 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_825 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_834 ();
 sky130_as_sc_hs__fill_2 FILLER_0_195_838 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_841 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_857 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_873 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_195_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_195_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_195_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_196_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_196_213 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_225 ();
 sky130_as_sc_hs__fill_1 FILLER_0_196_251 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_268 ();
 sky130_as_sc_hs__fill_1 FILLER_0_196_27 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_283 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_29 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_291 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_299 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_328 ();
 sky130_as_sc_hs__fill_1 FILLER_0_196_363 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_365 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_375 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_381 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_421 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_438 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_444 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_472 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_530 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_552 ();
 sky130_as_sc_hs__fill_1 FILLER_0_196_587 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_593 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_597 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_61 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_619 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_696 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_712 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_727 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_748 ();
 sky130_as_sc_hs__fill_1 FILLER_0_196_755 ();
 sky130_as_sc_hs__fill_1 FILLER_0_196_757 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_777 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_800 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_196_840 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_844 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_85 ();
 sky130_as_sc_hs__fill_8 FILLER_0_196_860 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_196_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_196_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_196_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_1173 ();
 sky130_as_sc_hs__fill_8 FILLER_0_197_1177 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_1185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_1207 ();
 sky130_as_sc_hs__fill_8 FILLER_0_197_1223 ();
 sky130_as_sc_hs__fill_1 FILLER_0_197_1231 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_197_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_221 ();
 sky130_as_sc_hs__fill_8 FILLER_0_197_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_233 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_238 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_242 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_197_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_197_321 ();
 sky130_as_sc_hs__fill_1 FILLER_0_197_335 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_337 ();
 sky130_as_sc_hs__fill_1 FILLER_0_197_341 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_349 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_35 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_385 ();
 sky130_as_sc_hs__fill_1 FILLER_0_197_389 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_401 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_417 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_425 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_454 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_471 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_494 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_197_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_556 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_569 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_197_580 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_613 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_636 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_646 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_669 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_697 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_723 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_733 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_741 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_766 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_770 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_781 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_804 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_846 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_850 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_866 ();
 sky130_as_sc_hs__fill_8 FILLER_0_197_882 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_89 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_890 ();
 sky130_as_sc_hs__fill_2 FILLER_0_197_894 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_197_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_197_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_197_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_101 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_1032 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_1168 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_1184 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_1200 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_198_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_250 ();
 sky130_as_sc_hs__fill_1 FILLER_0_198_266 ();
 sky130_as_sc_hs__fill_1 FILLER_0_198_27 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_286 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_297 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_301 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_305 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_320 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_339 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_376 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_404 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_414 ();
 sky130_as_sc_hs__fill_1 FILLER_0_198_429 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_435 ();
 sky130_as_sc_hs__fill_1 FILLER_0_198_439 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_442 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_451 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_474 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_485 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_528 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_533 ();
 sky130_as_sc_hs__fill_1 FILLER_0_198_537 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_540 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_554 ();
 sky130_as_sc_hs__fill_1 FILLER_0_198_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_583 ();
 sky130_as_sc_hs__fill_1 FILLER_0_198_587 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_632 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_642 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_663 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_667 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_678 ();
 sky130_as_sc_hs__fill_1 FILLER_0_198_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_752 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_762 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_766 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_770 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_774 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_778 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_782 ();
 sky130_as_sc_hs__fill_1 FILLER_0_198_803 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_198_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_198_845 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_85 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_865 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_198_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_198_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_198_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_199_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_221 ();
 sky130_as_sc_hs__fill_8 FILLER_0_199_225 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_233 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_237 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_258 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_295 ();
 sky130_as_sc_hs__fill_1 FILLER_0_199_299 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_332 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_337 ();
 sky130_as_sc_hs__fill_1 FILLER_0_199_341 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_361 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_371 ();
 sky130_as_sc_hs__fill_1 FILLER_0_199_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_415 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_446 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_457 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_463 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_480 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_484 ();
 sky130_as_sc_hs__fill_1 FILLER_0_199_495 ();
 sky130_as_sc_hs__fill_1 FILLER_0_199_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_522 ();
 sky130_as_sc_hs__fill_1 FILLER_0_199_543 ();
 sky130_as_sc_hs__fill_1 FILLER_0_199_55 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_585 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_593 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_598 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_608 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_614 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_663 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_681 ();
 sky130_as_sc_hs__fill_1 FILLER_0_199_685 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_707 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_711 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_73 ();
 sky130_as_sc_hs__fill_1 FILLER_0_199_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_778 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_782 ();
 sky130_as_sc_hs__fill_8 FILLER_0_199_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_793 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_797 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_846 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_850 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_866 ();
 sky130_as_sc_hs__fill_8 FILLER_0_199_882 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_89 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_890 ();
 sky130_as_sc_hs__fill_2 FILLER_0_199_894 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_199_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_199_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_199_985 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_100 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1025 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_104 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1065 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_108 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1121 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1193 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_12 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_19_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_1273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_136 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_142 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_146 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_15 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_150 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_154 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_19 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_191 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_195 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_200 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_204 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_210 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_214 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_218 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_225 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_229 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_23 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_235 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_243 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_247 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_251 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_255 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_262 ();
 sky130_as_sc_hs__fill_8 FILLER_0_19_266 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_274 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_28 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_281 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_32 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_337 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_344 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_364 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_37 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_391 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_393 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_397 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_400 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_43 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_430 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_434 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_47 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_478 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_482 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_495 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_518 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_527 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_532 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_546 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_554 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_558 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_561 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_576 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_584 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_600 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_606 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_612 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_625 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_630 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_634 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_638 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_64 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_643 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_647 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_664 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_671 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_678 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_68 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_682 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_686 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_699 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_703 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_708 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_72 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_76 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_783 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_793 ();
 sky130_as_sc_hs__decap_4 FILLER_0_19_8 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_80 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_805 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_809 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_84 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_860 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_88 ();
 sky130_as_sc_hs__fill_1 FILLER_0_19_890 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_92 ();
 sky130_as_sc_hs__decap_3 FILLER_0_19_922 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_96 ();
 sky130_as_sc_hs__fill_2 FILLER_0_19_961 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_965 ();
 sky130_as_sc_hs__decap_16 FILLER_0_19_981 ();
 sky130_as_sc_hs__fill_8 FILLER_0_19_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_1_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_1025 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_105 ();
 sky130_as_sc_hs__decap_3 FILLER_0_1_1065 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_1084 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_1088 ();
 sky130_as_sc_hs__decap_3 FILLER_0_1_109 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_11 ();
 sky130_as_sc_hs__decap_3 FILLER_0_1_1117 ();
 sky130_as_sc_hs__fill_8 FILLER_0_1_1121 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_1129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_113 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_1157 ();
 sky130_as_sc_hs__fill_8 FILLER_0_1_1161 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_1169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_1196 ();
 sky130_as_sc_hs__fill_8 FILLER_0_1_1220 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_1228 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_1_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_129 ();
 sky130_as_sc_hs__fill_8 FILLER_0_1_145 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_15 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_153 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_157 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_167 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_182 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_186 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_223 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_225 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_245 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_1_277 ();
 sky130_as_sc_hs__fill_8 FILLER_0_1_281 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_289 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_29 ();
 sky130_as_sc_hs__fill_8 FILLER_0_1_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_303 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_307 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_33 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_335 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_337 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_353 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_357 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_371 ();
 sky130_as_sc_hs__fill_8 FILLER_0_1_383 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_391 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_415 ();
 sky130_as_sc_hs__fill_8 FILLER_0_1_432 ();
 sky130_as_sc_hs__decap_3 FILLER_0_1_440 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_457 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_461 ();
 sky130_as_sc_hs__decap_3 FILLER_0_1_472 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_49 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_503 ();
 sky130_as_sc_hs__fill_8 FILLER_0_1_505 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_513 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_539 ();
 sky130_as_sc_hs__fill_8 FILLER_0_1_569 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_577 ();
 sky130_as_sc_hs__decap_3 FILLER_0_1_608 ();
 sky130_as_sc_hs__decap_3 FILLER_0_1_636 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_65 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_668 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_702 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_707 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_711 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_727 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_745 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_761 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_777 ();
 sky130_as_sc_hs__decap_3 FILLER_0_1_781 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_789 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_815 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_819 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_835 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_839 ();
 sky130_as_sc_hs__fill_8 FILLER_0_1_841 ();
 sky130_as_sc_hs__decap_4 FILLER_0_1_849 ();
 sky130_as_sc_hs__decap_3 FILLER_0_1_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_1_883 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_887 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_916 ();
 sky130_as_sc_hs__fill_1 FILLER_0_1_932 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_969 ();
 sky130_as_sc_hs__fill_8 FILLER_0_1_97 ();
 sky130_as_sc_hs__decap_16 FILLER_0_1_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_200_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_197 ();
 sky130_as_sc_hs__fill_8 FILLER_0_200_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_265 ();
 sky130_as_sc_hs__fill_1 FILLER_0_200_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_303 ();
 sky130_as_sc_hs__fill_1 FILLER_0_200_307 ();
 sky130_as_sc_hs__fill_8 FILLER_0_200_309 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_317 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_321 ();
 sky130_as_sc_hs__fill_1 FILLER_0_200_331 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_340 ();
 sky130_as_sc_hs__fill_1 FILLER_0_200_363 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_365 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_381 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_386 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_390 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_410 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_429 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_435 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_439 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_200_462 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_504 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_576 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_582 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_624 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_628 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_642 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_698 ();
 sky130_as_sc_hs__fill_1 FILLER_0_200_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_734 ();
 sky130_as_sc_hs__fill_8 FILLER_0_200_738 ();
 sky130_as_sc_hs__fill_1 FILLER_0_200_746 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_754 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_761 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_765 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_769 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_77 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_783 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_799 ();
 sky130_as_sc_hs__fill_1 FILLER_0_200_803 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_806 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_810 ();
 sky130_as_sc_hs__fill_8 FILLER_0_200_813 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_821 ();
 sky130_as_sc_hs__fill_1 FILLER_0_200_825 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_842 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_846 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_85 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_862 ();
 sky130_as_sc_hs__fill_2 FILLER_0_200_866 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_200_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_200_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_200_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_201_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_221 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_225 ();
 sky130_as_sc_hs__fill_1 FILLER_0_201_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_262 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_266 ();
 sky130_as_sc_hs__fill_8 FILLER_0_201_270 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_294 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_201_316 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_342 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_346 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_350 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_354 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_358 ();
 sky130_as_sc_hs__fill_1 FILLER_0_201_367 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_401 ();
 sky130_as_sc_hs__fill_1 FILLER_0_201_405 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_424 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_465 ();
 sky130_as_sc_hs__fill_1 FILLER_0_201_495 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_531 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_535 ();
 sky130_as_sc_hs__fill_1 FILLER_0_201_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_551 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_555 ();
 sky130_as_sc_hs__fill_1 FILLER_0_201_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_201_586 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_614 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_622 ();
 sky130_as_sc_hs__fill_8 FILLER_0_201_653 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_661 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_665 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_673 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_685 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_725 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_748 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_752 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_781 ();
 sky130_as_sc_hs__fill_2 FILLER_0_201_785 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_789 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_805 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_821 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_837 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_841 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_857 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_873 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_201_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_201_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_201_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_202_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_247 ();
 sky130_as_sc_hs__fill_1 FILLER_0_202_251 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_253 ();
 sky130_as_sc_hs__fill_1 FILLER_0_202_266 ();
 sky130_as_sc_hs__fill_1 FILLER_0_202_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_275 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_279 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_283 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_301 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_305 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_328 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_339 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_361 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_433 ();
 sky130_as_sc_hs__fill_1 FILLER_0_202_437 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_202_465 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_474 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_512 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_516 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_522 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_528 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_557 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_562 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_566 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_571 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_589 ();
 sky130_as_sc_hs__fill_8 FILLER_0_202_593 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_606 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_616 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_642 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_653 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_657 ();
 sky130_as_sc_hs__fill_1 FILLER_0_202_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_693 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_715 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_719 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_741 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_202_781 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_785 ();
 sky130_as_sc_hs__fill_8 FILLER_0_202_801 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_809 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_81 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_813 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_829 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_845 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_85 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_865 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_202_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_202_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_202_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_203_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_255 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_259 ();
 sky130_as_sc_hs__fill_1 FILLER_0_203_286 ();
 sky130_as_sc_hs__fill_1 FILLER_0_203_295 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_315 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_325 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_35 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_364 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_381 ();
 sky130_as_sc_hs__fill_1 FILLER_0_203_385 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_388 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_414 ();
 sky130_as_sc_hs__fill_1 FILLER_0_203_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_435 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_439 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_443 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_449 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_453 ();
 sky130_as_sc_hs__fill_1 FILLER_0_203_457 ();
 sky130_as_sc_hs__fill_1 FILLER_0_203_465 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_501 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_510 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_514 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_518 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_522 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_526 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_547 ();
 sky130_as_sc_hs__fill_1 FILLER_0_203_55 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_557 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_569 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_581 ();
 sky130_as_sc_hs__fill_1 FILLER_0_203_585 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_605 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_614 ();
 sky130_as_sc_hs__fill_1 FILLER_0_203_636 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_642 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_646 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_650 ();
 sky130_as_sc_hs__fill_8 FILLER_0_203_692 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_700 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_704 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_709 ();
 sky130_as_sc_hs__fill_1 FILLER_0_203_713 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_724 ();
 sky130_as_sc_hs__fill_1 FILLER_0_203_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_746 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_761 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_765 ();
 sky130_as_sc_hs__fill_1 FILLER_0_203_769 ();
 sky130_as_sc_hs__fill_2 FILLER_0_203_775 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_779 ();
 sky130_as_sc_hs__fill_1 FILLER_0_203_783 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_785 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_801 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_817 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_833 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_837 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_841 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_857 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_873 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_203_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_203_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_203_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_204_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_213 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_248 ();
 sky130_as_sc_hs__fill_1 FILLER_0_204_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_262 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_266 ();
 sky130_as_sc_hs__fill_1 FILLER_0_204_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_304 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_313 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_327 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_333 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_337 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_341 ();
 sky130_as_sc_hs__fill_1 FILLER_0_204_347 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_405 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_418 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_433 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_437 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_441 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_463 ();
 sky130_as_sc_hs__fill_1 FILLER_0_204_475 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_204_481 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_512 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_516 ();
 sky130_as_sc_hs__fill_8 FILLER_0_204_520 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_528 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_533 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_537 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_553 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_589 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_61 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_619 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_641 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_653 ();
 sky130_as_sc_hs__fill_1 FILLER_0_204_669 ();
 sky130_as_sc_hs__fill_8 FILLER_0_204_691 ();
 sky130_as_sc_hs__fill_1 FILLER_0_204_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_728 ();
 sky130_as_sc_hs__fill_2 FILLER_0_204_732 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_753 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_77 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_784 ();
 sky130_as_sc_hs__fill_8 FILLER_0_204_800 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_808 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_81 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_813 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_829 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_845 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_85 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_865 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_204_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_204_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_204_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_205_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_14 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_225 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_241 ();
 sky130_as_sc_hs__fill_1 FILLER_0_205_245 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_264 ();
 sky130_as_sc_hs__fill_8 FILLER_0_205_268 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_276 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_285 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_297 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_30 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_318 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_334 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_350 ();
 sky130_as_sc_hs__fill_1 FILLER_0_205_372 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_425 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_449 ();
 sky130_as_sc_hs__fill_8 FILLER_0_205_46 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_468 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_472 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_480 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_484 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_488 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_501 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_505 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_509 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_525 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_54 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_547 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_557 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_585 ();
 sky130_as_sc_hs__fill_8 FILLER_0_205_589 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_597 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_601 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_609 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_613 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_617 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_638 ();
 sky130_as_sc_hs__fill_1 FILLER_0_205_642 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_645 ();
 sky130_as_sc_hs__fill_8 FILLER_0_205_661 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_669 ();
 sky130_as_sc_hs__fill_8 FILLER_0_205_673 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_683 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_699 ();
 sky130_as_sc_hs__fill_8 FILLER_0_205_720 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_205_753 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_779 ();
 sky130_as_sc_hs__fill_1 FILLER_0_205_783 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_785 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_801 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_817 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_833 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_837 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_841 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_857 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_873 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_205_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_205_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_205_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_206_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_213 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_229 ();
 sky130_as_sc_hs__fill_1 FILLER_0_206_27 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_272 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_3 ();
 sky130_as_sc_hs__fill_8 FILLER_0_206_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_206_328 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_206_382 ();
 sky130_as_sc_hs__fill_8 FILLER_0_206_386 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_394 ();
 sky130_as_sc_hs__fill_1 FILLER_0_206_400 ();
 sky130_as_sc_hs__fill_8 FILLER_0_206_406 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_414 ();
 sky130_as_sc_hs__fill_2 FILLER_0_206_418 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_421 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_437 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_206_453 ();
 sky130_as_sc_hs__fill_2 FILLER_0_206_474 ();
 sky130_as_sc_hs__fill_2 FILLER_0_206_490 ();
 sky130_as_sc_hs__fill_2 FILLER_0_206_494 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_498 ();
 sky130_as_sc_hs__fill_8 FILLER_0_206_503 ();
 sky130_as_sc_hs__fill_2 FILLER_0_206_511 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_529 ();
 sky130_as_sc_hs__fill_1 FILLER_0_206_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_206_558 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_562 ();
 sky130_as_sc_hs__fill_8 FILLER_0_206_578 ();
 sky130_as_sc_hs__fill_2 FILLER_0_206_586 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_589 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_605 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_61 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_621 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_637 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_641 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_645 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_661 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_677 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_693 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_697 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_701 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_717 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_733 ();
 sky130_as_sc_hs__fill_2 FILLER_0_206_754 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_757 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_77 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_773 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_789 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_805 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_809 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_81 ();
 sky130_as_sc_hs__fill_8 FILLER_0_206_813 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_206_825 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_833 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_85 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_865 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_206_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_206_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_206_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_1156 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_1172 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_207_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_225 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_241 ();
 sky130_as_sc_hs__fill_1 FILLER_0_207_257 ();
 sky130_as_sc_hs__fill_8 FILLER_0_207_268 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_276 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_207_285 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_292 ();
 sky130_as_sc_hs__fill_2 FILLER_0_207_296 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_3 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_35 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_356 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_207_374 ();
 sky130_as_sc_hs__fill_2 FILLER_0_207_378 ();
 sky130_as_sc_hs__fill_8 FILLER_0_207_382 ();
 sky130_as_sc_hs__fill_2 FILLER_0_207_390 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_393 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_409 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_425 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_441 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_445 ();
 sky130_as_sc_hs__fill_8 FILLER_0_207_449 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_457 ();
 sky130_as_sc_hs__fill_2 FILLER_0_207_480 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_484 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_500 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_51 ();
 sky130_as_sc_hs__fill_8 FILLER_0_207_521 ();
 sky130_as_sc_hs__fill_8 FILLER_0_207_531 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_539 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_543 ();
 sky130_as_sc_hs__fill_1 FILLER_0_207_55 ();
 sky130_as_sc_hs__fill_8 FILLER_0_207_551 ();
 sky130_as_sc_hs__fill_1 FILLER_0_207_559 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_57 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_577 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_593 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_609 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_613 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_617 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_633 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_649 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_665 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_669 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_673 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_689 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_705 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_721 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_725 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_73 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_745 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_761 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_777 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_781 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_785 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_801 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_817 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_833 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_837 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_841 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_857 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_873 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_207_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_207_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_207_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_208_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_213 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_229 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_245 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_249 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_253 ();
 sky130_as_sc_hs__fill_1 FILLER_0_208_269 ();
 sky130_as_sc_hs__fill_1 FILLER_0_208_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_289 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_305 ();
 sky130_as_sc_hs__fill_8 FILLER_0_208_309 ();
 sky130_as_sc_hs__fill_1 FILLER_0_208_317 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_323 ();
 sky130_as_sc_hs__fill_2 FILLER_0_208_327 ();
 sky130_as_sc_hs__fill_8 FILLER_0_208_331 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_339 ();
 sky130_as_sc_hs__fill_2 FILLER_0_208_343 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_347 ();
 sky130_as_sc_hs__fill_1 FILLER_0_208_363 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_365 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_371 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_387 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_403 ();
 sky130_as_sc_hs__fill_1 FILLER_0_208_419 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_421 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_437 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_45 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_453 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_469 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_473 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_477 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_493 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_509 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_525 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_529 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_533 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_549 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_565 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_581 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_585 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_589 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_605 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_61 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_621 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_637 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_641 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_645 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_661 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_677 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_693 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_697 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_701 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_717 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_733 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_749 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_753 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_757 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_77 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_773 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_789 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_805 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_809 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_81 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_813 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_829 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_845 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_85 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_865 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_208_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_208_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_208_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_1065 ();
 sky130_as_sc_hs__fill_8 FILLER_0_209_1081 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_1089 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_1100 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_1116 ();
 sky130_as_sc_hs__fill_8 FILLER_0_209_1121 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_1129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_113 ();
 sky130_as_sc_hs__fill_2 FILLER_0_209_1133 ();
 sky130_as_sc_hs__fill_8 FILLER_0_209_1154 ();
 sky130_as_sc_hs__fill_1 FILLER_0_209_1162 ();
 sky130_as_sc_hs__fill_1 FILLER_0_209_1175 ();
 sky130_as_sc_hs__fill_8 FILLER_0_209_1177 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_1185 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_1189 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_1194 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_1210 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_1226 ();
 sky130_as_sc_hs__fill_2 FILLER_0_209_1230 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_209_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_225 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_241 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_277 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_297 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_3 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_313 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_329 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_333 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_35 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_353 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_369 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_385 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_389 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_393 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_409 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_425 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_441 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_445 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_449 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_465 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_481 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_497 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_501 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_51 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_521 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_537 ();
 sky130_as_sc_hs__fill_1 FILLER_0_209_55 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_553 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_557 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_57 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_577 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_593 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_609 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_613 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_617 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_633 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_649 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_665 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_669 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_673 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_689 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_705 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_721 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_725 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_73 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_745 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_761 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_777 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_781 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_785 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_801 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_817 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_833 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_837 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_841 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_857 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_873 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_889 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_89 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_893 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_897 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_913 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_929 ();
 sky130_as_sc_hs__decap_4 FILLER_0_209_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_209_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_209_985 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_10 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1037 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_105 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1093 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_110 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1181 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_119 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_14 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_151 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_162 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_166 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_176 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_18 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_182 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_194 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_197 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_201 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_204 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_208 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_217 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_22 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_247 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_251 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_268 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_272 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_276 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_286 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_29 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_299 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_323 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_34 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_343 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_365 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_38 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_382 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_388 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_394 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_402 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_416 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_429 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_43 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_435 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_457 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_47 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_474 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_501 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_509 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_513 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_529 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_533 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_540 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_554 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_559 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_56 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_589 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_60 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_636 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_643 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_66 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_661 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_697 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_7 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_70 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_701 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_710 ();
 sky130_as_sc_hs__decap_4 FILLER_0_20_73 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_755 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_788 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_79 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_795 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_799 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_811 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_83 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_840 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_844 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_848 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_852 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_866 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_89 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_890 ();
 sky130_as_sc_hs__decap_3 FILLER_0_20_899 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_923 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_93 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_933 ();
 sky130_as_sc_hs__fill_1 FILLER_0_20_947 ();
 sky130_as_sc_hs__fill_2 FILLER_0_20_97 ();
 sky130_as_sc_hs__fill_8 FILLER_0_20_972 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_20_997 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_1033 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_1045 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_105 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_1061 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_1069 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_1075 ();
 sky130_as_sc_hs__fill_1 FILLER_0_210_1091 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_1093 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_11 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_1120 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_1128 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_1143 ();
 sky130_as_sc_hs__fill_1 FILLER_0_210_1169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_210_1193 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_120 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_1228 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_124 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_1244 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_1261 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_141 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_149 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_15 ();
 sky130_as_sc_hs__fill_1 FILLER_0_210_153 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_158 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_162 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_178 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_186 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_190 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_201 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_217 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_225 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_23 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_233 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_245 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_253 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_265 ();
 sky130_as_sc_hs__fill_1 FILLER_0_210_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_272 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_276 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_292 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_313 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_317 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_333 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_341 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_349 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_353 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_361 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_365 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_37 ();
 sky130_as_sc_hs__fill_1 FILLER_0_210_381 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_386 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_390 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_406 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_414 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_418 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_425 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_429 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_445 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_45 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_453 ();
 sky130_as_sc_hs__fill_1 FILLER_0_210_457 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_462 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_466 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_474 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_477 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_49 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_493 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_499 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_503 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_519 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_527 ();
 sky130_as_sc_hs__fill_1 FILLER_0_210_531 ();
 sky130_as_sc_hs__fill_1 FILLER_0_210_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_538 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_542 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_558 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_574 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_582 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_586 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_589 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_605 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_621 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_637 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_641 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_645 ();
 sky130_as_sc_hs__fill_8 FILLER_0_210_65 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_661 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_677 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_693 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_697 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_701 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_717 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_73 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_733 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_749 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_753 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_757 ();
 sky130_as_sc_hs__fill_1 FILLER_0_210_77 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_773 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_789 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_805 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_809 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_82 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_829 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_210_85 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_865 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_885 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_89 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_901 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_210_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_210_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_210_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_1004 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_1009 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_1025 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_1033 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_1037 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_105 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_1055 ();
 sky130_as_sc_hs__fill_1 FILLER_0_211_1063 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_1065 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_1073 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_109 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_1093 ();
 sky130_as_sc_hs__fill_1 FILLER_0_211_11 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_1102 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_1118 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_113 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_1137 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_1145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_1149 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_1173 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_1177 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_1185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_1205 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_121 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_1221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_1229 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_1249 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_1257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_1270 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_1274 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_141 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_157 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_165 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_185 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_193 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_219 ();
 sky130_as_sc_hs__fill_1 FILLER_0_211_223 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_253 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_269 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_277 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_29 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_297 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_305 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_333 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_337 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_345 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_365 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_381 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_389 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_409 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_417 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_429 ();
 sky130_as_sc_hs__fill_1 FILLER_0_211_447 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_449 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_45 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_465 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_473 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_493 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_501 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_505 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_523 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_53 ();
 sky130_as_sc_hs__fill_1 FILLER_0_211_531 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_533 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_541 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_561 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_577 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_585 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_605 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_609 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_613 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_617 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_624 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_640 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_645 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_653 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_657 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_662 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_670 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_673 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_689 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_701 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_717 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_725 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_729 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_733 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_738 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_754 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_757 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_776 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_785 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_801 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_809 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_81 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_816 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_832 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_841 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_85 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_852 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_885 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_890 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_894 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_897 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_913 ();
 sky130_as_sc_hs__decap_3 FILLER_0_211_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_928 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_944 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_953 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_961 ();
 sky130_as_sc_hs__fill_8 FILLER_0_211_966 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_974 ();
 sky130_as_sc_hs__fill_2 FILLER_0_211_978 ();
 sky130_as_sc_hs__decap_16 FILLER_0_211_981 ();
 sky130_as_sc_hs__decap_4 FILLER_0_211_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_21_1002 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_1006 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_21_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1041 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_21_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1065 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_108 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_21_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_21_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_117 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1193 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_12 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1209 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_122 ();
 sky130_as_sc_hs__decap_4 FILLER_0_21_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_1249 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_126 ();
 sky130_as_sc_hs__fill_8 FILLER_0_21_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_21_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_130 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_137 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_142 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_16 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_165 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_173 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_194 ();
 sky130_as_sc_hs__decap_4 FILLER_0_21_20 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_230 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_254 ();
 sky130_as_sc_hs__decap_4 FILLER_0_21_26 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_262 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_269 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_275 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_279 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_286 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_300 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_306 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_32 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_333 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_36 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_369 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_391 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_40 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_439 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_44 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_449 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_462 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_48 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_484 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_501 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_52 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_532 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_559 ();
 sky130_as_sc_hs__decap_4 FILLER_0_21_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_585 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_607 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_626 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_63 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_663 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_667 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_67 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_673 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_685 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_707 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_71 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_729 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_735 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_76 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_767 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_773 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_789 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_8 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_803 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_807 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_818 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_822 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_830 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_85 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_860 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_868 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_879 ();
 sky130_as_sc_hs__decap_3 FILLER_0_21_883 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_89 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_910 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_923 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_93 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_951 ();
 sky130_as_sc_hs__fill_1 FILLER_0_21_961 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_97 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_970 ();
 sky130_as_sc_hs__fill_2 FILLER_0_21_974 ();
 sky130_as_sc_hs__decap_16 FILLER_0_21_978 ();
 sky130_as_sc_hs__fill_8 FILLER_0_21_994 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1013 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_102 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1053 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_106 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1093 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_11 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_110 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_114 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1237 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_1261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_131 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_136 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_15 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_156 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_160 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_19 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_192 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_227 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_232 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_24 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_241 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_248 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_257 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_269 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_302 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_326 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_33 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_334 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_344 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_365 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_37 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_392 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_40 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_403 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_419 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_426 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_435 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_44 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_443 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_448 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_48 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_491 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_495 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_502 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_508 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_512 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_53 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_531 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_533 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_544 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_550 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_555 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_559 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_573 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_584 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_60 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_600 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_606 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_610 ();
 sky130_as_sc_hs__decap_4 FILLER_0_22_624 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_628 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_631 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_64 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_653 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_674 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_678 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_68 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_698 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_72 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_722 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_726 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_76 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_776 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_80 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_806 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_848 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_866 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_877 ();
 sky130_as_sc_hs__decap_3 FILLER_0_22_89 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_920 ();
 sky130_as_sc_hs__fill_1 FILLER_0_22_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_94 ();
 sky130_as_sc_hs__fill_8 FILLER_0_22_970 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_978 ();
 sky130_as_sc_hs__fill_2 FILLER_0_22_98 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_22_997 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_10 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_102 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1065 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_108 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1121 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1177 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_23_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_15 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_152 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_165 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_175 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_179 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_186 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_19 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_190 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_194 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_206 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_210 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_214 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_23 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_259 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_27 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_296 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_307 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_31 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_311 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_333 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_345 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_35 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_353 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_369 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_383 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_39 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_393 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_418 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_43 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_430 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_435 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_449 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_458 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_462 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_465 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_47 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_479 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_486 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_503 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_513 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_529 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_536 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_540 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_543 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_547 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_559 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_561 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_604 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_61 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_617 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_64 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_643 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_647 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_677 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_681 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_685 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_689 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_70 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_711 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_727 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_738 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_74 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_742 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_746 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_754 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_775 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_78 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_789 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_793 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_801 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_82 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_88 ();
 sky130_as_sc_hs__decap_3 FILLER_0_23_902 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_913 ();
 sky130_as_sc_hs__decap_4 FILLER_0_23_92 ();
 sky130_as_sc_hs__fill_1 FILLER_0_23_947 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_957 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_961 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_965 ();
 sky130_as_sc_hs__fill_2 FILLER_0_23_98 ();
 sky130_as_sc_hs__decap_16 FILLER_0_23_981 ();
 sky130_as_sc_hs__fill_8 FILLER_0_23_997 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_100 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1093 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_11 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1125 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_114 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_129 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_132 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_136 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_145 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_15 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_159 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_166 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_174 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_182 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_186 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_19 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_190 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_202 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_206 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_209 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_228 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_23 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_240 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_269 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_29 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_297 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_319 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_325 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_33 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_348 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_352 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_363 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_37 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_370 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_386 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_400 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_436 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_450 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_46 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_492 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_50 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_506 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_519 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_53 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_554 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_565 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_57 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_578 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_584 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_61 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_610 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_627 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_643 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_65 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_650 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_69 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_696 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_72 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_720 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_747 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_755 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_76 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_80 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_803 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_809 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_818 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_834 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_874 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_878 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_882 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_886 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_890 ();
 sky130_as_sc_hs__decap_3 FILLER_0_24_902 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_915 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_919 ();
 sky130_as_sc_hs__fill_1 FILLER_0_24_923 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_930 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_934 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_950 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_954 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_958 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_96 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_962 ();
 sky130_as_sc_hs__fill_8 FILLER_0_24_966 ();
 sky130_as_sc_hs__decap_4 FILLER_0_24_974 ();
 sky130_as_sc_hs__fill_2 FILLER_0_24_978 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_24_997 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_1041 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_25_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_25_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_25_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_1177 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_118 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_1193 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_12 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_1213 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_25_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_25_1273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_129 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_135 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_148 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_16 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_20 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_216 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_25_24 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_241 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_245 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_254 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_262 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_268 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_272 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_293 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_315 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_334 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_337 ();
 sky130_as_sc_hs__decap_4 FILLER_0_25_355 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_359 ();
 sky130_as_sc_hs__decap_4 FILLER_0_25_375 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_379 ();
 sky130_as_sc_hs__decap_4 FILLER_0_25_393 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_404 ();
 sky130_as_sc_hs__decap_4 FILLER_0_25_410 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_414 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_417 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_433 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_445 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_454 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_458 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_462 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_479 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_493 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_499 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_510 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_515 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_519 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_528 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_540 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_55 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_559 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_561 ();
 sky130_as_sc_hs__decap_4 FILLER_0_25_57 ();
 sky130_as_sc_hs__decap_4 FILLER_0_25_599 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_603 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_606 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_61 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_615 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_622 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_627 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_655 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_665 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_677 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_681 ();
 sky130_as_sc_hs__decap_4 FILLER_0_25_69 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_7 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_705 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_712 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_716 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_741 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_745 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_755 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_76 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_761 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_769 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_785 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_80 ();
 sky130_as_sc_hs__fill_1 FILLER_0_25_830 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_836 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_849 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_853 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_865 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_87 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_881 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_893 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_902 ();
 sky130_as_sc_hs__decap_3 FILLER_0_25_933 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_946 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_950 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_953 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_957 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_961 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_965 ();
 sky130_as_sc_hs__fill_2 FILLER_0_25_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_973 ();
 sky130_as_sc_hs__decap_16 FILLER_0_25_989 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_10 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_26_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_26_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1109 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_111 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_26_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_26_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_26_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_1261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_132 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_14 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_155 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_165 ();
 sky130_as_sc_hs__decap_4 FILLER_0_26_18 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_190 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_207 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_225 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_24 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_245 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_251 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_280 ();
 sky130_as_sc_hs__decap_4 FILLER_0_26_29 ();
 sky130_as_sc_hs__decap_4 FILLER_0_26_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_304 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_314 ();
 sky130_as_sc_hs__decap_4 FILLER_0_26_318 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_322 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_33 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_333 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_355 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_373 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_409 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_418 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_430 ();
 sky130_as_sc_hs__decap_4 FILLER_0_26_458 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_46 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_462 ();
 sky130_as_sc_hs__decap_4 FILLER_0_26_470 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_501 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_524 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_530 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_541 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_551 ();
 sky130_as_sc_hs__decap_4 FILLER_0_26_557 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_569 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_589 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_598 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_639 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_653 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_678 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_698 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_713 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_731 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_753 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_77 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_809 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_823 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_866 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_869 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_912 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_923 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_929 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_933 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_949 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_953 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_957 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_961 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_965 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_969 ();
 sky130_as_sc_hs__fill_1 FILLER_0_26_97 ();
 sky130_as_sc_hs__fill_2 FILLER_0_26_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_26_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_26_997 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_1006 ();
 sky130_as_sc_hs__decap_16 FILLER_0_27_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_27_1025 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_104 ();
 sky130_as_sc_hs__decap_16 FILLER_0_27_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_27_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_27_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_27_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_27_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_27_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_27_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_113 ();
 sky130_as_sc_hs__decap_4 FILLER_0_27_1137 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_1141 ();
 sky130_as_sc_hs__fill_8 FILLER_0_27_1163 ();
 sky130_as_sc_hs__decap_4 FILLER_0_27_1171 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_1175 ();
 sky130_as_sc_hs__decap_16 FILLER_0_27_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_27_1193 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_12 ();
 sky130_as_sc_hs__decap_16 FILLER_0_27_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_27_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_27_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_27_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_27_1265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_127 ();
 sky130_as_sc_hs__decap_4 FILLER_0_27_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_134 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_138 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_27_16 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_165 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_173 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_192 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_206 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_22 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_26 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_264 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_268 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_291 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_295 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_299 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_30 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_317 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_325 ();
 sky130_as_sc_hs__decap_4 FILLER_0_27_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_34 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_341 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_344 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_369 ();
 sky130_as_sc_hs__decap_4 FILLER_0_27_382 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_388 ();
 sky130_as_sc_hs__decap_4 FILLER_0_27_432 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_443 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_449 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_474 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_488 ();
 sky130_as_sc_hs__decap_4 FILLER_0_27_498 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_505 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_528 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_53 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_546 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_57 ();
 sky130_as_sc_hs__decap_4 FILLER_0_27_577 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_583 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_602 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_608 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_634 ();
 sky130_as_sc_hs__decap_4 FILLER_0_27_64 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_644 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_649 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_700 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_726 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_733 ();
 sky130_as_sc_hs__decap_3 FILLER_0_27_743 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_751 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_755 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_789 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_79 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_797 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_8 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_811 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_822 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_835 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_860 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_864 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_895 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_90 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_915 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_936 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_942 ();
 sky130_as_sc_hs__fill_1 FILLER_0_27_946 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_966 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_970 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_974 ();
 sky130_as_sc_hs__fill_2 FILLER_0_27_978 ();
 sky130_as_sc_hs__decap_16 FILLER_0_27_982 ();
 sky130_as_sc_hs__fill_8 FILLER_0_27_998 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1005 ();
 sky130_as_sc_hs__fill_8 FILLER_0_28_1021 ();
 sky130_as_sc_hs__decap_4 FILLER_0_28_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_28_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1093 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_11 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_110 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_28_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1165 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_28_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_28_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_28_127 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_131 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_139 ();
 sky130_as_sc_hs__decap_4 FILLER_0_28_141 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_145 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_15 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_153 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_190 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_20 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_212 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_226 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_24 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_275 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_279 ();
 sky130_as_sc_hs__decap_4 FILLER_0_28_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_306 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_313 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_317 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_326 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_33 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_332 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_336 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_352 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_369 ();
 sky130_as_sc_hs__decap_4 FILLER_0_28_381 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_395 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_400 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_41 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_414 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_430 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_473 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_483 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_531 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_533 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_540 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_560 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_566 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_586 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_602 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_606 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_619 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_628 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_63 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_673 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_69 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_705 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_735 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_739 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_754 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_775 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_790 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_804 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_856 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_863 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_882 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_902 ();
 sky130_as_sc_hs__decap_3 FILLER_0_28_911 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_922 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_93 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_937 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_955 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_959 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_963 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_967 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_971 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_975 ();
 sky130_as_sc_hs__fill_1 FILLER_0_28_979 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_981 ();
 sky130_as_sc_hs__fill_2 FILLER_0_28_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_28_989 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_1006 ();
 sky130_as_sc_hs__decap_16 FILLER_0_29_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_29_1025 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_1029 ();
 sky130_as_sc_hs__fill_8 FILLER_0_29_1050 ();
 sky130_as_sc_hs__decap_4 FILLER_0_29_1058 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_29_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_29_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_29_1097 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_11 ();
 sky130_as_sc_hs__decap_4 FILLER_0_29_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_29_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_29_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_29_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_29_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_1173 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_29_1197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_29_1213 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_1229 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_29_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_29_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_29_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_29_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_15 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_163 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_174 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_182 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_189 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_19 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_193 ();
 sky130_as_sc_hs__fill_1 FILLER_0_29_218 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_23 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_263 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_27 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_286 ();
 sky130_as_sc_hs__fill_1 FILLER_0_29_290 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_311 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_330 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_334 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_347 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_367 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_374 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_379 ();
 sky130_as_sc_hs__decap_4 FILLER_0_29_401 ();
 sky130_as_sc_hs__fill_1 FILLER_0_29_405 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_416 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_427 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_446 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_453 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_46 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_486 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_501 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_505 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_516 ();
 sky130_as_sc_hs__fill_1 FILLER_0_29_543 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_549 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_557 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_561 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_565 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_579 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_583 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_587 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_599 ();
 sky130_as_sc_hs__fill_1 FILLER_0_29_643 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_649 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_663 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_670 ();
 sky130_as_sc_hs__fill_1 FILLER_0_29_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_709 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_748 ();
 sky130_as_sc_hs__fill_1 FILLER_0_29_775 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_822 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_889 ();
 sky130_as_sc_hs__fill_1 FILLER_0_29_921 ();
 sky130_as_sc_hs__decap_3 FILLER_0_29_930 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_962 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_966 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_970 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_974 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_978 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_982 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_986 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_990 ();
 sky130_as_sc_hs__fill_2 FILLER_0_29_994 ();
 sky130_as_sc_hs__fill_8 FILLER_0_29_998 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_1029 ();
 sky130_as_sc_hs__fill_1 FILLER_0_2_1033 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_1037 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_1049 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_1053 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_1057 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_1074 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_1090 ();
 sky130_as_sc_hs__fill_8 FILLER_0_2_1098 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_11 ();
 sky130_as_sc_hs__fill_1 FILLER_0_2_1106 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_1111 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_1115 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_1131 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_1135 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_1157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_117 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_1200 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_1224 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_1240 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_1256 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_15 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_189 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_193 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_201 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_209 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_213 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_229 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_23 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_245 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_249 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_253 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_269 ();
 sky130_as_sc_hs__fill_1 FILLER_0_2_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_285 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_29 ();
 sky130_as_sc_hs__fill_8 FILLER_0_2_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_301 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_305 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_309 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_325 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_341 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_357 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_361 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_365 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_377 ();
 sky130_as_sc_hs__fill_8 FILLER_0_2_393 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_401 ();
 sky130_as_sc_hs__fill_1 FILLER_0_2_421 ();
 sky130_as_sc_hs__fill_8 FILLER_0_2_442 ();
 sky130_as_sc_hs__fill_8 FILLER_0_2_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_450 ();
 sky130_as_sc_hs__fill_8 FILLER_0_2_462 ();
 sky130_as_sc_hs__fill_1 FILLER_0_2_470 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_2_485 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_492 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_508 ();
 sky130_as_sc_hs__fill_8 FILLER_0_2_524 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_53 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_533 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_549 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_565 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_569 ();
 sky130_as_sc_hs__fill_1 FILLER_0_2_575 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_58 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_581 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_610 ();
 sky130_as_sc_hs__fill_1 FILLER_0_2_617 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_645 ();
 sky130_as_sc_hs__fill_1 FILLER_0_2_649 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_656 ();
 sky130_as_sc_hs__fill_1 FILLER_0_2_660 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_666 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_693 ();
 sky130_as_sc_hs__fill_1 FILLER_0_2_697 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_701 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_720 ();
 sky130_as_sc_hs__fill_8 FILLER_0_2_736 ();
 sky130_as_sc_hs__fill_8 FILLER_0_2_74 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_744 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_753 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_757 ();
 sky130_as_sc_hs__fill_8 FILLER_0_2_773 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_781 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_790 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_809 ();
 sky130_as_sc_hs__fill_2 FILLER_0_2_82 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_832 ();
 sky130_as_sc_hs__fill_1 FILLER_0_2_848 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_2_869 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_908 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_2_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_2_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_2_997 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_1001 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1005 ();
 sky130_as_sc_hs__fill_8 FILLER_0_30_1021 ();
 sky130_as_sc_hs__decap_4 FILLER_0_30_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_30_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1093 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_11 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_30_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_30_1197 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_120 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_30_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_30_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_136 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_145 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_15 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_158 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_162 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_166 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_180 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_19 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_222 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_231 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_250 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_275 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_279 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_294 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_320 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_330 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_334 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_353 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_370 ();
 sky130_as_sc_hs__decap_4 FILLER_0_30_387 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_398 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_404 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_418 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_43 ();
 sky130_as_sc_hs__decap_4 FILLER_0_30_445 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_47 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_490 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_501 ();
 sky130_as_sc_hs__decap_4 FILLER_0_30_513 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_517 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_520 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_524 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_528 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_565 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_572 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_584 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_601 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_61 ();
 sky130_as_sc_hs__decap_4 FILLER_0_30_619 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_630 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_641 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_645 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_681 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_7 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_720 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_734 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_74 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_745 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_757 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_770 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_776 ();
 sky130_as_sc_hs__decap_3 FILLER_0_30_796 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_80 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_811 ();
 sky130_as_sc_hs__decap_4 FILLER_0_30_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_867 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_89 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_892 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_898 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_912 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_92 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_949 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_959 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_96 ();
 sky130_as_sc_hs__fill_1 FILLER_0_30_973 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_978 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_985 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_989 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_993 ();
 sky130_as_sc_hs__fill_2 FILLER_0_30_997 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_1007 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_1009 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1013 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1029 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1045 ();
 sky130_as_sc_hs__decap_4 FILLER_0_31_105 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1081 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_31_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_31_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1193 ();
 sky130_as_sc_hs__decap_4 FILLER_0_31_12 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_31_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_31_1249 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_125 ();
 sky130_as_sc_hs__fill_8 FILLER_0_31_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_31_1273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_134 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_140 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_144 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_148 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_155 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_16 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_183 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_19 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_23 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_264 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_278 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_31 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_326 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_332 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_353 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_370 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_378 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_388 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_393 ();
 sky130_as_sc_hs__decap_4 FILLER_0_31_415 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_419 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_435 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_439 ();
 sky130_as_sc_hs__decap_4 FILLER_0_31_462 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_466 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_469 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_477 ();
 sky130_as_sc_hs__decap_4 FILLER_0_31_486 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_492 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_496 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_500 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_505 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_545 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_55 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_554 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_561 ();
 sky130_as_sc_hs__decap_4 FILLER_0_31_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_577 ();
 sky130_as_sc_hs__decap_4 FILLER_0_31_610 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_622 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_626 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_630 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_667 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_673 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_708 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_716 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_722 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_726 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_729 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_745 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_8 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_83 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_870 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_874 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_902 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_915 ();
 sky130_as_sc_hs__decap_3 FILLER_0_31_949 ();
 sky130_as_sc_hs__decap_4 FILLER_0_31_95 ();
 sky130_as_sc_hs__fill_2 FILLER_0_31_957 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_963 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_983 ();
 sky130_as_sc_hs__fill_1 FILLER_0_31_988 ();
 sky130_as_sc_hs__decap_4 FILLER_0_32_10 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_1013 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1017 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_32_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1109 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_111 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_32_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_32_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_32_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_32_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_146 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_16 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_168 ();
 sky130_as_sc_hs__decap_4 FILLER_0_32_181 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_187 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_20 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_202 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_206 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_210 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_216 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_221 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_231 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_238 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_24 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_246 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_295 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_299 ();
 sky130_as_sc_hs__decap_4 FILLER_0_32_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_303 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_307 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_318 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_340 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_344 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_387 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_391 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_416 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_426 ();
 sky130_as_sc_hs__decap_4 FILLER_0_32_43 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_443 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_450 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_47 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_50 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_508 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_519 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_530 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_541 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_554 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_567 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_579 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_597 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_608 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_628 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_642 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_645 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_661 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_686 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_69 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_705 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_709 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_732 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_76 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_80 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_809 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_817 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_828 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_853 ();
 sky130_as_sc_hs__decap_3 FILLER_0_32_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_864 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_882 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_894 ();
 sky130_as_sc_hs__fill_2 FILLER_0_32_898 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_909 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_919 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_939 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_959 ();
 sky130_as_sc_hs__fill_1 FILLER_0_32_979 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_10 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_1017 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_1021 ();
 sky130_as_sc_hs__decap_16 FILLER_0_33_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_33_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_33_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_33_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_33_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_33_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_33_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_33_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_33_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_33_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_33_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_33_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_33_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_33_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_33_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_1229 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_33_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_33_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_33_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_33_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_138 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_14 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_146 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_160 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_18 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_184 ();
 sky130_as_sc_hs__fill_1 FILLER_0_33_191 ();
 sky130_as_sc_hs__fill_1 FILLER_0_33_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_203 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_207 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_22 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_26 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_276 ();
 sky130_as_sc_hs__fill_1 FILLER_0_33_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_287 ();
 sky130_as_sc_hs__fill_1 FILLER_0_33_296 ();
 sky130_as_sc_hs__decap_4 FILLER_0_33_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_302 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_306 ();
 sky130_as_sc_hs__fill_1 FILLER_0_33_310 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_321 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_325 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_331 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_347 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_374 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_393 ();
 sky130_as_sc_hs__fill_1 FILLER_0_33_40 ();
 sky130_as_sc_hs__decap_4 FILLER_0_33_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_419 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_445 ();
 sky130_as_sc_hs__decap_4 FILLER_0_33_464 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_486 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_490 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_510 ();
 sky130_as_sc_hs__fill_1 FILLER_0_33_522 ();
 sky130_as_sc_hs__fill_1 FILLER_0_33_528 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_537 ();
 sky130_as_sc_hs__fill_1 FILLER_0_33_549 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_566 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_575 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_584 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_599 ();
 sky130_as_sc_hs__fill_1 FILLER_0_33_615 ();
 sky130_as_sc_hs__decap_4 FILLER_0_33_62 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_635 ();
 sky130_as_sc_hs__fill_1 FILLER_0_33_671 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_682 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_694 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_698 ();
 sky130_as_sc_hs__fill_1 FILLER_0_33_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_714 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_720 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_724 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_729 ();
 sky130_as_sc_hs__fill_1 FILLER_0_33_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_733 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_741 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_745 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_749 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_790 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_824 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_84 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_846 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_885 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_889 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_893 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_916 ();
 sky130_as_sc_hs__decap_3 FILLER_0_33_93 ();
 sky130_as_sc_hs__fill_2 FILLER_0_33_98 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_10 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_1020 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_1024 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_1028 ();
 sky130_as_sc_hs__decap_4 FILLER_0_34_1032 ();
 sky130_as_sc_hs__decap_16 FILLER_0_34_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_34_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_34_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_34_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_34_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_34_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_34_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_34_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_34_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_34_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_34_1168 ();
 sky130_as_sc_hs__decap_16 FILLER_0_34_1184 ();
 sky130_as_sc_hs__decap_4 FILLER_0_34_1200 ();
 sky130_as_sc_hs__decap_16 FILLER_0_34_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_34_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_34_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_34_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_34_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_34_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_14 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_34_163 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_224 ();
 sky130_as_sc_hs__fill_1 FILLER_0_34_233 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_243 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_297 ();
 sky130_as_sc_hs__decap_4 FILLER_0_34_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_301 ();
 sky130_as_sc_hs__fill_1 FILLER_0_34_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_320 ();
 sky130_as_sc_hs__decap_3 FILLER_0_34_332 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_350 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_39 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_390 ();
 sky130_as_sc_hs__decap_3 FILLER_0_34_434 ();
 sky130_as_sc_hs__decap_3 FILLER_0_34_439 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_464 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_34_503 ();
 sky130_as_sc_hs__decap_4 FILLER_0_34_538 ();
 sky130_as_sc_hs__decap_4 FILLER_0_34_559 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_565 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_610 ();
 sky130_as_sc_hs__fill_1 FILLER_0_34_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_628 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_632 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_636 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_640 ();
 sky130_as_sc_hs__decap_3 FILLER_0_34_645 ();
 sky130_as_sc_hs__decap_4 FILLER_0_34_653 ();
 sky130_as_sc_hs__fill_1 FILLER_0_34_657 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_669 ();
 sky130_as_sc_hs__fill_1 FILLER_0_34_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_722 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_743 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_747 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_751 ();
 sky130_as_sc_hs__fill_1 FILLER_0_34_755 ();
 sky130_as_sc_hs__fill_1 FILLER_0_34_757 ();
 sky130_as_sc_hs__fill_1 FILLER_0_34_763 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_769 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_790 ();
 sky130_as_sc_hs__fill_1 FILLER_0_34_794 ();
 sky130_as_sc_hs__fill_1 FILLER_0_34_800 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_806 ();
 sky130_as_sc_hs__decap_3 FILLER_0_34_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_817 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_821 ();
 sky130_as_sc_hs__fill_1 FILLER_0_34_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_854 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_866 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_901 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_91 ();
 sky130_as_sc_hs__decap_3 FILLER_0_34_921 ();
 sky130_as_sc_hs__fill_1 FILLER_0_34_930 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_952 ();
 sky130_as_sc_hs__fill_2 FILLER_0_34_973 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_1026 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_1030 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_1034 ();
 sky130_as_sc_hs__decap_16 FILLER_0_35_1038 ();
 sky130_as_sc_hs__fill_8 FILLER_0_35_1054 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_35_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_35_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_35_1097 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_11 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_111 ();
 sky130_as_sc_hs__decap_4 FILLER_0_35_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_35_1121 ();
 sky130_as_sc_hs__decap_4 FILLER_0_35_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_35_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_35_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_35_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_35_1177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_119 ();
 sky130_as_sc_hs__decap_16 FILLER_0_35_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_35_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_35_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_1229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_35_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_35_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_35_1265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_127 ();
 sky130_as_sc_hs__decap_4 FILLER_0_35_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_14 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_153 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_157 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_165 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_176 ();
 sky130_as_sc_hs__decap_4 FILLER_0_35_185 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_191 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_215 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_219 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_223 ();
 sky130_as_sc_hs__decap_4 FILLER_0_35_23 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_263 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_29 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_315 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_33 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_333 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_342 ();
 sky130_as_sc_hs__decap_4 FILLER_0_35_349 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_353 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_369 ();
 sky130_as_sc_hs__decap_4 FILLER_0_35_378 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_38 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_384 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_388 ();
 sky130_as_sc_hs__decap_4 FILLER_0_35_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_404 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_42 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_422 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_431 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_436 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_464 ();
 sky130_as_sc_hs__decap_4 FILLER_0_35_474 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_480 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_484 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_488 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_492 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_501 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_518 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_523 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_558 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_587 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_596 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_62 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_628 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_632 ();
 sky130_as_sc_hs__decap_4 FILLER_0_35_652 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_658 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_66 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_662 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_666 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_679 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_683 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_692 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_696 ();
 sky130_as_sc_hs__decap_4 FILLER_0_35_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_700 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_704 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_710 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_714 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_718 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_734 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_738 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_759 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_781 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_80 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_803 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_826 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_830 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_834 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_851 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_855 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_868 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_895 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_90 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_906 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_912 ();
 sky130_as_sc_hs__decap_3 FILLER_0_35_949 ();
 sky130_as_sc_hs__fill_1 FILLER_0_35_972 ();
 sky130_as_sc_hs__fill_2 FILLER_0_35_978 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_1008 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_1032 ();
 sky130_as_sc_hs__decap_16 FILLER_0_36_1037 ();
 sky130_as_sc_hs__fill_8 FILLER_0_36_1053 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_1061 ();
 sky130_as_sc_hs__fill_8 FILLER_0_36_1082 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_1090 ();
 sky130_as_sc_hs__decap_16 FILLER_0_36_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_36_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_36_1125 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_113 ();
 sky130_as_sc_hs__decap_4 FILLER_0_36_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_36_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_36_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_36_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_36_1197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_12 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_36_1205 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_36_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_36_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_36_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_1257 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_126 ();
 sky130_as_sc_hs__decap_16 FILLER_0_36_1261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_135 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_148 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_152 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_156 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_160 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_164 ();
 sky130_as_sc_hs__fill_1 FILLER_0_36_195 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_197 ();
 sky130_as_sc_hs__decap_4 FILLER_0_36_205 ();
 sky130_as_sc_hs__fill_1 FILLER_0_36_209 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_240 ();
 sky130_as_sc_hs__fill_1 FILLER_0_36_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_250 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_26 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_263 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_267 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_274 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_285 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_289 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_293 ();
 sky130_as_sc_hs__fill_1 FILLER_0_36_297 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_322 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_326 ();
 sky130_as_sc_hs__decap_4 FILLER_0_36_330 ();
 sky130_as_sc_hs__fill_1 FILLER_0_36_334 ();
 sky130_as_sc_hs__fill_1 FILLER_0_36_342 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_361 ();
 sky130_as_sc_hs__decap_4 FILLER_0_36_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_376 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_380 ();
 sky130_as_sc_hs__decap_4 FILLER_0_36_402 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_416 ();
 sky130_as_sc_hs__decap_4 FILLER_0_36_421 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_43 ();
 sky130_as_sc_hs__decap_4 FILLER_0_36_432 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_438 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_468 ();
 sky130_as_sc_hs__decap_4 FILLER_0_36_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_528 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_533 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_548 ();
 sky130_as_sc_hs__decap_4 FILLER_0_36_556 ();
 sky130_as_sc_hs__fill_1 FILLER_0_36_570 ();
 sky130_as_sc_hs__fill_1 FILLER_0_36_576 ();
 sky130_as_sc_hs__fill_1 FILLER_0_36_582 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_606 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_624 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_635 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_67 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_710 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_714 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_718 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_735 ();
 sky130_as_sc_hs__decap_4 FILLER_0_36_74 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_754 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_766 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_770 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_8 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_80 ();
 sky130_as_sc_hs__fill_1 FILLER_0_36_811 ();
 sky130_as_sc_hs__fill_1 FILLER_0_36_821 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_36_867 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_869 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_892 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_957 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_978 ();
 sky130_as_sc_hs__decap_3 FILLER_0_36_985 ();
 sky130_as_sc_hs__fill_2 FILLER_0_36_99 ();
 sky130_as_sc_hs__fill_1 FILLER_0_36_998 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_1005 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_1009 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_1038 ();
 sky130_as_sc_hs__decap_16 FILLER_0_37_1042 ();
 sky130_as_sc_hs__decap_4 FILLER_0_37_1058 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_37_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_37_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_37_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_37_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_37_1121 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_37_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_37_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_37_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_37_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_37_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_37_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_37_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_37_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_37_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_37_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_37_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_134 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_15 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_162 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_178 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_185 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_219 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_223 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_238 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_242 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_246 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_250 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_263 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_27 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_274 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_293 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_297 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_301 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_310 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_321 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_345 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_357 ();
 sky130_as_sc_hs__decap_4 FILLER_0_37_382 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_388 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_401 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_407 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_419 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_428 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_439 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_449 ();
 sky130_as_sc_hs__decap_4 FILLER_0_37_485 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_491 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_500 ();
 sky130_as_sc_hs__decap_4 FILLER_0_37_513 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_517 ();
 sky130_as_sc_hs__decap_4 FILLER_0_37_535 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_569 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_595 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_612 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_617 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_653 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_681 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_687 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_709 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_713 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_726 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_729 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_746 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_768 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_785 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_789 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_804 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_815 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_860 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_87 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_876 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_902 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_37_93 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_949 ();
 sky130_as_sc_hs__fill_1 FILLER_0_37_953 ();
 sky130_as_sc_hs__decap_3 FILLER_0_37_966 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_1010 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_1033 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_1037 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_1041 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_1045 ();
 sky130_as_sc_hs__decap_16 FILLER_0_38_1049 ();
 sky130_as_sc_hs__decap_4 FILLER_0_38_105 ();
 sky130_as_sc_hs__decap_16 FILLER_0_38_1065 ();
 sky130_as_sc_hs__fill_8 FILLER_0_38_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_38_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_38_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_38_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_38_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_38_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_38_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_38_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_38_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_38_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_38_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_38_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_38_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_1257 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_126 ();
 sky130_as_sc_hs__decap_16 FILLER_0_38_1261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_137 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_146 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_180 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_186 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_190 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_194 ();
 sky130_as_sc_hs__decap_4 FILLER_0_38_197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_20 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_201 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_204 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_223 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_231 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_235 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_251 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_268 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_282 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_38_34 ();
 sky130_as_sc_hs__decap_4 FILLER_0_38_342 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_353 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_363 ();
 sky130_as_sc_hs__decap_4 FILLER_0_38_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_386 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_396 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_419 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_421 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_428 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_441 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_464 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_474 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_49 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_500 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_515 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_520 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_524 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_528 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_546 ();
 sky130_as_sc_hs__decap_4 FILLER_0_38_552 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_558 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_562 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_567 ();
 sky130_as_sc_hs__decap_4 FILLER_0_38_581 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_585 ();
 sky130_as_sc_hs__decap_4 FILLER_0_38_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_59 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_593 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_606 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_611 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_629 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_645 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_651 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_66 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_686 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_690 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_694 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_731 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_738 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_74 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_745 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_757 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_772 ();
 sky130_as_sc_hs__decap_4 FILLER_0_38_792 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_796 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_799 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_811 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_817 ();
 sky130_as_sc_hs__decap_4 FILLER_0_38_843 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_849 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_854 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_867 ();
 sky130_as_sc_hs__decap_3 FILLER_0_38_92 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_923 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_940 ();
 sky130_as_sc_hs__fill_2 FILLER_0_38_974 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_981 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_987 ();
 sky130_as_sc_hs__fill_1 FILLER_0_38_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_39_10 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_1006 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_1027 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_1031 ();
 sky130_as_sc_hs__decap_4 FILLER_0_39_105 ();
 sky130_as_sc_hs__fill_8 FILLER_0_39_1052 ();
 sky130_as_sc_hs__decap_4 FILLER_0_39_1060 ();
 sky130_as_sc_hs__decap_16 FILLER_0_39_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_39_1081 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_39_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_39_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_39_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_39_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_39_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_39_1169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_117 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_39_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_39_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_39_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_39_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_39_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_39_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_39_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_39_1273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_131 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_142 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_160 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_202 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_210 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_251 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_263 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_274 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_293 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_297 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_30 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_301 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_305 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_313 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_317 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_321 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_325 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_329 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_333 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_337 ();
 sky130_as_sc_hs__decap_4 FILLER_0_39_341 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_377 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_389 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_411 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_426 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_440 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_446 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_481 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_515 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_536 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_542 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_547 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_559 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_566 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_571 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_577 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_584 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_598 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_615 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_638 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_649 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_655 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_70 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_704 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_74 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_762 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_776 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_78 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_780 ();
 sky130_as_sc_hs__decap_4 FILLER_0_39_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_791 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_82 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_833 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_850 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_856 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_894 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_897 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_914 ();
 sky130_as_sc_hs__fill_2 FILLER_0_39_950 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_982 ();
 sky130_as_sc_hs__decap_3 FILLER_0_39_988 ();
 sky130_as_sc_hs__fill_1 FILLER_0_39_99 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_1173 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_1177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_1186 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_1194 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_1211 ();
 sky130_as_sc_hs__fill_8 FILLER_0_3_1217 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_3_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_225 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_241 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_277 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_297 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_3 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_313 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_329 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_333 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_35 ();
 sky130_as_sc_hs__fill_8 FILLER_0_3_353 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_361 ();
 sky130_as_sc_hs__fill_8 FILLER_0_3_368 ();
 sky130_as_sc_hs__fill_1 FILLER_0_3_386 ();
 sky130_as_sc_hs__fill_8 FILLER_0_3_398 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_406 ();
 sky130_as_sc_hs__fill_1 FILLER_0_3_410 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_421 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_439 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_454 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_470 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_3_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_51 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_530 ();
 sky130_as_sc_hs__fill_8 FILLER_0_3_546 ();
 sky130_as_sc_hs__fill_1 FILLER_0_3_55 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_554 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_3_597 ();
 sky130_as_sc_hs__fill_1 FILLER_0_3_603 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_609 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_636 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_655 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_663 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_670 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_673 ();
 sky130_as_sc_hs__fill_8 FILLER_0_3_681 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_689 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_713 ();
 sky130_as_sc_hs__fill_8 FILLER_0_3_717 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_725 ();
 sky130_as_sc_hs__fill_8 FILLER_0_3_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_73 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_741 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_772 ();
 sky130_as_sc_hs__fill_1 FILLER_0_3_783 ();
 sky130_as_sc_hs__fill_1 FILLER_0_3_825 ();
 sky130_as_sc_hs__fill_8 FILLER_0_3_830 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_838 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_841 ();
 sky130_as_sc_hs__fill_1 FILLER_0_3_845 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_89 ();
 sky130_as_sc_hs__fill_2 FILLER_0_3_894 ();
 sky130_as_sc_hs__fill_1 FILLER_0_3_901 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_921 ();
 sky130_as_sc_hs__fill_8 FILLER_0_3_937 ();
 sky130_as_sc_hs__decap_4 FILLER_0_3_945 ();
 sky130_as_sc_hs__decap_3 FILLER_0_3_949 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_3_985 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_1034 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_1037 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_1041 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_1045 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_1049 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_105 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_1053 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_1057 ();
 sky130_as_sc_hs__decap_16 FILLER_0_40_1061 ();
 sky130_as_sc_hs__fill_8 FILLER_0_40_1077 ();
 sky130_as_sc_hs__decap_4 FILLER_0_40_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_1089 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_40_1113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_40_1129 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_40_1149 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_116 ();
 sky130_as_sc_hs__decap_16 FILLER_0_40_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_40_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_40_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_12 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_40_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_40_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_40_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_40_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_40_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_129 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_138 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_171 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_175 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_180 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_184 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_205 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_209 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_227 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_231 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_240 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_25 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_251 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_279 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_291 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_297 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_331 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_335 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_339 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_343 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_361 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_371 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_375 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_387 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_39 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_403 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_417 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_437 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_454 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_46 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_473 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_495 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_528 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_546 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_555 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_577 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_586 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_605 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_613 ();
 sky130_as_sc_hs__decap_4 FILLER_0_40_622 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_626 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_63 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_642 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_666 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_681 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_713 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_730 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_734 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_738 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_742 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_746 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_751 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_755 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_765 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_772 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_801 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_82 ();
 sky130_as_sc_hs__fill_1 FILLER_0_40_832 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_866 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_882 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_889 ();
 sky130_as_sc_hs__decap_3 FILLER_0_40_90 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_915 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_922 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_929 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_969 ();
 sky130_as_sc_hs__fill_2 FILLER_0_40_986 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_1006 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_1042 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_1046 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_1050 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_1054 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_1058 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_41_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_41_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_41_1097 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_11 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_41_1121 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_41_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_41_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_41_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_41_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_41_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_41_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_41_1249 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_126 ();
 sky130_as_sc_hs__fill_8 FILLER_0_41_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_132 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_136 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_154 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_158 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_162 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_169 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_175 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_191 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_203 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_230 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_307 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_314 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_342 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_355 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_366 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_37 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_374 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_382 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_388 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_398 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_402 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_405 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_417 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_42 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_433 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_453 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_462 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_488 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_496 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_500 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_513 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_531 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_547 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_553 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_557 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_569 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_576 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_595 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_606 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_612 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_622 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_628 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_670 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_7 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_706 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_711 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_718 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_726 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_729 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_735 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_749 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_764 ();
 sky130_as_sc_hs__decap_3 FILLER_0_41_779 ();
 sky130_as_sc_hs__decap_4 FILLER_0_41_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_791 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_795 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_822 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_829 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_846 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_87 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_905 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_927 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_94 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_968 ();
 sky130_as_sc_hs__fill_2 FILLER_0_41_98 ();
 sky130_as_sc_hs__fill_1 FILLER_0_41_984 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_103 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_1045 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_1049 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_1053 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_1057 ();
 sky130_as_sc_hs__decap_16 FILLER_0_42_1061 ();
 sky130_as_sc_hs__fill_8 FILLER_0_42_1077 ();
 sky130_as_sc_hs__decap_4 FILLER_0_42_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_1089 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_42_1114 ();
 sky130_as_sc_hs__decap_16 FILLER_0_42_1130 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_114 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_1146 ();
 sky130_as_sc_hs__decap_16 FILLER_0_42_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_42_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_42_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_42_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_42_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_42_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_42_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_42_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_42_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_131 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_141 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_174 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_185 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_193 ();
 sky130_as_sc_hs__decap_4 FILLER_0_42_202 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_206 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_214 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_218 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_226 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_230 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_285 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_299 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_303 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_307 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_330 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_379 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_388 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_399 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_419 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_430 ();
 sky130_as_sc_hs__decap_4 FILLER_0_42_44 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_455 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_48 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_486 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_492 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_499 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_510 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_521 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_540 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_565 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_593 ();
 sky130_as_sc_hs__decap_4 FILLER_0_42_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_613 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_643 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_65 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_664 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_689 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_693 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_705 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_724 ();
 sky130_as_sc_hs__decap_4 FILLER_0_42_73 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_751 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_762 ();
 sky130_as_sc_hs__decap_4 FILLER_0_42_785 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_792 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_796 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_809 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_818 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_867 ();
 sky130_as_sc_hs__fill_1 FILLER_0_42_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_875 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_896 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_903 ();
 sky130_as_sc_hs__decap_3 FILLER_0_42_940 ();
 sky130_as_sc_hs__fill_2 FILLER_0_42_959 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_1052 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_1056 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_1060 ();
 sky130_as_sc_hs__decap_16 FILLER_0_43_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_43_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_43_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_43_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_43_1121 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_43_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_43_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_43_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_43_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_43_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_43_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_43_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_43_1233 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_124 ();
 sky130_as_sc_hs__decap_16 FILLER_0_43_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_43_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_43_1273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_132 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_148 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_166 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_174 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_187 ();
 sky130_as_sc_hs__decap_4 FILLER_0_43_195 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_201 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_212 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_218 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_222 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_225 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_233 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_252 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_256 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_262 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_279 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_287 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_319 ();
 sky130_as_sc_hs__decap_4 FILLER_0_43_323 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_327 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_335 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_342 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_355 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_375 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_393 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_40 ();
 sky130_as_sc_hs__decap_4 FILLER_0_43_408 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_412 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_428 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_446 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_500 ();
 sky130_as_sc_hs__decap_4 FILLER_0_43_513 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_53 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_550 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_588 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_595 ();
 sky130_as_sc_hs__decap_4 FILLER_0_43_609 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_615 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_629 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_63 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_635 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_639 ();
 sky130_as_sc_hs__decap_4 FILLER_0_43_643 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_669 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_677 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_686 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_690 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_699 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_713 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_72 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_724 ();
 sky130_as_sc_hs__decap_4 FILLER_0_43_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_735 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_739 ();
 sky130_as_sc_hs__decap_4 FILLER_0_43_743 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_759 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_763 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_78 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_804 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_82 ();
 sky130_as_sc_hs__decap_3 FILLER_0_43_824 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_850 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_865 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_890 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_932 ();
 sky130_as_sc_hs__decap_4 FILLER_0_43_96 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_971 ();
 sky130_as_sc_hs__fill_1 FILLER_0_43_981 ();
 sky130_as_sc_hs__fill_2 FILLER_0_43_987 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_10 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_101 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_1034 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_1062 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_1066 ();
 sky130_as_sc_hs__decap_16 FILLER_0_44_1070 ();
 sky130_as_sc_hs__decap_4 FILLER_0_44_1086 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_1090 ();
 sky130_as_sc_hs__decap_16 FILLER_0_44_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_44_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_44_1125 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_113 ();
 sky130_as_sc_hs__decap_4 FILLER_0_44_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_44_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_44_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_44_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_44_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_44_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_44_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_44_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_44_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_44_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_128 ();
 sky130_as_sc_hs__decap_4 FILLER_0_44_146 ();
 sky130_as_sc_hs__fill_1 FILLER_0_44_150 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_153 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_157 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_171 ();
 sky130_as_sc_hs__fill_1 FILLER_0_44_18 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_194 ();
 sky130_as_sc_hs__fill_1 FILLER_0_44_215 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_24 ();
 sky130_as_sc_hs__fill_1 FILLER_0_44_251 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_304 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_319 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_351 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_365 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_392 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_403 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_44_428 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_443 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_451 ();
 sky130_as_sc_hs__fill_1 FILLER_0_44_490 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_511 ();
 sky130_as_sc_hs__decap_4 FILLER_0_44_516 ();
 sky130_as_sc_hs__fill_1 FILLER_0_44_543 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_549 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_554 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_562 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_566 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_585 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_614 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_618 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_622 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_645 ();
 sky130_as_sc_hs__fill_1 FILLER_0_44_661 ();
 sky130_as_sc_hs__fill_1 FILLER_0_44_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_728 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_745 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_765 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_769 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_778 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_804 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_840 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_847 ();
 sky130_as_sc_hs__fill_1 FILLER_0_44_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_44_867 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_888 ();
 sky130_as_sc_hs__decap_3 FILLER_0_44_894 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_902 ();
 sky130_as_sc_hs__fill_1 FILLER_0_44_923 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_946 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_962 ();
 sky130_as_sc_hs__fill_2 FILLER_0_44_973 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_100 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_1014 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_104 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_1052 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_1056 ();
 sky130_as_sc_hs__decap_4 FILLER_0_45_1060 ();
 sky130_as_sc_hs__decap_16 FILLER_0_45_1065 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_108 ();
 sky130_as_sc_hs__decap_16 FILLER_0_45_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_45_1097 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_11 ();
 sky130_as_sc_hs__decap_4 FILLER_0_45_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_45_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_45_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_45_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_45_1169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_117 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_45_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_45_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_45_1209 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_121 ();
 sky130_as_sc_hs__decap_4 FILLER_0_45_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_45_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_45_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_45_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_45_1273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_132 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_138 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_142 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_146 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_150 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_164 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_182 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_194 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_203 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_211 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_222 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_235 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_249 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_256 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_260 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_28 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_290 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_294 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_312 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_318 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_326 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_334 ();
 sky130_as_sc_hs__decap_4 FILLER_0_45_342 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_348 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_361 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_367 ();
 sky130_as_sc_hs__decap_4 FILLER_0_45_373 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_377 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_380 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_384 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_388 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_432 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_439 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_457 ();
 sky130_as_sc_hs__decap_4 FILLER_0_45_466 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_470 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_473 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_487 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_495 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_50 ();
 sky130_as_sc_hs__decap_4 FILLER_0_45_510 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_529 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_566 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_581 ();
 sky130_as_sc_hs__decap_4 FILLER_0_45_585 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_597 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_605 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_650 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_67 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_673 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_684 ();
 sky130_as_sc_hs__decap_4 FILLER_0_45_704 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_75 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_756 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_812 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_84 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_869 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_889 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_895 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_913 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_92 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_929 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_949 ();
 sky130_as_sc_hs__fill_1 FILLER_0_45_958 ();
 sky130_as_sc_hs__fill_2 FILLER_0_45_96 ();
 sky130_as_sc_hs__decap_3 FILLER_0_45_983 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_1023 ();
 sky130_as_sc_hs__fill_1 FILLER_0_46_1035 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_1050 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_1054 ();
 sky130_as_sc_hs__decap_16 FILLER_0_46_1058 ();
 sky130_as_sc_hs__decap_16 FILLER_0_46_1074 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_1090 ();
 sky130_as_sc_hs__decap_16 FILLER_0_46_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_46_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_46_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_46_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_46_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_46_1165 ();
 sky130_as_sc_hs__decap_4 FILLER_0_46_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_46_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_46_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_46_1205 ();
 sky130_as_sc_hs__fill_1 FILLER_0_46_122 ();
 sky130_as_sc_hs__decap_16 FILLER_0_46_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_46_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_46_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_46_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_46_15 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_161 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_166 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_170 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_183 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_187 ();
 sky130_as_sc_hs__fill_1 FILLER_0_46_207 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_213 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_218 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_223 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_232 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_236 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_240 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_248 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_26 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_268 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_29 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_290 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_318 ();
 sky130_as_sc_hs__fill_1 FILLER_0_46_327 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_333 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_337 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_381 ();
 sky130_as_sc_hs__decap_4 FILLER_0_46_392 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_416 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_426 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_443 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_472 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_496 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_516 ();
 sky130_as_sc_hs__decap_4 FILLER_0_46_526 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_533 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_547 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_571 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_579 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_613 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_618 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_634 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_642 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_66 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_669 ();
 sky130_as_sc_hs__fill_1 FILLER_0_46_677 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_683 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_687 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_691 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_695 ();
 sky130_as_sc_hs__fill_1 FILLER_0_46_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_720 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_724 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_728 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_732 ();
 sky130_as_sc_hs__decap_4 FILLER_0_46_74 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_757 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_791 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_80 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_813 ();
 sky130_as_sc_hs__fill_1 FILLER_0_46_820 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_831 ();
 sky130_as_sc_hs__fill_1 FILLER_0_46_867 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_873 ();
 sky130_as_sc_hs__fill_2 FILLER_0_46_925 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_95 ();
 sky130_as_sc_hs__fill_1 FILLER_0_46_965 ();
 sky130_as_sc_hs__fill_1 FILLER_0_46_979 ();
 sky130_as_sc_hs__decap_3 FILLER_0_46_989 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_1002 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_1024 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_1043 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_1047 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_1051 ();
 sky130_as_sc_hs__fill_8 FILLER_0_47_1055 ();
 sky130_as_sc_hs__decap_4 FILLER_0_47_106 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_1063 ();
 sky130_as_sc_hs__decap_16 FILLER_0_47_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_47_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_47_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_47_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_47_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_47_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_47_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_47_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_47_1177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_47_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_47_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_47_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_47_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_47_1249 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_125 ();
 sky130_as_sc_hs__fill_8 FILLER_0_47_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_47_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_136 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_140 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_154 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_159 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_169 ();
 sky130_as_sc_hs__decap_4 FILLER_0_47_190 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_194 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_23 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_238 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_246 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_250 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_262 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_281 ();
 sky130_as_sc_hs__decap_4 FILLER_0_47_303 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_307 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_320 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_346 ();
 sky130_as_sc_hs__decap_4 FILLER_0_47_353 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_357 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_414 ();
 sky130_as_sc_hs__decap_4 FILLER_0_47_442 ();
 sky130_as_sc_hs__decap_4 FILLER_0_47_459 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_463 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_47 ();
 sky130_as_sc_hs__decap_4 FILLER_0_47_474 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_478 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_481 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_485 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_513 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_534 ();
 sky130_as_sc_hs__decap_4 FILLER_0_47_543 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_549 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_569 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_583 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_596 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_613 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_622 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_628 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_649 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_655 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_659 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_666 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_683 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_707 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_715 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_726 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_734 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_76 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_776 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_782 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_839 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_860 ();
 sky130_as_sc_hs__decap_3 FILLER_0_47_883 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_891 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_913 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_945 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_951 ();
 sky130_as_sc_hs__fill_1 FILLER_0_47_962 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_972 ();
 sky130_as_sc_hs__fill_2 FILLER_0_47_99 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_1001 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_1035 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_1046 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_1050 ();
 sky130_as_sc_hs__decap_16 FILLER_0_48_1054 ();
 sky130_as_sc_hs__decap_16 FILLER_0_48_1070 ();
 sky130_as_sc_hs__decap_4 FILLER_0_48_1086 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_1090 ();
 sky130_as_sc_hs__decap_16 FILLER_0_48_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_48_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_48_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_48_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_48_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_48_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_48_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_48_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_48_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_48_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_48_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_48_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_48_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_141 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_172 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_193 ();
 sky130_as_sc_hs__decap_4 FILLER_0_48_207 ();
 sky130_as_sc_hs__decap_4 FILLER_0_48_213 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_22 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_234 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_251 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_257 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_270 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_274 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_278 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_29 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_302 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_326 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_336 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_347 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_351 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_355 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_373 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_378 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_390 ();
 sky130_as_sc_hs__decap_4 FILLER_0_48_400 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_404 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_418 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_426 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_460 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_465 ();
 sky130_as_sc_hs__decap_4 FILLER_0_48_469 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_515 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_54 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_549 ();
 sky130_as_sc_hs__decap_4 FILLER_0_48_555 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_559 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_567 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_572 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_586 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_593 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_605 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_633 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_653 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_677 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_68 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_696 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_706 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_717 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_748 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_76 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_776 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_794 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_807 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_82 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_826 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_851 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_878 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_913 ();
 sky130_as_sc_hs__decap_3 FILLER_0_48_921 ();
 sky130_as_sc_hs__fill_2 FILLER_0_48_954 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_986 ();
 sky130_as_sc_hs__fill_1 FILLER_0_48_99 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_1017 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_1044 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_1048 ();
 sky130_as_sc_hs__fill_8 FILLER_0_49_1052 ();
 sky130_as_sc_hs__decap_4 FILLER_0_49_1060 ();
 sky130_as_sc_hs__decap_16 FILLER_0_49_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_49_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_49_1097 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_111 ();
 sky130_as_sc_hs__decap_4 FILLER_0_49_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_49_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_49_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_49_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_49_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_49_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_49_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_49_1209 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_122 ();
 sky130_as_sc_hs__decap_4 FILLER_0_49_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_49_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_49_1249 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_126 ();
 sky130_as_sc_hs__fill_8 FILLER_0_49_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_49_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_135 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_14 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_140 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_159 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_165 ();
 sky130_as_sc_hs__decap_4 FILLER_0_49_169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_173 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_176 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_180 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_188 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_202 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_214 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_222 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_240 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_246 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_291 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_295 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_299 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_305 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_309 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_323 ();
 sky130_as_sc_hs__decap_4 FILLER_0_49_329 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_333 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_347 ();
 sky130_as_sc_hs__decap_4 FILLER_0_49_372 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_388 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_414 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_428 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_43 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_443 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_464 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_490 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_518 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_525 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_54 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_548 ();
 sky130_as_sc_hs__decap_4 FILLER_0_49_554 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_569 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_595 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_605 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_630 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_636 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_643 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_65 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_688 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_718 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_748 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_75 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_775 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_781 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_798 ();
 sky130_as_sc_hs__decap_4 FILLER_0_49_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_826 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_832 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_838 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_858 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_894 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_897 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_950 ();
 sky130_as_sc_hs__fill_2 FILLER_0_49_966 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_978 ();
 sky130_as_sc_hs__decap_3 FILLER_0_49_98 ();
 sky130_as_sc_hs__fill_1 FILLER_0_49_999 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1181 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1209 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1225 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1241 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_4_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_213 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_229 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_245 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_249 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_253 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_269 ();
 sky130_as_sc_hs__fill_1 FILLER_0_4_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_285 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_301 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_305 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_309 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_325 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_341 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_357 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_375 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_389 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_405 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_409 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_418 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_450 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_454 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_473 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_477 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_485 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_489 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_511 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_515 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_528 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_533 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_537 ();
 sky130_as_sc_hs__fill_8 FILLER_0_4_553 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_574 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_585 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_61 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_616 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_633 ();
 sky130_as_sc_hs__fill_1 FILLER_0_4_637 ();
 sky130_as_sc_hs__fill_1 FILLER_0_4_645 ();
 sky130_as_sc_hs__fill_1 FILLER_0_4_665 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_679 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_683 ();
 sky130_as_sc_hs__fill_1 FILLER_0_4_691 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_724 ();
 sky130_as_sc_hs__fill_8 FILLER_0_4_740 ();
 sky130_as_sc_hs__fill_1 FILLER_0_4_755 ();
 sky130_as_sc_hs__fill_8 FILLER_0_4_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_765 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_769 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_775 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_779 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_789 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_793 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_825 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_833 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_837 ();
 sky130_as_sc_hs__decap_4 FILLER_0_4_841 ();
 sky130_as_sc_hs__fill_1 FILLER_0_4_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_848 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_852 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_861 ();
 sky130_as_sc_hs__fill_1 FILLER_0_4_869 ();
 sky130_as_sc_hs__fill_1 FILLER_0_4_878 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_910 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_914 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_918 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_922 ();
 sky130_as_sc_hs__fill_2 FILLER_0_4_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_929 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_945 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_961 ();
 sky130_as_sc_hs__decap_3 FILLER_0_4_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_4_997 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_10 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_1011 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_1037 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_1041 ();
 sky130_as_sc_hs__decap_16 FILLER_0_50_1045 ();
 sky130_as_sc_hs__decap_16 FILLER_0_50_1061 ();
 sky130_as_sc_hs__fill_8 FILLER_0_50_1077 ();
 sky130_as_sc_hs__decap_4 FILLER_0_50_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_50_1093 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_110 ();
 sky130_as_sc_hs__decap_16 FILLER_0_50_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_50_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_50_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_50_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_50_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_50_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_50_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_50_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_50_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_50_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_50_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_50_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_139 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_146 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_155 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_173 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_195 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_222 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_231 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_248 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_26 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_289 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_50_301 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_305 ();
 sky130_as_sc_hs__decap_4 FILLER_0_50_314 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_318 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_321 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_325 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_334 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_344 ();
 sky130_as_sc_hs__decap_4 FILLER_0_50_357 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_361 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_365 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_383 ();
 sky130_as_sc_hs__decap_4 FILLER_0_50_405 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_411 ();
 sky130_as_sc_hs__decap_4 FILLER_0_50_429 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_433 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_446 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_456 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_475 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_482 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_522 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_530 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_533 ();
 sky130_as_sc_hs__decap_4 FILLER_0_50_541 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_545 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_556 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_568 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_581 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_602 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_606 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_634 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_640 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_654 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_659 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_663 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_670 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_699 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_721 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_794 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_810 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_817 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_842 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_873 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_885 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_890 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_901 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_916 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_923 ();
 sky130_as_sc_hs__decap_3 FILLER_0_50_938 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_945 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_95 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_970 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_981 ();
 sky130_as_sc_hs__fill_1 FILLER_0_50_99 ();
 sky130_as_sc_hs__fill_2 FILLER_0_50_991 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_1007 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_1009 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_1039 ();
 sky130_as_sc_hs__decap_16 FILLER_0_51_1043 ();
 sky130_as_sc_hs__decap_4 FILLER_0_51_1059 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_1063 ();
 sky130_as_sc_hs__decap_16 FILLER_0_51_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_51_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_51_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_51_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_51_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_51_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_51_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_51_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_51_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_51_1193 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_120 ();
 sky130_as_sc_hs__decap_16 FILLER_0_51_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_51_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_51_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_51_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_51_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_51_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_147 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_160 ();
 sky130_as_sc_hs__decap_4 FILLER_0_51_184 ();
 sky130_as_sc_hs__decap_4 FILLER_0_51_190 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_194 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_197 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_206 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_212 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_225 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_285 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_289 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_3 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_30 ();
 sky130_as_sc_hs__decap_4 FILLER_0_51_312 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_316 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_319 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_333 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_362 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_375 ();
 sky130_as_sc_hs__decap_4 FILLER_0_51_385 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_389 ();
 sky130_as_sc_hs__decap_4 FILLER_0_51_393 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_397 ();
 sky130_as_sc_hs__decap_4 FILLER_0_51_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_414 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_423 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_427 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_431 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_445 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_465 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_469 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_48 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_481 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_485 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_531 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_537 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_551 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_591 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_595 ();
 sky130_as_sc_hs__decap_4 FILLER_0_51_599 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_603 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_625 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_63 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_642 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_646 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_654 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_660 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_664 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_668 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_687 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_71 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_712 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_719 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_723 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_733 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_739 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_76 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_781 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_799 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_80 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_818 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_826 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_84 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_841 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_847 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_868 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_914 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_924 ();
 sky130_as_sc_hs__fill_2 FILLER_0_51_93 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_941 ();
 sky130_as_sc_hs__fill_1 FILLER_0_51_946 ();
 sky130_as_sc_hs__decap_3 FILLER_0_51_953 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_101 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_1012 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_1031 ();
 sky130_as_sc_hs__fill_1 FILLER_0_52_1035 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_1037 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_1041 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_1045 ();
 sky130_as_sc_hs__decap_16 FILLER_0_52_1049 ();
 sky130_as_sc_hs__decap_16 FILLER_0_52_1065 ();
 sky130_as_sc_hs__fill_8 FILLER_0_52_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_52_1093 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_110 ();
 sky130_as_sc_hs__decap_16 FILLER_0_52_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_52_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_52_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_52_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_52_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_52_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_52_119 ();
 sky130_as_sc_hs__decap_4 FILLER_0_52_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_52_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_52_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_52_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_52_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_52_1261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_130 ();
 sky130_as_sc_hs__decap_4 FILLER_0_52_14 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_154 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_158 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_168 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_175 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_183 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_20 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_219 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_227 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_232 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_24 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_243 ();
 sky130_as_sc_hs__fill_1 FILLER_0_52_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_264 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_268 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_280 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_289 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_29 ();
 sky130_as_sc_hs__fill_1 FILLER_0_52_297 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_321 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_344 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_351 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_377 ();
 sky130_as_sc_hs__fill_1 FILLER_0_52_389 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_410 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_417 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_42 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_52_438 ();
 sky130_as_sc_hs__fill_1 FILLER_0_52_449 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_455 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_463 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_467 ();
 sky130_as_sc_hs__fill_1 FILLER_0_52_506 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_51 ();
 sky130_as_sc_hs__fill_1 FILLER_0_52_531 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_541 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_56 ();
 sky130_as_sc_hs__fill_1 FILLER_0_52_574 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_585 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_602 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_606 ();
 sky130_as_sc_hs__fill_1 FILLER_0_52_611 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_625 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_642 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_645 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_658 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_692 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_696 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_705 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_724 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_75 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_753 ();
 sky130_as_sc_hs__fill_1 FILLER_0_52_780 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_796 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_841 ();
 sky130_as_sc_hs__fill_1 FILLER_0_52_845 ();
 sky130_as_sc_hs__fill_1 FILLER_0_52_85 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_865 ();
 sky130_as_sc_hs__decap_3 FILLER_0_52_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_52_973 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_1002 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_1022 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_1026 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_1030 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_1034 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_1038 ();
 sky130_as_sc_hs__decap_16 FILLER_0_53_1042 ();
 sky130_as_sc_hs__decap_4 FILLER_0_53_1058 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_53_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_53_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_53_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_53_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_53_1121 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_53_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_53_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_53_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_53_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_53_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_53_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_53_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_53_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_53_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_53_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_53_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_13 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_136 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_140 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_153 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_159 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_165 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_17 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_174 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_235 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_249 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_260 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_281 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_304 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_324 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_335 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_354 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_370 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_391 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_403 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_435 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_449 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_464 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_494 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_502 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_549 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_557 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_569 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_585 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_625 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_657 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_66 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_683 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_694 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_698 ();
 sky130_as_sc_hs__decap_4 FILLER_0_53_7 ();
 sky130_as_sc_hs__decap_3 FILLER_0_53_706 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_748 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_759 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_779 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_78 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_805 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_832 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_836 ();
 sky130_as_sc_hs__decap_4 FILLER_0_53_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_53_856 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_866 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_894 ();
 sky130_as_sc_hs__fill_2 FILLER_0_53_953 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_10 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_1031 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_1035 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_54_1041 ();
 sky130_as_sc_hs__decap_16 FILLER_0_54_1057 ();
 sky130_as_sc_hs__decap_16 FILLER_0_54_1073 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_54_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_54_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_54_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_54_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_54_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_54_1165 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_54_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_54_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_54_1205 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_122 ();
 sky130_as_sc_hs__decap_16 FILLER_0_54_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_54_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_54_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_54_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_133 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_141 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_158 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_189 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_19 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_203 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_235 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_248 ();
 sky130_as_sc_hs__decap_4 FILLER_0_54_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_259 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_263 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_290 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_294 ();
 sky130_as_sc_hs__decap_4 FILLER_0_54_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_318 ();
 sky130_as_sc_hs__decap_4 FILLER_0_54_332 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_336 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_339 ();
 sky130_as_sc_hs__decap_4 FILLER_0_54_351 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_355 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_363 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_377 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_383 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_39 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_392 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_401 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_416 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_443 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_450 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_456 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_462 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_472 ();
 sky130_as_sc_hs__decap_4 FILLER_0_54_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_481 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_484 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_488 ();
 sky130_as_sc_hs__decap_4 FILLER_0_54_49 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_492 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_501 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_517 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_528 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_543 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_55 ();
 sky130_as_sc_hs__decap_4 FILLER_0_54_550 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_554 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_557 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_561 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_565 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_585 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_602 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_624 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_631 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_641 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_649 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_653 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_657 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_678 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_69 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_7 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_734 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_75 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_794 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_825 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_829 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_83 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_833 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_845 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_85 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_90 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_922 ();
 sky130_as_sc_hs__decap_3 FILLER_0_54_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_951 ();
 sky130_as_sc_hs__fill_1 FILLER_0_54_963 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_978 ();
 sky130_as_sc_hs__fill_2 FILLER_0_54_99 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_1022 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_1026 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_1030 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_1034 ();
 sky130_as_sc_hs__decap_16 FILLER_0_55_1038 ();
 sky130_as_sc_hs__fill_8 FILLER_0_55_1054 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_55_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_55_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_55_1097 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_111 ();
 sky130_as_sc_hs__decap_4 FILLER_0_55_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_55_1121 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_55_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_55_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_55_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_55_1177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_55_1193 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_12 ();
 sky130_as_sc_hs__decap_16 FILLER_0_55_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_55_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_55_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_55_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_55_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_55_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_132 ();
 sky130_as_sc_hs__decap_4 FILLER_0_55_136 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_147 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_151 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_155 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_164 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_183 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_207 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_21 ();
 sky130_as_sc_hs__decap_4 FILLER_0_55_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_232 ();
 sky130_as_sc_hs__decap_4 FILLER_0_55_236 ();
 sky130_as_sc_hs__decap_4 FILLER_0_55_242 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_262 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_266 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_277 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_281 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_286 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_292 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_304 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_308 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_327 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_332 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_347 ();
 sky130_as_sc_hs__decap_4 FILLER_0_55_35 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_376 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_384 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_39 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_391 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_398 ();
 sky130_as_sc_hs__decap_4 FILLER_0_55_408 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_412 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_415 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_433 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_437 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_454 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_470 ();
 sky130_as_sc_hs__decap_4 FILLER_0_55_488 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_492 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_495 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_513 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_52 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_526 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_532 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_561 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_575 ();
 sky130_as_sc_hs__decap_4 FILLER_0_55_588 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_606 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_610 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_627 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_638 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_648 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_67 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_677 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_681 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_685 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_701 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_705 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_71 ();
 sky130_as_sc_hs__decap_3 FILLER_0_55_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_729 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_761 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_778 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_8 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_817 ();
 sky130_as_sc_hs__decap_4 FILLER_0_55_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_827 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_864 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_890 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_90 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_910 ();
 sky130_as_sc_hs__fill_1 FILLER_0_55_931 ();
 sky130_as_sc_hs__fill_2 FILLER_0_55_953 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_1026 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_1030 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_1034 ();
 sky130_as_sc_hs__decap_16 FILLER_0_56_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_56_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_56_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_56_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_56_1093 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_110 ();
 sky130_as_sc_hs__decap_16 FILLER_0_56_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_56_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_56_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_56_1149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_116 ();
 sky130_as_sc_hs__decap_16 FILLER_0_56_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_56_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_56_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_56_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_56_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_56_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_56_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_56_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_56_146 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_150 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_158 ();
 sky130_as_sc_hs__decap_4 FILLER_0_56_162 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_188 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_192 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_197 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_226 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_268 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_292 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_299 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_306 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_309 ();
 sky130_as_sc_hs__decap_4 FILLER_0_56_326 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_337 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_34 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_363 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_374 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_40 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_418 ();
 sky130_as_sc_hs__decap_4 FILLER_0_56_442 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_446 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_465 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_477 ();
 sky130_as_sc_hs__decap_4 FILLER_0_56_48 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_500 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_511 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_52 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_529 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_551 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_574 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_608 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_612 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_616 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_664 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_672 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_676 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_695 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_699 ();
 sky130_as_sc_hs__decap_4 FILLER_0_56_70 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_716 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_741 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_754 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_793 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_821 ();
 sky130_as_sc_hs__decap_3 FILLER_0_56_846 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_56_934 ();
 sky130_as_sc_hs__fill_1 FILLER_0_56_979 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_1007 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_1033 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_1037 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_104 ();
 sky130_as_sc_hs__decap_16 FILLER_0_57_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_57_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_57_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_57_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_57_1097 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_11 ();
 sky130_as_sc_hs__decap_4 FILLER_0_57_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_57_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_57_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_57_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_57_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_57_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_57_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_57_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_57_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_57_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_57_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_57_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_57_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_128 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_133 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_152 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_196 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_212 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_247 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_264 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_281 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_29 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_296 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_319 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_335 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_337 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_345 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_355 ();
 sky130_as_sc_hs__decap_4 FILLER_0_57_361 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_368 ();
 sky130_as_sc_hs__decap_4 FILLER_0_57_380 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_384 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_387 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_397 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_401 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_405 ();
 sky130_as_sc_hs__decap_4 FILLER_0_57_417 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_428 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_432 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_444 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_449 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_467 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_481 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_492 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_496 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_500 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_505 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_513 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_52 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_557 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_582 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_586 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_590 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_614 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_627 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_647 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_661 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_668 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_696 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_721 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_727 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_759 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_777 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_798 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_819 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_827 ();
 sky130_as_sc_hs__fill_2 FILLER_0_57_833 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_907 ();
 sky130_as_sc_hs__fill_1 FILLER_0_57_951 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_96 ();
 sky130_as_sc_hs__decap_3 FILLER_0_57_994 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_1007 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_1033 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_1041 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_1045 ();
 sky130_as_sc_hs__decap_16 FILLER_0_58_1049 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_105 ();
 sky130_as_sc_hs__decap_16 FILLER_0_58_1065 ();
 sky130_as_sc_hs__fill_8 FILLER_0_58_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_1089 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_58_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_58_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_58_1125 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_113 ();
 sky130_as_sc_hs__decap_4 FILLER_0_58_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_58_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_58_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_58_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_58_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_58_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_58_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_58_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_58_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_58_1261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_127 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_165 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_174 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_184 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_188 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_192 ();
 sky130_as_sc_hs__decap_4 FILLER_0_58_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_203 ();
 sky130_as_sc_hs__decap_4 FILLER_0_58_217 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_238 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_249 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_277 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_287 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_304 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_344 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_351 ();
 sky130_as_sc_hs__decap_4 FILLER_0_58_357 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_361 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_365 ();
 sky130_as_sc_hs__decap_4 FILLER_0_58_374 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_378 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_389 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_39 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_407 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_437 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_443 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_451 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_463 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_474 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_48 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_482 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_515 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_520 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_538 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_554 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_568 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_598 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_616 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_622 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_645 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_649 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_668 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_672 ();
 sky130_as_sc_hs__decap_4 FILLER_0_58_69 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_697 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_7 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_711 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_722 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_748 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_75 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_780 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_79 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_796 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_802 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_809 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_822 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_854 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_861 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_867 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_869 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_90 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_921 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_938 ();
 sky130_as_sc_hs__fill_2 FILLER_0_58_964 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_971 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_977 ();
 sky130_as_sc_hs__decap_3 FILLER_0_58_981 ();
 sky130_as_sc_hs__fill_1 FILLER_0_58_997 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_10 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_1014 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_1038 ();
 sky130_as_sc_hs__decap_16 FILLER_0_59_1042 ();
 sky130_as_sc_hs__decap_4 FILLER_0_59_1058 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_59_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_59_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_59_1097 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_111 ();
 sky130_as_sc_hs__decap_4 FILLER_0_59_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_59_1121 ();
 sky130_as_sc_hs__decap_4 FILLER_0_59_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_59_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_59_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_59_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_59_1177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_119 ();
 sky130_as_sc_hs__decap_16 FILLER_0_59_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_59_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_59_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_59_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_59_1249 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_126 ();
 sky130_as_sc_hs__fill_8 FILLER_0_59_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_59_1273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_132 ();
 sky130_as_sc_hs__decap_4 FILLER_0_59_148 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_152 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_155 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_159 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_182 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_188 ();
 sky130_as_sc_hs__decap_4 FILLER_0_59_19 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_192 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_196 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_200 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_230 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_234 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_238 ();
 sky130_as_sc_hs__decap_4 FILLER_0_59_242 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_25 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_259 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_263 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_281 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_289 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_294 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_298 ();
 sky130_as_sc_hs__decap_4 FILLER_0_59_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_302 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_306 ();
 sky130_as_sc_hs__decap_4 FILLER_0_59_320 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_327 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_337 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_351 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_425 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_44 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_464 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_473 ();
 sky130_as_sc_hs__decap_4 FILLER_0_59_50 ();
 sky130_as_sc_hs__decap_4 FILLER_0_59_518 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_522 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_541 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_549 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_561 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_615 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_623 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_637 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_660 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_683 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_703 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_707 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_713 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_733 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_770 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_790 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_839 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_851 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_86 ();
 sky130_as_sc_hs__fill_1 FILLER_0_59_915 ();
 sky130_as_sc_hs__decap_3 FILLER_0_59_949 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_958 ();
 sky130_as_sc_hs__fill_2 FILLER_0_59_977 ();
 sky130_as_sc_hs__decap_4 FILLER_0_5_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_5_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_5_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_5_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_5_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_5_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_5_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_5_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_5_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_5_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_225 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_241 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_5_273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_277 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_297 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_3 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_313 ();
 sky130_as_sc_hs__decap_4 FILLER_0_5_329 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_333 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_35 ();
 sky130_as_sc_hs__fill_8 FILLER_0_5_353 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_361 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_374 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_398 ();
 sky130_as_sc_hs__fill_1 FILLER_0_5_437 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_457 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_491 ();
 sky130_as_sc_hs__fill_1 FILLER_0_5_495 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_501 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_5_51 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_526 ();
 sky130_as_sc_hs__fill_8 FILLER_0_5_546 ();
 sky130_as_sc_hs__fill_1 FILLER_0_5_55 ();
 sky130_as_sc_hs__decap_4 FILLER_0_5_554 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_591 ();
 sky130_as_sc_hs__fill_1 FILLER_0_5_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_621 ();
 sky130_as_sc_hs__fill_1 FILLER_0_5_671 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_708 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_733 ();
 sky130_as_sc_hs__fill_1 FILLER_0_5_745 ();
 sky130_as_sc_hs__fill_1 FILLER_0_5_783 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_785 ();
 sky130_as_sc_hs__fill_1 FILLER_0_5_817 ();
 sky130_as_sc_hs__fill_1 FILLER_0_5_822 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_836 ();
 sky130_as_sc_hs__fill_1 FILLER_0_5_868 ();
 sky130_as_sc_hs__fill_1 FILLER_0_5_873 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_89 ();
 sky130_as_sc_hs__fill_1 FILLER_0_5_895 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_905 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_915 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_927 ();
 sky130_as_sc_hs__decap_3 FILLER_0_5_931 ();
 sky130_as_sc_hs__fill_8 FILLER_0_5_942 ();
 sky130_as_sc_hs__fill_2 FILLER_0_5_950 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_5_985 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_10 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_1031 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_1035 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_60_1041 ();
 sky130_as_sc_hs__decap_16 FILLER_0_60_1057 ();
 sky130_as_sc_hs__decap_16 FILLER_0_60_1073 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_60_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_60_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_60_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_60_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_60_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_60_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_60_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_60_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_60_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_60_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_60_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_60_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_60_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_139 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_14 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_156 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_167 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_208 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_221 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_275 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_29 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_295 ();
 sky130_as_sc_hs__decap_4 FILLER_0_60_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_301 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_307 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_317 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_330 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_347 ();
 sky130_as_sc_hs__decap_4 FILLER_0_60_358 ();
 sky130_as_sc_hs__decap_4 FILLER_0_60_370 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_394 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_411 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_417 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_42 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_425 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_451 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_474 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_482 ();
 sky130_as_sc_hs__decap_4 FILLER_0_60_491 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_495 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_498 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_50 ();
 sky130_as_sc_hs__decap_4 FILLER_0_60_511 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_515 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_531 ();
 sky130_as_sc_hs__decap_4 FILLER_0_60_533 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_537 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_544 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_550 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_556 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_563 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_583 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_605 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_624 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_628 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_664 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_698 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_701 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_705 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_732 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_736 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_757 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_761 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_78 ();
 sky130_as_sc_hs__decap_4 FILLER_0_60_794 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_800 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_804 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_808 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_825 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_844 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_850 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_856 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_867 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_873 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_893 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_917 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_923 ();
 sky130_as_sc_hs__fill_2 FILLER_0_60_925 ();
 sky130_as_sc_hs__fill_1 FILLER_0_60_936 ();
 sky130_as_sc_hs__decap_3 FILLER_0_60_99 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_10 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_1026 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_1030 ();
 sky130_as_sc_hs__decap_16 FILLER_0_61_1034 ();
 sky130_as_sc_hs__fill_8 FILLER_0_61_1050 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_1058 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_61_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_61_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_61_1097 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_111 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_61_1121 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_61_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_61_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_61_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_61_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_61_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_61_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_61_1249 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_126 ();
 sky130_as_sc_hs__fill_8 FILLER_0_61_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_1273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_131 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_137 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_14 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_143 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_147 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_156 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_160 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_17 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_180 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_184 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_203 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_21 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_220 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_236 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_248 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_260 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_266 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_281 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_290 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_30 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_321 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_332 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_351 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_393 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_401 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_407 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_420 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_449 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_465 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_471 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_480 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_491 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_496 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_500 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_505 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_519 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_536 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_540 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_55 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_554 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_561 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_568 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_572 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_575 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_579 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_587 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_609 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_627 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_633 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_637 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_652 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_656 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_669 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_673 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_677 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_680 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_686 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_708 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_714 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_718 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_722 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_772 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_795 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_803 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_809 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_81 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_813 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_820 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_846 ();
 sky130_as_sc_hs__decap_4 FILLER_0_61_87 ();
 sky130_as_sc_hs__fill_2 FILLER_0_61_871 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_913 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_941 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_949 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_975 ();
 sky130_as_sc_hs__decap_3 FILLER_0_61_98 ();
 sky130_as_sc_hs__fill_1 FILLER_0_61_983 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_1014 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_1018 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_1022 ();
 sky130_as_sc_hs__fill_8 FILLER_0_62_1026 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_1034 ();
 sky130_as_sc_hs__decap_16 FILLER_0_62_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_62_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_62_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_62_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_62_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_62_1109 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_111 ();
 sky130_as_sc_hs__decap_16 FILLER_0_62_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_62_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_62_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_62_1165 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_62_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_62_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_62_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_62_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_62_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_62_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_62_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_128 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_15 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_166 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_175 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_195 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_210 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_217 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_224 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_235 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_243 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_250 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_253 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_271 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_29 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_292 ();
 sky130_as_sc_hs__decap_4 FILLER_0_62_298 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_304 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_319 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_323 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_347 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_354 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_37 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_389 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_399 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_414 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_440 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_459 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_466 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_477 ();
 sky130_as_sc_hs__decap_4 FILLER_0_62_48 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_491 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_498 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_524 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_552 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_587 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_602 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_640 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_645 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_655 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_681 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_685 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_699 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_739 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_748 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_752 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_769 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_773 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_777 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_783 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_792 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_851 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_874 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_922 ();
 sky130_as_sc_hs__decap_4 FILLER_0_62_94 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_945 ();
 sky130_as_sc_hs__fill_2 FILLER_0_62_978 ();
 sky130_as_sc_hs__fill_1 FILLER_0_62_98 ();
 sky130_as_sc_hs__decap_3 FILLER_0_62_990 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_1003 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_1007 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_1009 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_1013 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_1017 ();
 sky130_as_sc_hs__decap_16 FILLER_0_63_1021 ();
 sky130_as_sc_hs__decap_16 FILLER_0_63_1037 ();
 sky130_as_sc_hs__fill_8 FILLER_0_63_1053 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_63_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_63_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_63_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_63_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_63_1121 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_63_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_63_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_63_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_63_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_63_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_63_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_63_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_63_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_63_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_63_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_63_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_146 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_159 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_164 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_189 ();
 sky130_as_sc_hs__decap_4 FILLER_0_63_197 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_235 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_251 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_257 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_277 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_321 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_334 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_342 ();
 sky130_as_sc_hs__decap_4 FILLER_0_63_352 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_38 ();
 sky130_as_sc_hs__decap_4 FILLER_0_63_381 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_385 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_388 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_393 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_420 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_440 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_470 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_478 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_485 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_49 ();
 sky130_as_sc_hs__decap_4 FILLER_0_63_510 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_516 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_520 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_529 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_541 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_574 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_613 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_622 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_627 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_632 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_64 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_660 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_677 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_681 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_70 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_704 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_708 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_712 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_716 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_722 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_726 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_742 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_762 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_771 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_775 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_795 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_816 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_837 ();
 sky130_as_sc_hs__decap_4 FILLER_0_63_86 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_876 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_897 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_923 ();
 sky130_as_sc_hs__fill_1 FILLER_0_63_932 ();
 sky130_as_sc_hs__fill_2 FILLER_0_63_958 ();
 sky130_as_sc_hs__decap_3 FILLER_0_63_984 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_1010 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1014 ();
 sky130_as_sc_hs__decap_4 FILLER_0_64_1030 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_1034 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1037 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_104 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_64_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_64_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_64_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1205 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_122 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_64_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_64_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_127 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_131 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_135 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_150 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_160 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_177 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_181 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_212 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_220 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_264 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_278 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_287 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_29 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_295 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_304 ();
 sky130_as_sc_hs__decap_4 FILLER_0_64_309 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_313 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_316 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_335 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_373 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_380 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_400 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_421 ();
 sky130_as_sc_hs__decap_4 FILLER_0_64_440 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_444 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_474 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_482 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_487 ();
 sky130_as_sc_hs__decap_4 FILLER_0_64_496 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_502 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_530 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_549 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_574 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_586 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_594 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_603 ();
 sky130_as_sc_hs__decap_4 FILLER_0_64_607 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_61 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_611 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_614 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_685 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_689 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_693 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_727 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_731 ();
 sky130_as_sc_hs__decap_4 FILLER_0_64_74 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_753 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_766 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_796 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_80 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_807 ();
 sky130_as_sc_hs__decap_4 FILLER_0_64_813 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_817 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_833 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_862 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_877 ();
 sky130_as_sc_hs__fill_2 FILLER_0_64_899 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_906 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_915 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_930 ();
 sky130_as_sc_hs__decap_3 FILLER_0_64_96 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_979 ();
 sky130_as_sc_hs__fill_1 FILLER_0_64_986 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_1000 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_1004 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_1009 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_1013 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_1018 ();
 sky130_as_sc_hs__decap_16 FILLER_0_65_1022 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_103 ();
 sky130_as_sc_hs__decap_16 FILLER_0_65_1038 ();
 sky130_as_sc_hs__fill_8 FILLER_0_65_1054 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_65_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_65_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_65_1097 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_110 ();
 sky130_as_sc_hs__decap_4 FILLER_0_65_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_65_1121 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_65_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_65_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_65_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_65_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_65_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_65_1209 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_121 ();
 sky130_as_sc_hs__decap_4 FILLER_0_65_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_65_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_65_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_65_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_65_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_128 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_136 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_166 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_174 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_187 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_19 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_198 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_210 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_216 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_230 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_239 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_245 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_255 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_270 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_276 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_281 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_291 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_297 ();
 sky130_as_sc_hs__decap_4 FILLER_0_65_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_301 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_305 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_328 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_352 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_391 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_397 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_41 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_445 ();
 sky130_as_sc_hs__decap_4 FILLER_0_65_453 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_457 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_48 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_494 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_505 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_550 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_558 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_571 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_617 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_637 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_65 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_657 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_661 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_669 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_681 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_685 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_706 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_710 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_714 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_718 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_722 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_733 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_737 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_783 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_823 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_846 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_852 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_86 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_875 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_895 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_897 ();
 sky130_as_sc_hs__decap_3 FILLER_0_65_910 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_918 ();
 sky130_as_sc_hs__fill_1 FILLER_0_65_951 ();
 sky130_as_sc_hs__fill_2 FILLER_0_65_962 ();
 sky130_as_sc_hs__decap_16 FILLER_0_66_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_66_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_66_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_66_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_66_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_66_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_66_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_66_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_66_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_66_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_66_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_66_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_66_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_66_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_66_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_66_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_66_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_66_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_66_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_66_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_66_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_151 ();
 sky130_as_sc_hs__decap_3 FILLER_0_66_158 ();
 sky130_as_sc_hs__decap_4 FILLER_0_66_163 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_167 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_195 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_197 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_239 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_245 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_251 ();
 sky130_as_sc_hs__decap_3 FILLER_0_66_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_29 ();
 sky130_as_sc_hs__decap_3 FILLER_0_66_305 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_66_321 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_326 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_330 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_339 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_350 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_40 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_419 ();
 sky130_as_sc_hs__decap_3 FILLER_0_66_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_452 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_458 ();
 sky130_as_sc_hs__decap_4 FILLER_0_66_469 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_473 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_482 ();
 sky130_as_sc_hs__decap_3 FILLER_0_66_499 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_517 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_530 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_597 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_632 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_643 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_666 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_696 ();
 sky130_as_sc_hs__decap_3 FILLER_0_66_720 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_73 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_755 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_757 ();
 sky130_as_sc_hs__decap_4 FILLER_0_66_761 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_765 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_772 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_80 ();
 sky130_as_sc_hs__decap_3 FILLER_0_66_804 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_899 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_972 ();
 sky130_as_sc_hs__fill_2 FILLER_0_66_978 ();
 sky130_as_sc_hs__fill_1 FILLER_0_66_997 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_1000 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_1004 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_1009 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_1013 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_1017 ();
 sky130_as_sc_hs__decap_16 FILLER_0_67_1021 ();
 sky130_as_sc_hs__decap_16 FILLER_0_67_1037 ();
 sky130_as_sc_hs__fill_8 FILLER_0_67_1053 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_67_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_67_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_67_1097 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_110 ();
 sky130_as_sc_hs__decap_4 FILLER_0_67_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_67_1121 ();
 sky130_as_sc_hs__decap_4 FILLER_0_67_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_67_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_67_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_67_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_67_1177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_119 ();
 sky130_as_sc_hs__decap_16 FILLER_0_67_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_67_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_67_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_1229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_67_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_67_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_67_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_67_1273 ();
 sky130_as_sc_hs__decap_4 FILLER_0_67_132 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_136 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_144 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_164 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_174 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_189 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_19 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_194 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_214 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_257 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_264 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_294 ();
 sky130_as_sc_hs__decap_4 FILLER_0_67_342 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_348 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_352 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_364 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_372 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_387 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_393 ();
 sky130_as_sc_hs__decap_4 FILLER_0_67_400 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_411 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_422 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_435 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_44 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_447 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_449 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_468 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_479 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_50 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_513 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_528 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_533 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_542 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_559 ();
 sky130_as_sc_hs__decap_4 FILLER_0_67_566 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_570 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_573 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_581 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_591 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_595 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_626 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_644 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_668 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_744 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_755 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_759 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_781 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_812 ();
 sky130_as_sc_hs__decap_4 FILLER_0_67_816 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_822 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_866 ();
 sky130_as_sc_hs__decap_3 FILLER_0_67_870 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_875 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_881 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_907 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_917 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_92 ();
 sky130_as_sc_hs__fill_1 FILLER_0_67_926 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_958 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_98 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_992 ();
 sky130_as_sc_hs__fill_2 FILLER_0_67_996 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_1001 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_1005 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_68_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_68_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_68_1056 ();
 sky130_as_sc_hs__decap_16 FILLER_0_68_1072 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_108 ();
 sky130_as_sc_hs__decap_4 FILLER_0_68_1088 ();
 sky130_as_sc_hs__decap_16 FILLER_0_68_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_68_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_68_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_68_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_68_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_68_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_68_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_68_1197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_12 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_68_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_68_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_68_1237 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_68_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_68_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_134 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_151 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_156 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_160 ();
 sky130_as_sc_hs__decap_4 FILLER_0_68_169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_173 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_176 ();
 sky130_as_sc_hs__decap_4 FILLER_0_68_190 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_215 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_228 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_234 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_244 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_250 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_257 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_26 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_270 ();
 sky130_as_sc_hs__decap_4 FILLER_0_68_279 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_285 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_294 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_306 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_318 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_322 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_336 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_365 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_369 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_37 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_375 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_413 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_426 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_448 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_461 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_475 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_494 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_516 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_530 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_552 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_573 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_586 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_599 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_605 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_642 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_665 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_686 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_699 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_7 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_706 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_710 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_714 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_720 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_724 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_728 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_740 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_744 ();
 sky130_as_sc_hs__decap_3 FILLER_0_68_748 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_771 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_805 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_840 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_844 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_848 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_866 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_874 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_884 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_923 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_925 ();
 sky130_as_sc_hs__fill_1 FILLER_0_68_956 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_978 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_985 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_989 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_99 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_993 ();
 sky130_as_sc_hs__fill_2 FILLER_0_68_997 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_10 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_1007 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_1013 ();
 sky130_as_sc_hs__decap_16 FILLER_0_69_1017 ();
 sky130_as_sc_hs__decap_16 FILLER_0_69_1033 ();
 sky130_as_sc_hs__fill_8 FILLER_0_69_1049 ();
 sky130_as_sc_hs__decap_4 FILLER_0_69_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_69_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_69_1081 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_1097 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_111 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_1118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_69_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_69_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_69_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_69_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_69_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_69_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_69_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_69_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_69_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_69_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_69_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_69_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_142 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_155 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_184 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_212 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_230 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_238 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_242 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_246 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_250 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_254 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_268 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_286 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_292 ();
 sky130_as_sc_hs__decap_4 FILLER_0_69_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_69_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_306 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_320 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_332 ();
 sky130_as_sc_hs__decap_4 FILLER_0_69_337 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_341 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_366 ();
 sky130_as_sc_hs__decap_4 FILLER_0_69_385 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_389 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_402 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_406 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_410 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_414 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_436 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_44 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_449 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_468 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_502 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_510 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_530 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_569 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_575 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_601 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_609 ();
 sky130_as_sc_hs__decap_4 FILLER_0_69_625 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_629 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_637 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_649 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_657 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_665 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_683 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_7 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_713 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_724 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_733 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_754 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_758 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_770 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_804 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_82 ();
 sky130_as_sc_hs__fill_1 FILLER_0_69_846 ();
 sky130_as_sc_hs__decap_3 FILLER_0_69_893 ();
 sky130_as_sc_hs__fill_2 FILLER_0_69_94 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_6_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_213 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_229 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_245 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_249 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_253 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_269 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_285 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_301 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_305 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_309 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_325 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_341 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_357 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_361 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_375 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_391 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_395 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_401 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_405 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_421 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_45 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_452 ();
 sky130_as_sc_hs__fill_8 FILLER_0_6_468 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_481 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_492 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_503 ();
 sky130_as_sc_hs__fill_2 FILLER_0_6_514 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_523 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_531 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_542 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_6_562 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_571 ();
 sky130_as_sc_hs__fill_2 FILLER_0_6_586 ();
 sky130_as_sc_hs__fill_2 FILLER_0_6_603 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_61 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_638 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_664 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_684 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_697 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_706 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_712 ();
 sky130_as_sc_hs__fill_2 FILLER_0_6_761 ();
 sky130_as_sc_hs__fill_2 FILLER_0_6_765 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_769 ();
 sky130_as_sc_hs__decap_4 FILLER_0_6_77 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_809 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_81 ();
 sky130_as_sc_hs__decap_3 FILLER_0_6_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_857 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_867 ();
 sky130_as_sc_hs__fill_1 FILLER_0_6_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_6_874 ();
 sky130_as_sc_hs__fill_2 FILLER_0_6_885 ();
 sky130_as_sc_hs__fill_8 FILLER_0_6_972 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_6_997 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_100 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_1022 ();
 sky130_as_sc_hs__fill_8 FILLER_0_70_1026 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_1034 ();
 sky130_as_sc_hs__decap_16 FILLER_0_70_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_70_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_70_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_70_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_70_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_70_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_70_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_70_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_70_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_70_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_70_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_70_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_70_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_70_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_70_1237 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_124 ();
 sky130_as_sc_hs__decap_4 FILLER_0_70_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_70_1261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_130 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_141 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_158 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_174 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_183 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_203 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_210 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_228 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_25 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_253 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_276 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_287 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_29 ();
 sky130_as_sc_hs__decap_4 FILLER_0_70_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_331 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_335 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_339 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_348 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_360 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_365 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_378 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_386 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_418 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_429 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_435 ();
 sky130_as_sc_hs__decap_4 FILLER_0_70_442 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_446 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_503 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_520 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_538 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_575 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_594 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_602 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_617 ();
 sky130_as_sc_hs__decap_4 FILLER_0_70_621 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_627 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_631 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_635 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_641 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_699 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_7 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_706 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_711 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_728 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_732 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_753 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_778 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_799 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_811 ();
 sky130_as_sc_hs__decap_4 FILLER_0_70_818 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_822 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_825 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_83 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_834 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_840 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_85 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_869 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_881 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_887 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_923 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_925 ();
 sky130_as_sc_hs__fill_1 FILLER_0_70_94 ();
 sky130_as_sc_hs__fill_2 FILLER_0_70_956 ();
 sky130_as_sc_hs__decap_3 FILLER_0_70_977 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_1017 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_1021 ();
 sky130_as_sc_hs__decap_16 FILLER_0_71_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_71_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_71_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_71_1065 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_108 ();
 sky130_as_sc_hs__decap_16 FILLER_0_71_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_71_1097 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_11 ();
 sky130_as_sc_hs__decap_4 FILLER_0_71_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_71_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_71_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_71_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_71_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_71_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_71_1193 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_120 ();
 sky130_as_sc_hs__decap_16 FILLER_0_71_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_71_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_71_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_71_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_71_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_71_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_129 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_134 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_138 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_147 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_15 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_166 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_169 ();
 sky130_as_sc_hs__decap_4 FILLER_0_71_186 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_190 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_193 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_208 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_215 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_231 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_258 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_271 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_276 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_291 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_297 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_313 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_320 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_34 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_342 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_351 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_362 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_383 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_406 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_420 ();
 sky130_as_sc_hs__decap_4 FILLER_0_71_432 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_495 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_502 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_505 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_523 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_551 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_577 ();
 sky130_as_sc_hs__decap_4 FILLER_0_71_606 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_612 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_635 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_64 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_643 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_648 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_658 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_669 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_696 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_718 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_722 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_745 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_749 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_753 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_783 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_849 ();
 sky130_as_sc_hs__decap_3 FILLER_0_71_853 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_87 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_874 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_885 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_913 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_951 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_958 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_965 ();
 sky130_as_sc_hs__fill_1 FILLER_0_71_976 ();
 sky130_as_sc_hs__fill_2 FILLER_0_71_987 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_10 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_1021 ();
 sky130_as_sc_hs__fill_8 FILLER_0_72_1025 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_72_1037 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_104 ();
 sky130_as_sc_hs__decap_16 FILLER_0_72_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_72_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_72_1085 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_1089 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_72_1110 ();
 sky130_as_sc_hs__decap_16 FILLER_0_72_1126 ();
 sky130_as_sc_hs__decap_4 FILLER_0_72_1142 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_1146 ();
 sky130_as_sc_hs__decap_16 FILLER_0_72_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_72_1165 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_72_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_72_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_72_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_72_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_72_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_72_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_72_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_157 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_171 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_189 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_195 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_202 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_222 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_237 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_249 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_25 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_278 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_29 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_291 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_307 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_318 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_322 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_331 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_400 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_418 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_442 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_473 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_49 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_492 ();
 sky130_as_sc_hs__decap_4 FILLER_0_72_505 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_509 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_528 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_533 ();
 sky130_as_sc_hs__decap_4 FILLER_0_72_555 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_559 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_581 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_601 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_609 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_615 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_625 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_643 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_653 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_706 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_71 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_721 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_736 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_778 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_786 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_793 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_800 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_808 ();
 sky130_as_sc_hs__fill_2 FILLER_0_72_847 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_85 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_869 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_938 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_951 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_964 ();
 sky130_as_sc_hs__decap_3 FILLER_0_72_977 ();
 sky130_as_sc_hs__fill_1 FILLER_0_72_98 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_1006 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_102 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_1021 ();
 sky130_as_sc_hs__decap_16 FILLER_0_73_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_73_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_73_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_73_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_73_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_73_1097 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_11 ();
 sky130_as_sc_hs__decap_4 FILLER_0_73_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_73_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_73_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_73_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_73_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_73_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_73_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_73_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_73_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_73_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_73_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_73_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_73_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_128 ();
 sky130_as_sc_hs__fill_1 FILLER_0_73_150 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_156 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_174 ();
 sky130_as_sc_hs__decap_4 FILLER_0_73_183 ();
 sky130_as_sc_hs__fill_1 FILLER_0_73_187 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_210 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_217 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_23 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_240 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_249 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_257 ();
 sky130_as_sc_hs__fill_1 FILLER_0_73_266 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_298 ();
 sky130_as_sc_hs__fill_1 FILLER_0_73_307 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_323 ();
 sky130_as_sc_hs__fill_1 FILLER_0_73_335 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_345 ();
 sky130_as_sc_hs__fill_1 FILLER_0_73_352 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_358 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_362 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_366 ();
 sky130_as_sc_hs__decap_4 FILLER_0_73_385 ();
 sky130_as_sc_hs__fill_1 FILLER_0_73_389 ();
 sky130_as_sc_hs__fill_1 FILLER_0_73_403 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_412 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_42 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_440 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_457 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_489 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_505 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_534 ();
 sky130_as_sc_hs__decap_4 FILLER_0_73_546 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_569 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_625 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_639 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_643 ();
 sky130_as_sc_hs__fill_1 FILLER_0_73_647 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_658 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_670 ();
 sky130_as_sc_hs__fill_1 FILLER_0_73_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_687 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_718 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_722 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_726 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_739 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_743 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_770 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_774 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_778 ();
 sky130_as_sc_hs__fill_1 FILLER_0_73_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_794 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_806 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_821 ();
 sky130_as_sc_hs__decap_4 FILLER_0_73_825 ();
 sky130_as_sc_hs__fill_1 FILLER_0_73_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_832 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_836 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_846 ();
 sky130_as_sc_hs__fill_2 FILLER_0_73_850 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_854 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_86 ();
 sky130_as_sc_hs__fill_1 FILLER_0_73_901 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_922 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_94 ();
 sky130_as_sc_hs__decap_3 FILLER_0_73_949 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_1010 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_1028 ();
 sky130_as_sc_hs__decap_4 FILLER_0_74_1032 ();
 sky130_as_sc_hs__decap_16 FILLER_0_74_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_74_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_74_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_74_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_74_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_74_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_74_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_74_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_74_1149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_115 ();
 sky130_as_sc_hs__decap_16 FILLER_0_74_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_74_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_74_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_74_1205 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_122 ();
 sky130_as_sc_hs__decap_16 FILLER_0_74_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_74_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_74_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_74_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_74_128 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_132 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_135 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_16 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_172 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_187 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_20 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_221 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_237 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_24 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_259 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_284 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_294 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_298 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_307 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_314 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_320 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_333 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_353 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_363 ();
 sky130_as_sc_hs__decap_4 FILLER_0_74_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_371 ();
 sky130_as_sc_hs__decap_4 FILLER_0_74_390 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_396 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_421 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_428 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_43 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_435 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_475 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_490 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_52 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_525 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_551 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_567 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_58 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_585 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_594 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_624 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_661 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_727 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_754 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_757 ();
 sky130_as_sc_hs__decap_3 FILLER_0_74_766 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_77 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_792 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_832 ();
 sky130_as_sc_hs__decap_4 FILLER_0_74_836 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_902 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_908 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_918 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_922 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_940 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_945 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_951 ();
 sky130_as_sc_hs__fill_2 FILLER_0_74_978 ();
 sky130_as_sc_hs__fill_1 FILLER_0_74_996 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_1005 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_1017 ();
 sky130_as_sc_hs__decap_16 FILLER_0_75_1038 ();
 sky130_as_sc_hs__fill_8 FILLER_0_75_1054 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_75_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_75_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_75_1097 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_111 ();
 sky130_as_sc_hs__decap_4 FILLER_0_75_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_75_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_75_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_75_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_75_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_75_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_75_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_75_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_75_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_1229 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_75_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_75_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_75_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_75_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_13 ();
 sky130_as_sc_hs__decap_4 FILLER_0_75_141 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_152 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_200 ();
 sky130_as_sc_hs__decap_4 FILLER_0_75_208 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_212 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_215 ();
 sky130_as_sc_hs__decap_4 FILLER_0_75_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_231 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_235 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_239 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_286 ();
 sky130_as_sc_hs__decap_4 FILLER_0_75_295 ();
 sky130_as_sc_hs__decap_4 FILLER_0_75_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_301 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_305 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_319 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_328 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_332 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_379 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_38 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_383 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_407 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_419 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_427 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_449 ();
 sky130_as_sc_hs__decap_4 FILLER_0_75_461 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_467 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_486 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_505 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_513 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_531 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_561 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_570 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_576 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_587 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_611 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_62 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_638 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_651 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_658 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_669 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_683 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_700 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_727 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_745 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_815 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_83 ();
 sky130_as_sc_hs__fill_1 FILLER_0_75_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_869 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_873 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_894 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_9 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_919 ();
 sky130_as_sc_hs__fill_2 FILLER_0_75_953 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_96 ();
 sky130_as_sc_hs__decap_3 FILLER_0_75_988 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_102 ();
 sky130_as_sc_hs__fill_8 FILLER_0_76_1027 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_1035 ();
 sky130_as_sc_hs__decap_16 FILLER_0_76_1041 ();
 sky130_as_sc_hs__decap_16 FILLER_0_76_1057 ();
 sky130_as_sc_hs__decap_16 FILLER_0_76_1073 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_76_1093 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_110 ();
 sky130_as_sc_hs__decap_16 FILLER_0_76_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_76_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_76_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_76_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_76_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_76_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_76_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_76_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_76_1221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_76_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_76_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_76_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_157 ();
 sky130_as_sc_hs__decap_4 FILLER_0_76_165 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_172 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_186 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_207 ();
 sky130_as_sc_hs__decap_4 FILLER_0_76_214 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_218 ();
 sky130_as_sc_hs__decap_4 FILLER_0_76_226 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_247 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_299 ();
 sky130_as_sc_hs__decap_4 FILLER_0_76_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_307 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_314 ();
 sky130_as_sc_hs__decap_4 FILLER_0_76_321 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_327 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_346 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_362 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_380 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_395 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_42 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_445 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_456 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_46 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_465 ();
 sky130_as_sc_hs__decap_4 FILLER_0_76_520 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_531 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_557 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_594 ();
 sky130_as_sc_hs__decap_4 FILLER_0_76_605 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_609 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_634 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_641 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_661 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_665 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_674 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_678 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_682 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_699 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_7 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_736 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_742 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_80 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_811 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_813 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_827 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_858 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_867 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_877 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_882 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_896 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_901 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_905 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_919 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_923 ();
 sky130_as_sc_hs__fill_1 FILLER_0_76_933 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_947 ();
 sky130_as_sc_hs__fill_2 FILLER_0_76_95 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_966 ();
 sky130_as_sc_hs__decap_3 FILLER_0_76_977 ();
 sky130_as_sc_hs__decap_4 FILLER_0_77_10 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_1005 ();
 sky130_as_sc_hs__decap_4 FILLER_0_77_1009 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_1013 ();
 sky130_as_sc_hs__fill_8 FILLER_0_77_1020 ();
 sky130_as_sc_hs__decap_4 FILLER_0_77_1028 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_1032 ();
 sky130_as_sc_hs__decap_16 FILLER_0_77_1042 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_77_1058 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_77_1065 ();
 sky130_as_sc_hs__fill_8 FILLER_0_77_1081 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_1089 ();
 sky130_as_sc_hs__fill_8 FILLER_0_77_1110 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_1118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_77_1121 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_77_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_77_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_77_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_77_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_77_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_77_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_77_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_1229 ();
 sky130_as_sc_hs__decap_4 FILLER_0_77_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_77_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_77_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_77_1265 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_127 ();
 sky130_as_sc_hs__decap_4 FILLER_0_77_1273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_14 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_140 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_144 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_17 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_180 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_196 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_259 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_26 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_269 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_277 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_285 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_294 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_322 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_334 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_342 ();
 sky130_as_sc_hs__decap_4 FILLER_0_77_364 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_368 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_381 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_40 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_427 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_431 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_435 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_439 ();
 sky130_as_sc_hs__decap_4 FILLER_0_77_483 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_489 ();
 sky130_as_sc_hs__decap_4 FILLER_0_77_498 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_519 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_559 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_565 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_588 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_642 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_669 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_707 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_727 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_762 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_795 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_816 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_828 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_839 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_849 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_857 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_882 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_893 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_916 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_941 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_945 ();
 sky130_as_sc_hs__fill_1 FILLER_0_77_951 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_958 ();
 sky130_as_sc_hs__decap_3 FILLER_0_77_97 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_984 ();
 sky130_as_sc_hs__fill_2 FILLER_0_77_988 ();
 sky130_as_sc_hs__fill_8 FILLER_0_78_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_78_1021 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_1025 ();
 sky130_as_sc_hs__fill_1 FILLER_0_78_1035 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_1052 ();
 sky130_as_sc_hs__decap_16 FILLER_0_78_1056 ();
 sky130_as_sc_hs__fill_1 FILLER_0_78_107 ();
 sky130_as_sc_hs__decap_16 FILLER_0_78_1072 ();
 sky130_as_sc_hs__decap_4 FILLER_0_78_1088 ();
 sky130_as_sc_hs__decap_16 FILLER_0_78_1093 ();
 sky130_as_sc_hs__fill_1 FILLER_0_78_11 ();
 sky130_as_sc_hs__decap_16 FILLER_0_78_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_78_1125 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_113 ();
 sky130_as_sc_hs__decap_4 FILLER_0_78_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_78_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_78_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_78_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_78_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_78_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_78_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_78_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_78_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_78_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_141 ();
 sky130_as_sc_hs__fill_1 FILLER_0_78_150 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_170 ();
 sky130_as_sc_hs__fill_1 FILLER_0_78_195 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_210 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_219 ();
 sky130_as_sc_hs__decap_4 FILLER_0_78_22 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_224 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_228 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_280 ();
 sky130_as_sc_hs__decap_4 FILLER_0_78_287 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_29 ();
 sky130_as_sc_hs__fill_1 FILLER_0_78_291 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_294 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_337 ();
 sky130_as_sc_hs__fill_1 FILLER_0_78_344 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_355 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_377 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_392 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_408 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_418 ();
 sky130_as_sc_hs__fill_1 FILLER_0_78_437 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_443 ();
 sky130_as_sc_hs__decap_4 FILLER_0_78_470 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_506 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_528 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_541 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_567 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_57 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_585 ();
 sky130_as_sc_hs__decap_4 FILLER_0_78_593 ();
 sky130_as_sc_hs__fill_1 FILLER_0_78_597 ();
 sky130_as_sc_hs__decap_4 FILLER_0_78_605 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_61 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_611 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_65 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_658 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_662 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_675 ();
 sky130_as_sc_hs__fill_1 FILLER_0_78_683 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_69 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_698 ();
 sky130_as_sc_hs__fill_1 FILLER_0_78_701 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_741 ();
 sky130_as_sc_hs__decap_4 FILLER_0_78_78 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_804 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_833 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_860 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_864 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_869 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_887 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_89 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_909 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_915 ();
 sky130_as_sc_hs__fill_1 FILLER_0_78_919 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_93 ();
 sky130_as_sc_hs__decap_3 FILLER_0_78_935 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_962 ();
 sky130_as_sc_hs__fill_1 FILLER_0_78_979 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_989 ();
 sky130_as_sc_hs__fill_2 FILLER_0_78_993 ();
 sky130_as_sc_hs__decap_16 FILLER_0_78_997 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_100 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_79_1009 ();
 sky130_as_sc_hs__fill_8 FILLER_0_79_1025 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_1033 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_1037 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_1042 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_1046 ();
 sky130_as_sc_hs__fill_8 FILLER_0_79_1052 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_106 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_1060 ();
 sky130_as_sc_hs__decap_16 FILLER_0_79_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_79_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_79_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_79_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_79_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_79_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_79_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_79_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_79_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_1229 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_79_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_79_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_79_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_128 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_132 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_147 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_161 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_175 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_179 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_223 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_236 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_259 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_27 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_303 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_310 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_324 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_380 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_384 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_398 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_409 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_417 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_43 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_454 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_477 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_483 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_494 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_503 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_510 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_516 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_526 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_530 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_533 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_599 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_608 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_612 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_617 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_621 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_624 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_637 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_644 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_650 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_657 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_666 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_678 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_72 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_727 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_733 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_741 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_78 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_783 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_794 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_823 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_839 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_84 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_852 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_864 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_868 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_872 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_906 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_914 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_918 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_922 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_93 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_933 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_940 ();
 sky130_as_sc_hs__fill_1 FILLER_0_79_944 ();
 sky130_as_sc_hs__decap_3 FILLER_0_79_949 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_79_963 ();
 sky130_as_sc_hs__fill_2 FILLER_0_79_973 ();
 sky130_as_sc_hs__decap_16 FILLER_0_79_977 ();
 sky130_as_sc_hs__fill_8 FILLER_0_79_993 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_1003 ();
 sky130_as_sc_hs__fill_1 FILLER_0_7_1007 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_7_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_225 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_241 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_277 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_297 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_3 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_313 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_329 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_333 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_35 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_353 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_357 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_370 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_383 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_393 ();
 sky130_as_sc_hs__fill_1 FILLER_0_7_415 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_421 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_444 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_449 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_457 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_461 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_474 ();
 sky130_as_sc_hs__fill_1 FILLER_0_7_478 ();
 sky130_as_sc_hs__fill_1 FILLER_0_7_484 ();
 sky130_as_sc_hs__fill_1 FILLER_0_7_503 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_51 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_520 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_533 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_540 ();
 sky130_as_sc_hs__fill_1 FILLER_0_7_544 ();
 sky130_as_sc_hs__fill_1 FILLER_0_7_547 ();
 sky130_as_sc_hs__fill_1 FILLER_0_7_55 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_606 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_613 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_631 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_665 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_669 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_673 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_689 ();
 sky130_as_sc_hs__fill_1 FILLER_0_7_693 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_716 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_726 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_729 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_753 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_767 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_776 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_790 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_820 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_824 ();
 sky130_as_sc_hs__decap_3 FILLER_0_7_837 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_845 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_872 ();
 sky130_as_sc_hs__fill_1 FILLER_0_7_876 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_89 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_890 ();
 sky130_as_sc_hs__fill_2 FILLER_0_7_897 ();
 sky130_as_sc_hs__fill_1 FILLER_0_7_923 ();
 sky130_as_sc_hs__fill_1 FILLER_0_7_942 ();
 sky130_as_sc_hs__decap_4 FILLER_0_7_948 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_963 ();
 sky130_as_sc_hs__decap_16 FILLER_0_7_979 ();
 sky130_as_sc_hs__fill_8 FILLER_0_7_995 ();
 sky130_as_sc_hs__decap_16 FILLER_0_80_1010 ();
 sky130_as_sc_hs__fill_8 FILLER_0_80_1026 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_1034 ();
 sky130_as_sc_hs__decap_16 FILLER_0_80_1075 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_1091 ();
 sky130_as_sc_hs__decap_16 FILLER_0_80_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_80_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_80_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_80_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_80_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_80_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_80_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_80_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_80_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_80_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_80_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_80_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_80_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_131 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_137 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_141 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_189 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_195 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_204 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_23 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_249 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_268 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_278 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_29 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_293 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_80_301 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_305 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_309 ();
 sky130_as_sc_hs__decap_4 FILLER_0_80_321 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_325 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_338 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_344 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_354 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_365 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_373 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_380 ();
 sky130_as_sc_hs__decap_4 FILLER_0_80_389 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_416 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_426 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_435 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_442 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_447 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_48 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_503 ();
 sky130_as_sc_hs__decap_4 FILLER_0_80_512 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_518 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_539 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_554 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_564 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_571 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_581 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_596 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_622 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_641 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_645 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_661 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_678 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_683 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_693 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_720 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_778 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_796 ();
 sky130_as_sc_hs__fill_1 FILLER_0_80_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_853 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_866 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_873 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_882 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_895 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_903 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_907 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_920 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_925 ();
 sky130_as_sc_hs__decap_4 FILLER_0_80_929 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_935 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_939 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_943 ();
 sky130_as_sc_hs__decap_4 FILLER_0_80_947 ();
 sky130_as_sc_hs__decap_16 FILLER_0_80_953 ();
 sky130_as_sc_hs__fill_8 FILLER_0_80_969 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_977 ();
 sky130_as_sc_hs__decap_3 FILLER_0_80_98 ();
 sky130_as_sc_hs__decap_4 FILLER_0_80_981 ();
 sky130_as_sc_hs__fill_2 FILLER_0_80_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_81_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_81_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_81_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_81_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_81_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_81_1273 ();
 sky130_as_sc_hs__decap_4 FILLER_0_81_152 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_158 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_167 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_174 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_178 ();
 sky130_as_sc_hs__decap_4 FILLER_0_81_187 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_191 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_199 ();
 sky130_as_sc_hs__decap_4 FILLER_0_81_208 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_214 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_223 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_230 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_234 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_243 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_252 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_263 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_27 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_292 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_296 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_315 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_329 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_337 ();
 sky130_as_sc_hs__decap_4 FILLER_0_81_345 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_351 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_355 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_359 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_36 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_363 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_367 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_376 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_388 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_393 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_42 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_447 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_460 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_469 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_476 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_480 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_484 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_488 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_492 ();
 sky130_as_sc_hs__decap_4 FILLER_0_81_50 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_510 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_529 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_559 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_566 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_585 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_592 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_596 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_609 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_636 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_65 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_655 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_670 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_713 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_717 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_721 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_733 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_737 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_741 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_790 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_796 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_826 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_83 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_830 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_845 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_849 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_856 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_894 ();
 sky130_as_sc_hs__fill_1 FILLER_0_81_90 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_926 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_930 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_934 ();
 sky130_as_sc_hs__fill_2 FILLER_0_81_950 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_953 ();
 sky130_as_sc_hs__decap_3 FILLER_0_81_96 ();
 sky130_as_sc_hs__decap_16 FILLER_0_81_992 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1000 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1016 ();
 sky130_as_sc_hs__decap_4 FILLER_0_82_1032 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_82_107 ();
 sky130_as_sc_hs__decap_4 FILLER_0_82_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_82_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_82_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1221 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_82_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_134 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_153 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_181 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_188 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_203 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_223 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_228 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_259 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_266 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_285 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_289 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_29 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_318 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_332 ();
 sky130_as_sc_hs__decap_4 FILLER_0_82_341 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_345 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_35 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_363 ();
 sky130_as_sc_hs__decap_4 FILLER_0_82_375 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_379 ();
 sky130_as_sc_hs__decap_4 FILLER_0_82_395 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_401 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_410 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_419 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_421 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_425 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_433 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_457 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_467 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_474 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_486 ();
 sky130_as_sc_hs__decap_4 FILLER_0_82_501 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_507 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_524 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_530 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_54 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_543 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_567 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_598 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_60 ();
 sky130_as_sc_hs__decap_4 FILLER_0_82_611 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_617 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_623 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_632 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_636 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_643 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_645 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_701 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_705 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_709 ();
 sky130_as_sc_hs__decap_4 FILLER_0_82_71 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_713 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_717 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_721 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_729 ();
 sky130_as_sc_hs__decap_4 FILLER_0_82_733 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_737 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_749 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_787 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_817 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_82 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_826 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_837 ();
 sky130_as_sc_hs__fill_1 FILLER_0_82_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_866 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_903 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_907 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_911 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_918 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_922 ();
 sky130_as_sc_hs__fill_2 FILLER_0_82_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_929 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_945 ();
 sky130_as_sc_hs__decap_16 FILLER_0_82_961 ();
 sky130_as_sc_hs__decap_3 FILLER_0_82_977 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_83_1009 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_1025 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_1042 ();
 sky130_as_sc_hs__fill_8 FILLER_0_83_1050 ();
 sky130_as_sc_hs__decap_4 FILLER_0_83_1058 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_83_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_83_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_83_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_83_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_83_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_83_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_83_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_83_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_83_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_83_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_83_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_83_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_83_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_83_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_83_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_83_1273 ();
 sky130_as_sc_hs__decap_4 FILLER_0_83_137 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_164 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_186 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_23 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_230 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_246 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_250 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_259 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_263 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_272 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_278 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_281 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_305 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_310 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_319 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_372 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_38 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_389 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_412 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_423 ();
 sky130_as_sc_hs__decap_4 FILLER_0_83_436 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_440 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_447 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_454 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_458 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_462 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_476 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_483 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_499 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_513 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_53 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_549 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_559 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_566 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_576 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_584 ();
 sky130_as_sc_hs__decap_4 FILLER_0_83_590 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_594 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_615 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_617 ();
 sky130_as_sc_hs__decap_4 FILLER_0_83_628 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_649 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_653 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_711 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_715 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_724 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_781 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_798 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_836 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_846 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_850 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_854 ();
 sky130_as_sc_hs__decap_3 FILLER_0_83_877 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_890 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_894 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_83_909 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_913 ();
 sky130_as_sc_hs__fill_8 FILLER_0_83_953 ();
 sky130_as_sc_hs__fill_1 FILLER_0_83_961 ();
 sky130_as_sc_hs__decap_16 FILLER_0_83_981 ();
 sky130_as_sc_hs__fill_8 FILLER_0_83_997 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_84_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_1056 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_1072 ();
 sky130_as_sc_hs__decap_4 FILLER_0_84_1088 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_1093 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_110 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_84_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_84_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_84_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_1257 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_126 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_131 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_151 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_167 ();
 sky130_as_sc_hs__decap_4 FILLER_0_84_179 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_183 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_207 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_221 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_233 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_25 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_288 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_304 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_315 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_327 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_333 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_339 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_360 ();
 sky130_as_sc_hs__decap_4 FILLER_0_84_370 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_376 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_380 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_394 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_41 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_419 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_421 ();
 sky130_as_sc_hs__decap_4 FILLER_0_84_437 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_453 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_471 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_493 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_50 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_522 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_528 ();
 sky130_as_sc_hs__decap_4 FILLER_0_84_533 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_537 ();
 sky130_as_sc_hs__decap_4 FILLER_0_84_544 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_548 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_575 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_587 ();
 sky130_as_sc_hs__decap_4 FILLER_0_84_594 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_598 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_611 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_623 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_627 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_63 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_643 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_659 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_663 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_672 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_69 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_697 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_713 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_730 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_734 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_738 ();
 sky130_as_sc_hs__decap_4 FILLER_0_84_742 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_748 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_776 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_790 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_796 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_809 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_82 ();
 sky130_as_sc_hs__fill_1 FILLER_0_84_856 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_865 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_885 ();
 sky130_as_sc_hs__decap_3 FILLER_0_84_90 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_922 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_930 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_946 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_962 ();
 sky130_as_sc_hs__fill_2 FILLER_0_84_978 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_84_997 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_85_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_85_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_85_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1177 ();
 sky130_as_sc_hs__decap_4 FILLER_0_85_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_85_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1233 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_124 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_85_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_85_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_128 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_150 ();
 sky130_as_sc_hs__decap_4 FILLER_0_85_156 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_160 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_186 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_203 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_212 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_22 ();
 sky130_as_sc_hs__decap_4 FILLER_0_85_230 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_246 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_26 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_267 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_281 ();
 sky130_as_sc_hs__decap_4 FILLER_0_85_290 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_294 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_297 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_30 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_314 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_350 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_357 ();
 sky130_as_sc_hs__decap_4 FILLER_0_85_373 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_415 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_419 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_423 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_431 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_44 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_442 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_454 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_475 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_479 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_488 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_494 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_503 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_85_509 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_513 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_521 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_531 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_543 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_550 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_592 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_596 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_600 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_608 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_62 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_626 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_644 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_656 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_660 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_669 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_678 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_682 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_686 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_703 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_715 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_726 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_733 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_741 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_773 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_778 ();
 sky130_as_sc_hs__fill_1 FILLER_0_85_78 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_803 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_807 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_811 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_815 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_832 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_854 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_890 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_894 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_897 ();
 sky130_as_sc_hs__decap_4 FILLER_0_85_905 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_909 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_927 ();
 sky130_as_sc_hs__decap_4 FILLER_0_85_948 ();
 sky130_as_sc_hs__fill_8 FILLER_0_85_953 ();
 sky130_as_sc_hs__fill_2 FILLER_0_85_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_85_981 ();
 sky130_as_sc_hs__decap_3 FILLER_0_85_99 ();
 sky130_as_sc_hs__fill_8 FILLER_0_85_997 ();
 sky130_as_sc_hs__fill_1 FILLER_0_86_100 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1013 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_1029 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_1034 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_86_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_86_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_86_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1205 ();
 sky130_as_sc_hs__fill_1 FILLER_0_86_121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_86_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_1261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_132 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_166 ();
 sky130_as_sc_hs__decap_4 FILLER_0_86_190 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_207 ();
 sky130_as_sc_hs__fill_1 FILLER_0_86_21 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_236 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_249 ();
 sky130_as_sc_hs__decap_4 FILLER_0_86_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_269 ();
 sky130_as_sc_hs__fill_1 FILLER_0_86_27 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_319 ();
 sky130_as_sc_hs__fill_1 FILLER_0_86_326 ();
 sky130_as_sc_hs__decap_4 FILLER_0_86_332 ();
 sky130_as_sc_hs__decap_4 FILLER_0_86_338 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_365 ();
 sky130_as_sc_hs__fill_1 FILLER_0_86_373 ();
 sky130_as_sc_hs__fill_1 FILLER_0_86_379 ();
 sky130_as_sc_hs__fill_1 FILLER_0_86_385 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_391 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_396 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_400 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_417 ();
 sky130_as_sc_hs__fill_1 FILLER_0_86_42 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_426 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_430 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_443 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_455 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_467 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_472 ();
 sky130_as_sc_hs__decap_4 FILLER_0_86_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_488 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_504 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_517 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_537 ();
 sky130_as_sc_hs__fill_1 FILLER_0_86_563 ();
 sky130_as_sc_hs__fill_1 FILLER_0_86_58 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_598 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_649 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_667 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_674 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_678 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_686 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_69 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_690 ();
 sky130_as_sc_hs__fill_1 FILLER_0_86_694 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_714 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_718 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_723 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_727 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_731 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_735 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_739 ();
 sky130_as_sc_hs__fill_1 FILLER_0_86_755 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_767 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_81 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_828 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_85 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_865 ();
 sky130_as_sc_hs__fill_2 FILLER_0_86_869 ();
 sky130_as_sc_hs__fill_8 FILLER_0_86_892 ();
 sky130_as_sc_hs__decap_4 FILLER_0_86_900 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_904 ();
 sky130_as_sc_hs__decap_4 FILLER_0_86_917 ();
 sky130_as_sc_hs__decap_3 FILLER_0_86_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_86_997 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_100 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_1005 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_1032 ();
 sky130_as_sc_hs__fill_8 FILLER_0_87_1050 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_1058 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_1062 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_1097 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_110 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_1177 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_1229 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_87_1265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_127 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_147 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_154 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_159 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_179 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_18 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_184 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_203 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_215 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_220 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_225 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_237 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_243 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_267 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_277 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_281 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_292 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_296 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_314 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_337 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_346 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_367 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_371 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_398 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_416 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_42 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_422 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_432 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_459 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_487 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_49 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_505 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_53 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_532 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_547 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_551 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_558 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_57 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_570 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_574 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_606 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_612 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_62 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_622 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_630 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_651 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_657 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_671 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_692 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_71 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_711 ();
 sky130_as_sc_hs__fill_1 FILLER_0_87_760 ();
 sky130_as_sc_hs__decap_3 FILLER_0_87_794 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_816 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_851 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_863 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_875 ();
 sky130_as_sc_hs__decap_4 FILLER_0_87_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_901 ();
 sky130_as_sc_hs__fill_8 FILLER_0_87_923 ();
 sky130_as_sc_hs__fill_2 FILLER_0_87_931 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_87_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_88_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_88_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_88_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_1145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_88_1149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_1153 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_1174 ();
 sky130_as_sc_hs__fill_8 FILLER_0_88_1190 ();
 sky130_as_sc_hs__decap_4 FILLER_0_88_1198 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_1202 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_88_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_132 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_138 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_141 ();
 sky130_as_sc_hs__decap_4 FILLER_0_88_160 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_164 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_167 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_171 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_195 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_220 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_224 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_245 ();
 sky130_as_sc_hs__decap_4 FILLER_0_88_253 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_257 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_270 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_286 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_293 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_300 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_304 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_314 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_323 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_333 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_337 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_35 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_351 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_373 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_386 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_391 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_421 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_43 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_444 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_473 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_482 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_487 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_504 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_531 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_537 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_541 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_550 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_557 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_571 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_575 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_587 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_594 ();
 sky130_as_sc_hs__decap_4 FILLER_0_88_605 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_609 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_622 ();
 sky130_as_sc_hs__decap_4 FILLER_0_88_626 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_630 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_633 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_637 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_64 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_643 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_654 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_658 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_672 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_678 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_682 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_699 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_70 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_730 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_734 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_738 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_742 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_746 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_76 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_80 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_800 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_804 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_832 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_862 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_882 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_90 ();
 sky130_as_sc_hs__decap_4 FILLER_0_88_919 ();
 sky130_as_sc_hs__fill_1 FILLER_0_88_923 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_94 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_88_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_88_977 ();
 sky130_as_sc_hs__fill_2 FILLER_0_88_98 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_88_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_1004 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_89_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_89_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1121 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_1169 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_117 ();
 sky130_as_sc_hs__decap_3 FILLER_0_89_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_89_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_89_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_89_169 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_17 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_198 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_21 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_231 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_24 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_281 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_308 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_327 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_337 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_346 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_350 ();
 sky130_as_sc_hs__decap_3 FILLER_0_89_379 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_390 ();
 sky130_as_sc_hs__decap_3 FILLER_0_89_398 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_405 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_416 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_435 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_44 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_447 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_453 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_457 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_476 ();
 sky130_as_sc_hs__decap_3 FILLER_0_89_491 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_505 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_509 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_517 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_615 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_644 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_655 ();
 sky130_as_sc_hs__decap_3 FILLER_0_89_682 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_690 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_702 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_706 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_710 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_714 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_726 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_733 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_761 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_765 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_769 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_79 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_808 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_812 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_816 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_821 ();
 sky130_as_sc_hs__decap_3 FILLER_0_89_837 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_846 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_856 ();
 sky130_as_sc_hs__fill_8 FILLER_0_89_865 ();
 sky130_as_sc_hs__fill_2 FILLER_0_89_873 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_880 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_889 ();
 sky130_as_sc_hs__decap_3 FILLER_0_89_893 ();
 sky130_as_sc_hs__fill_8 FILLER_0_89_897 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_90 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_905 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_909 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_920 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_936 ();
 sky130_as_sc_hs__fill_1 FILLER_0_89_94 ();
 sky130_as_sc_hs__fill_8 FILLER_0_89_953 ();
 sky130_as_sc_hs__decap_4 FILLER_0_89_961 ();
 sky130_as_sc_hs__decap_16 FILLER_0_89_988 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_101 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1013 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_1029 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_1033 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_1261 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_133 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_141 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_157 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_189 ();
 sky130_as_sc_hs__fill_8 FILLER_0_8_19 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_197 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_213 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_229 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_245 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_249 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_253 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_269 ();
 sky130_as_sc_hs__fill_1 FILLER_0_8_27 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_285 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_29 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_3 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_301 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_305 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_309 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_325 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_341 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_357 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_361 ();
 sky130_as_sc_hs__fill_1 FILLER_0_8_385 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_396 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_406 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_429 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_433 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_45 ();
 sky130_as_sc_hs__fill_1 FILLER_0_8_450 ();
 sky130_as_sc_hs__fill_1 FILLER_0_8_475 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_497 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_528 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_533 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_554 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_577 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_61 ();
 sky130_as_sc_hs__fill_1 FILLER_0_8_639 ();
 sky130_as_sc_hs__fill_1 FILLER_0_8_660 ();
 sky130_as_sc_hs__fill_1 FILLER_0_8_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_711 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_715 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_719 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_745 ();
 sky130_as_sc_hs__decap_4 FILLER_0_8_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_776 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_794 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_81 ();
 sky130_as_sc_hs__fill_1 FILLER_0_8_813 ();
 sky130_as_sc_hs__fill_1 FILLER_0_8_827 ();
 sky130_as_sc_hs__fill_1 FILLER_0_8_848 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_85 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_853 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_896 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_912 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_919 ();
 sky130_as_sc_hs__fill_1 FILLER_0_8_923 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_925 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_929 ();
 sky130_as_sc_hs__fill_2 FILLER_0_8_933 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_937 ();
 sky130_as_sc_hs__fill_8 FILLER_0_8_969 ();
 sky130_as_sc_hs__decap_3 FILLER_0_8_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_8_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_1013 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_1037 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_1054 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_1058 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_1074 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_109 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_1090 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_1149 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_115 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_1181 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_119 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_127 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_133 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_137 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_147 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_156 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_179 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_187 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_192 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_21 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_212 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_216 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_220 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_234 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_243 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_250 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_253 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_263 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_274 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_278 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_286 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_296 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_303 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_314 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_318 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_321 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_336 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_344 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_355 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_365 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_371 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_375 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_421 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_427 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_442 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_448 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_461 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_477 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_487 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_521 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_529 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_533 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_547 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_55 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_551 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_574 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_584 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_589 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_600 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_605 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_619 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_623 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_634 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_638 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_649 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_654 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_658 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_738 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_742 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_746 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_754 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_761 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_765 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_769 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_78 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_794 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_798 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_806 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_810 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_813 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_817 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_825 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_833 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_837 ();
 sky130_as_sc_hs__decap_3 FILLER_0_90_85 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_852 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_864 ();
 sky130_as_sc_hs__decap_4 FILLER_0_90_874 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_878 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_894 ();
 sky130_as_sc_hs__fill_2 FILLER_0_90_9 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_929 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_964 ();
 sky130_as_sc_hs__fill_1 FILLER_0_90_98 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_981 ();
 sky130_as_sc_hs__decap_16 FILLER_0_90_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_1005 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_1009 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_1013 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_1033 ();
 sky130_as_sc_hs__fill_8 FILLER_0_91_1049 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_1103 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_1119 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_1121 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_1177 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_119 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_91_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_1273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_132 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_136 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_155 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_166 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_174 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_190 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_206 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_215 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_223 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_230 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_236 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_255 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_262 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_278 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_291 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_297 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_306 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_313 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_331 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_337 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_367 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_375 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_389 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_397 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_405 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_409 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_425 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_432 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_439 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_45 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_464 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_476 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_503 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_510 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_518 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_522 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_526 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_530 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_539 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_549 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_553 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_556 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_569 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_574 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_594 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_613 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_617 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_629 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_637 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_667 ();
 sky130_as_sc_hs__decap_4 FILLER_0_91_67 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_671 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_673 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_677 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_681 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_690 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_694 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_700 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_706 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_71 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_710 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_726 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_74 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_749 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_753 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_778 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_78 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_797 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_801 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_822 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_846 ();
 sky130_as_sc_hs__fill_1 FILLER_0_91_895 ();
 sky130_as_sc_hs__decap_3 FILLER_0_91_92 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_926 ();
 sky130_as_sc_hs__fill_8 FILLER_0_91_942 ();
 sky130_as_sc_hs__fill_2 FILLER_0_91_950 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_969 ();
 sky130_as_sc_hs__decap_16 FILLER_0_91_985 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1000 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1016 ();
 sky130_as_sc_hs__decap_4 FILLER_0_92_1032 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1037 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_104 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_92_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_92_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_92_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_92_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1165 ();
 sky130_as_sc_hs__decap_4 FILLER_0_92_1181 ();
 sky130_as_sc_hs__fill_1 FILLER_0_92_1203 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_92_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_92_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_136 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_92_153 ();
 sky130_as_sc_hs__decap_3 FILLER_0_92_176 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_92_244 ();
 sky130_as_sc_hs__fill_1 FILLER_0_92_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_289 ();
 sky130_as_sc_hs__decap_4 FILLER_0_92_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_339 ();
 sky130_as_sc_hs__decap_3 FILLER_0_92_351 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_365 ();
 sky130_as_sc_hs__fill_1 FILLER_0_92_37 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_380 ();
 sky130_as_sc_hs__decap_3 FILLER_0_92_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_406 ();
 sky130_as_sc_hs__fill_1 FILLER_0_92_445 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_460 ();
 sky130_as_sc_hs__fill_1 FILLER_0_92_464 ();
 sky130_as_sc_hs__fill_1 FILLER_0_92_475 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_485 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_513 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_53 ();
 sky130_as_sc_hs__decap_3 FILLER_0_92_533 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_541 ();
 sky130_as_sc_hs__decap_4 FILLER_0_92_559 ();
 sky130_as_sc_hs__fill_1 FILLER_0_92_563 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_566 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_640 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_677 ();
 sky130_as_sc_hs__fill_1 FILLER_0_92_681 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_692 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_696 ();
 sky130_as_sc_hs__fill_1 FILLER_0_92_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_717 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_721 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_733 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_741 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_745 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_749 ();
 sky130_as_sc_hs__decap_3 FILLER_0_92_753 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_776 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_784 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_80 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_810 ();
 sky130_as_sc_hs__fill_1 FILLER_0_92_85 ();
 sky130_as_sc_hs__decap_3 FILLER_0_92_852 ();
 sky130_as_sc_hs__decap_3 FILLER_0_92_865 ();
 sky130_as_sc_hs__fill_8 FILLER_0_92_869 ();
 sky130_as_sc_hs__fill_1 FILLER_0_92_877 ();
 sky130_as_sc_hs__fill_8 FILLER_0_92_893 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_906 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_91 ();
 sky130_as_sc_hs__decap_4 FILLER_0_92_920 ();
 sky130_as_sc_hs__fill_8 FILLER_0_92_925 ();
 sky130_as_sc_hs__decap_3 FILLER_0_92_933 ();
 sky130_as_sc_hs__fill_2 FILLER_0_92_95 ();
 sky130_as_sc_hs__decap_16 FILLER_0_92_955 ();
 sky130_as_sc_hs__fill_8 FILLER_0_92_971 ();
 sky130_as_sc_hs__fill_1 FILLER_0_92_979 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_1007 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_1009 ();
 sky130_as_sc_hs__fill_8 FILLER_0_93_1025 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_1033 ();
 sky130_as_sc_hs__decap_4 FILLER_0_93_1059 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_1063 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_1065 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_107 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_93_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_93_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_1177 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_118 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_93_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_93_1265 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_127 ();
 sky130_as_sc_hs__decap_4 FILLER_0_93_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_139 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_149 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_154 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_179 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_195 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_199 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_208 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_223 ();
 sky130_as_sc_hs__decap_4 FILLER_0_93_230 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_234 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_252 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_262 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_271 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_276 ();
 sky130_as_sc_hs__decap_4 FILLER_0_93_281 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_285 ();
 sky130_as_sc_hs__decap_4 FILLER_0_93_298 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_313 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_317 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_337 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_355 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_363 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_387 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_417 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_42 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_428 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_447 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_449 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_460 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_491 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_505 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_538 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_544 ();
 sky130_as_sc_hs__decap_4 FILLER_0_93_553 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_557 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_57 ();
 sky130_as_sc_hs__decap_4 FILLER_0_93_576 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_580 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_583 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_602 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_613 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_627 ();
 sky130_as_sc_hs__decap_4 FILLER_0_93_635 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_667 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_673 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_689 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_698 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_7 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_707 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_711 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_727 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_750 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_754 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_758 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_762 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_766 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_770 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_774 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_778 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_782 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_789 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_793 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_797 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_801 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_815 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_819 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_838 ();
 sky130_as_sc_hs__fill_8 FILLER_0_93_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_849 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_861 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_877 ();
 sky130_as_sc_hs__fill_8 FILLER_0_93_886 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_894 ();
 sky130_as_sc_hs__decap_4 FILLER_0_93_897 ();
 sky130_as_sc_hs__fill_1 FILLER_0_93_901 ();
 sky130_as_sc_hs__fill_2 FILLER_0_93_907 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_932 ();
 sky130_as_sc_hs__decap_4 FILLER_0_93_948 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_953 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_975 ();
 sky130_as_sc_hs__decap_3 FILLER_0_93_99 ();
 sky130_as_sc_hs__decap_16 FILLER_0_93_991 ();
 sky130_as_sc_hs__fill_8 FILLER_0_94_1003 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_1011 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_1053 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_1069 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_1085 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_1089 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_1109 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_111 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_1197 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_120 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_1257 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_126 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_1261 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_157 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_162 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_166 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_185 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_19 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_208 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_213 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_227 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_231 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_240 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_244 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_258 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_266 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_277 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_296 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_320 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_334 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_338 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_341 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_350 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_356 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_360 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_375 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_389 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_393 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_405 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_425 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_43 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_474 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_477 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_483 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_506 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_517 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_524 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_528 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_533 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_537 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_540 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_549 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_567 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_574 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_585 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_59 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_594 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_598 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_627 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_66 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_664 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_668 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_672 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_70 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_709 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_726 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_730 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_743 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_747 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_751 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_755 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_799 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_811 ();
 sky130_as_sc_hs__fill_8 FILLER_0_94_813 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_853 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_867 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_874 ();
 sky130_as_sc_hs__fill_8 FILLER_0_94_915 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_92 ();
 sky130_as_sc_hs__fill_1 FILLER_0_94_923 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_94_957 ();
 sky130_as_sc_hs__fill_2 FILLER_0_94_97 ();
 sky130_as_sc_hs__decap_4 FILLER_0_94_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_977 ();
 sky130_as_sc_hs__decap_3 FILLER_0_94_981 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_1001 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_1005 ();
 sky130_as_sc_hs__fill_8 FILLER_0_95_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_1017 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_1021 ();
 sky130_as_sc_hs__decap_16 FILLER_0_95_1043 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_1059 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_1063 ();
 sky130_as_sc_hs__decap_16 FILLER_0_95_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_95_1081 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_1097 ();
 sky130_as_sc_hs__decap_16 FILLER_0_95_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_95_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_95_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_1173 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_1177 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_1181 ();
 sky130_as_sc_hs__decap_16 FILLER_0_95_1201 ();
 sky130_as_sc_hs__fill_8 FILLER_0_95_1217 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_95_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_95_1249 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_125 ();
 sky130_as_sc_hs__fill_8 FILLER_0_95_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_1273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_131 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_139 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_160 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_167 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_169 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_193 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_21 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_252 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_279 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_291 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_299 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_318 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_335 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_337 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_353 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_364 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_379 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_39 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_390 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_398 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_426 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_43 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_440 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_454 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_474 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_500 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_510 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_525 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_550 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_556 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_566 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_590 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_594 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_662 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_666 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_686 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_690 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_694 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_698 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_710 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_714 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_73 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_772 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_776 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_785 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_805 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_82 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_836 ();
 sky130_as_sc_hs__fill_8 FILLER_0_95_841 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_849 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_856 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_863 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_88 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_890 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_894 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_901 ();
 sky130_as_sc_hs__fill_8 FILLER_0_95_908 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_916 ();
 sky130_as_sc_hs__decap_3 FILLER_0_95_920 ();
 sky130_as_sc_hs__fill_8 FILLER_0_95_942 ();
 sky130_as_sc_hs__fill_2 FILLER_0_95_950 ();
 sky130_as_sc_hs__decap_4 FILLER_0_95_953 ();
 sky130_as_sc_hs__fill_1 FILLER_0_95_957 ();
 sky130_as_sc_hs__decap_16 FILLER_0_95_977 ();
 sky130_as_sc_hs__fill_8 FILLER_0_95_993 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_1001 ();
 sky130_as_sc_hs__fill_8 FILLER_0_96_1025 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_1033 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_1043 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_1059 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_1075 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_1091 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_1093 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_110 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_1125 ();
 sky130_as_sc_hs__decap_4 FILLER_0_96_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_96_1197 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_96_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_1257 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_1261 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_138 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_146 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_152 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_170 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_187 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_209 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_213 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_222 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_228 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_242 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_248 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_304 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_309 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_322 ();
 sky130_as_sc_hs__decap_4 FILLER_0_96_331 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_335 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_338 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_34 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_342 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_346 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_350 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_370 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_419 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_425 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_442 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_455 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_470 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_501 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_505 ();
 sky130_as_sc_hs__decap_4 FILLER_0_96_517 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_521 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_567 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_589 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_60 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_602 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_615 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_640 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_650 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_662 ();
 sky130_as_sc_hs__decap_4 FILLER_0_96_666 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_688 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_699 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_705 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_709 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_717 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_727 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_755 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_757 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_761 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_765 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_769 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_773 ();
 sky130_as_sc_hs__decap_4 FILLER_0_96_777 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_781 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_805 ();
 sky130_as_sc_hs__fill_8 FILLER_0_96_813 ();
 sky130_as_sc_hs__decap_4 FILLER_0_96_821 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_825 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_847 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_861 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_96_884 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_888 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_894 ();
 sky130_as_sc_hs__fill_1 FILLER_0_96_902 ();
 sky130_as_sc_hs__fill_8 FILLER_0_96_913 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_96_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_96_977 ();
 sky130_as_sc_hs__decap_16 FILLER_0_96_981 ();
 sky130_as_sc_hs__decap_4 FILLER_0_96_997 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_1002 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_1006 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_1025 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_104 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_1065 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_108 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_1081 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_1115 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_1119 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_1229 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_123 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_97_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_1273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_131 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_137 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_143 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_147 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_166 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_180 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_184 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_188 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_202 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_219 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_223 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_230 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_244 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_255 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_26 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_260 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_269 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_273 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_276 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_281 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_294 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_3 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_30 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_309 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_315 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_319 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_322 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_347 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_362 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_368 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_413 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_43 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_460 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_47 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_478 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_484 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_494 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_500 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_505 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_516 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_522 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_539 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_550 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_587 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_613 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_622 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_628 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_637 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_667 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_671 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_709 ();
 sky130_as_sc_hs__fill_1 FILLER_0_97_714 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_72 ();
 sky130_as_sc_hs__decap_3 FILLER_0_97_725 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_780 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_785 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_789 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_829 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_833 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_846 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_916 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_932 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_948 ();
 sky130_as_sc_hs__fill_8 FILLER_0_97_953 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_961 ();
 sky130_as_sc_hs__fill_2 FILLER_0_97_965 ();
 sky130_as_sc_hs__decap_4 FILLER_0_97_98 ();
 sky130_as_sc_hs__decap_16 FILLER_0_97_986 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_1010 ();
 sky130_as_sc_hs__fill_8 FILLER_0_98_1026 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_1034 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_1037 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_1053 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_1069 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_107 ();
 sky130_as_sc_hs__fill_1 FILLER_0_98_1091 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_1093 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_1109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_1125 ();
 sky130_as_sc_hs__fill_1 FILLER_0_98_114 ();
 sky130_as_sc_hs__decap_4 FILLER_0_98_1141 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_1145 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_1149 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_1165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_1181 ();
 sky130_as_sc_hs__decap_4 FILLER_0_98_1197 ();
 sky130_as_sc_hs__fill_1 FILLER_0_98_120 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_1201 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_1205 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_1221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_1237 ();
 sky130_as_sc_hs__decap_4 FILLER_0_98_1253 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_1257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_98_126 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_1261 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_137 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_146 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_164 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_169 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_17 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_183 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_188 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_192 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_197 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_211 ();
 sky130_as_sc_hs__fill_1 FILLER_0_98_220 ();
 sky130_as_sc_hs__decap_4 FILLER_0_98_236 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_253 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_26 ();
 sky130_as_sc_hs__decap_4 FILLER_0_98_262 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_29 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_3 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_309 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_321 ();
 sky130_as_sc_hs__fill_1 FILLER_0_98_334 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_360 ();
 sky130_as_sc_hs__decap_4 FILLER_0_98_370 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_376 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_407 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_418 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_42 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_443 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_46 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_461 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_473 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_477 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_486 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_50 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_514 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_580 ();
 sky130_as_sc_hs__fill_1 FILLER_0_98_587 ();
 sky130_as_sc_hs__fill_1 FILLER_0_98_608 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_641 ();
 sky130_as_sc_hs__fill_1 FILLER_0_98_650 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_69 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_698 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_706 ();
 sky130_as_sc_hs__fill_1 FILLER_0_98_757 ();
 sky130_as_sc_hs__decap_4 FILLER_0_98_77 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_785 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_789 ();
 sky130_as_sc_hs__fill_1 FILLER_0_98_81 ();
 sky130_as_sc_hs__decap_4 FILLER_0_98_813 ();
 sky130_as_sc_hs__fill_1 FILLER_0_98_817 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_85 ();
 sky130_as_sc_hs__fill_1 FILLER_0_98_867 ();
 sky130_as_sc_hs__decap_4 FILLER_0_98_869 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_873 ();
 sky130_as_sc_hs__fill_8 FILLER_0_98_884 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_892 ();
 sky130_as_sc_hs__decap_4 FILLER_0_98_898 ();
 sky130_as_sc_hs__fill_1 FILLER_0_98_902 ();
 sky130_as_sc_hs__fill_8 FILLER_0_98_913 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_921 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_925 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_941 ();
 sky130_as_sc_hs__decap_16 FILLER_0_98_957 ();
 sky130_as_sc_hs__decap_4 FILLER_0_98_973 ();
 sky130_as_sc_hs__decap_3 FILLER_0_98_977 ();
 sky130_as_sc_hs__fill_8 FILLER_0_98_981 ();
 sky130_as_sc_hs__fill_2 FILLER_0_98_989 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_1005 ();
 sky130_as_sc_hs__fill_8 FILLER_0_99_1009 ();
 sky130_as_sc_hs__decap_4 FILLER_0_99_1017 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_1021 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_1040 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_1044 ();
 sky130_as_sc_hs__decap_4 FILLER_0_99_1060 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_1081 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_99_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_1121 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_99_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_99_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_99_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_99_1273 ();
 sky130_as_sc_hs__fill_1 FILLER_0_99_130 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_141 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_151 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_160 ();
 sky130_as_sc_hs__fill_1 FILLER_0_99_199 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_205 ();
 sky130_as_sc_hs__fill_1 FILLER_0_99_225 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_276 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_281 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_298 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_308 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_317 ();
 sky130_as_sc_hs__fill_1 FILLER_0_99_330 ();
 sky130_as_sc_hs__decap_4 FILLER_0_99_337 ();
 sky130_as_sc_hs__decap_4 FILLER_0_99_353 ();
 sky130_as_sc_hs__fill_1 FILLER_0_99_357 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_360 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_364 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_368 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_382 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_42 ();
 sky130_as_sc_hs__fill_1 FILLER_0_99_431 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_457 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_462 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_476 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_488 ();
 sky130_as_sc_hs__fill_1 FILLER_0_99_495 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_501 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_505 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_526 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_57 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_575 ();
 sky130_as_sc_hs__fill_1 FILLER_0_99_601 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_612 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_645 ();
 sky130_as_sc_hs__fill_1 FILLER_0_99_671 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_729 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_774 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_797 ();
 sky130_as_sc_hs__fill_8 FILLER_0_99_801 ();
 sky130_as_sc_hs__fill_8 FILLER_0_99_828 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_836 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_857 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_861 ();
 sky130_as_sc_hs__fill_8 FILLER_0_99_868 ();
 sky130_as_sc_hs__decap_4 FILLER_0_99_876 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_880 ();
 sky130_as_sc_hs__decap_3 FILLER_0_99_893 ();
 sky130_as_sc_hs__decap_4 FILLER_0_99_91 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_923 ();
 sky130_as_sc_hs__fill_8 FILLER_0_99_939 ();
 sky130_as_sc_hs__decap_4 FILLER_0_99_947 ();
 sky130_as_sc_hs__fill_1 FILLER_0_99_95 ();
 sky130_as_sc_hs__fill_1 FILLER_0_99_951 ();
 sky130_as_sc_hs__decap_16 FILLER_0_99_953 ();
 sky130_as_sc_hs__decap_4 FILLER_0_99_969 ();
 sky130_as_sc_hs__fill_1 FILLER_0_99_973 ();
 sky130_as_sc_hs__fill_2 FILLER_0_99_98 ();
 sky130_as_sc_hs__fill_8 FILLER_0_99_997 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_1005 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1009 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1025 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1041 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_105 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_1057 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_1061 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1065 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1081 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_109 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1097 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_1113 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_1117 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1121 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_113 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1137 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1153 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_1169 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_1173 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1177 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1193 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1209 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_1225 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_1229 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1233 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_1249 ();
 sky130_as_sc_hs__fill_8 FILLER_0_9_1265 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_1273 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_129 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_145 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_161 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_165 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_169 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_185 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_19 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_201 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_217 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_221 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_225 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_241 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_257 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_273 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_277 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_281 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_297 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_3 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_313 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_329 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_333 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_337 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_35 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_353 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_357 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_382 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_391 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_398 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_406 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_428 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_432 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_445 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_454 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_458 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_462 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_473 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_51 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_513 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_517 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_539 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_545 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_55 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_554 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_558 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_561 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_57 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_587 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_607 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_617 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_645 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_657 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_668 ();
 sky130_as_sc_hs__fill_8 FILLER_0_9_673 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_686 ();
 sky130_as_sc_hs__decap_4 FILLER_0_9_722 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_726 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_73 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_737 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_753 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_757 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_774 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_783 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_812 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_838 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_841 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_851 ();
 sky130_as_sc_hs__decap_3 FILLER_0_9_855 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_89 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_890 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_894 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_897 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_918 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_925 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_929 ();
 sky130_as_sc_hs__fill_1 FILLER_0_9_951 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_953 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_957 ();
 sky130_as_sc_hs__fill_2 FILLER_0_9_961 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_965 ();
 sky130_as_sc_hs__decap_16 FILLER_0_9_981 ();
 sky130_as_sc_hs__fill_8 FILLER_0_9_997 ();
 sky130_as_sc_hs__decap_3 PHY_0 ();
 sky130_as_sc_hs__decap_3 PHY_1 ();
 sky130_as_sc_hs__decap_3 PHY_10 ();
 sky130_as_sc_hs__decap_3 PHY_100 ();
 sky130_as_sc_hs__decap_3 PHY_101 ();
 sky130_as_sc_hs__decap_3 PHY_102 ();
 sky130_as_sc_hs__decap_3 PHY_103 ();
 sky130_as_sc_hs__decap_3 PHY_104 ();
 sky130_as_sc_hs__decap_3 PHY_105 ();
 sky130_as_sc_hs__decap_3 PHY_106 ();
 sky130_as_sc_hs__decap_3 PHY_107 ();
 sky130_as_sc_hs__decap_3 PHY_108 ();
 sky130_as_sc_hs__decap_3 PHY_109 ();
 sky130_as_sc_hs__decap_3 PHY_11 ();
 sky130_as_sc_hs__decap_3 PHY_110 ();
 sky130_as_sc_hs__decap_3 PHY_111 ();
 sky130_as_sc_hs__decap_3 PHY_112 ();
 sky130_as_sc_hs__decap_3 PHY_113 ();
 sky130_as_sc_hs__decap_3 PHY_114 ();
 sky130_as_sc_hs__decap_3 PHY_115 ();
 sky130_as_sc_hs__decap_3 PHY_116 ();
 sky130_as_sc_hs__decap_3 PHY_117 ();
 sky130_as_sc_hs__decap_3 PHY_118 ();
 sky130_as_sc_hs__decap_3 PHY_119 ();
 sky130_as_sc_hs__decap_3 PHY_12 ();
 sky130_as_sc_hs__decap_3 PHY_120 ();
 sky130_as_sc_hs__decap_3 PHY_121 ();
 sky130_as_sc_hs__decap_3 PHY_122 ();
 sky130_as_sc_hs__decap_3 PHY_123 ();
 sky130_as_sc_hs__decap_3 PHY_124 ();
 sky130_as_sc_hs__decap_3 PHY_125 ();
 sky130_as_sc_hs__decap_3 PHY_126 ();
 sky130_as_sc_hs__decap_3 PHY_127 ();
 sky130_as_sc_hs__decap_3 PHY_128 ();
 sky130_as_sc_hs__decap_3 PHY_129 ();
 sky130_as_sc_hs__decap_3 PHY_13 ();
 sky130_as_sc_hs__decap_3 PHY_130 ();
 sky130_as_sc_hs__decap_3 PHY_131 ();
 sky130_as_sc_hs__decap_3 PHY_132 ();
 sky130_as_sc_hs__decap_3 PHY_133 ();
 sky130_as_sc_hs__decap_3 PHY_134 ();
 sky130_as_sc_hs__decap_3 PHY_135 ();
 sky130_as_sc_hs__decap_3 PHY_136 ();
 sky130_as_sc_hs__decap_3 PHY_137 ();
 sky130_as_sc_hs__decap_3 PHY_138 ();
 sky130_as_sc_hs__decap_3 PHY_139 ();
 sky130_as_sc_hs__decap_3 PHY_14 ();
 sky130_as_sc_hs__decap_3 PHY_140 ();
 sky130_as_sc_hs__decap_3 PHY_141 ();
 sky130_as_sc_hs__decap_3 PHY_142 ();
 sky130_as_sc_hs__decap_3 PHY_143 ();
 sky130_as_sc_hs__decap_3 PHY_144 ();
 sky130_as_sc_hs__decap_3 PHY_145 ();
 sky130_as_sc_hs__decap_3 PHY_146 ();
 sky130_as_sc_hs__decap_3 PHY_147 ();
 sky130_as_sc_hs__decap_3 PHY_148 ();
 sky130_as_sc_hs__decap_3 PHY_149 ();
 sky130_as_sc_hs__decap_3 PHY_15 ();
 sky130_as_sc_hs__decap_3 PHY_150 ();
 sky130_as_sc_hs__decap_3 PHY_151 ();
 sky130_as_sc_hs__decap_3 PHY_152 ();
 sky130_as_sc_hs__decap_3 PHY_153 ();
 sky130_as_sc_hs__decap_3 PHY_154 ();
 sky130_as_sc_hs__decap_3 PHY_155 ();
 sky130_as_sc_hs__decap_3 PHY_156 ();
 sky130_as_sc_hs__decap_3 PHY_157 ();
 sky130_as_sc_hs__decap_3 PHY_158 ();
 sky130_as_sc_hs__decap_3 PHY_159 ();
 sky130_as_sc_hs__decap_3 PHY_16 ();
 sky130_as_sc_hs__decap_3 PHY_160 ();
 sky130_as_sc_hs__decap_3 PHY_161 ();
 sky130_as_sc_hs__decap_3 PHY_162 ();
 sky130_as_sc_hs__decap_3 PHY_163 ();
 sky130_as_sc_hs__decap_3 PHY_164 ();
 sky130_as_sc_hs__decap_3 PHY_165 ();
 sky130_as_sc_hs__decap_3 PHY_166 ();
 sky130_as_sc_hs__decap_3 PHY_167 ();
 sky130_as_sc_hs__decap_3 PHY_168 ();
 sky130_as_sc_hs__decap_3 PHY_169 ();
 sky130_as_sc_hs__decap_3 PHY_17 ();
 sky130_as_sc_hs__decap_3 PHY_170 ();
 sky130_as_sc_hs__decap_3 PHY_171 ();
 sky130_as_sc_hs__decap_3 PHY_172 ();
 sky130_as_sc_hs__decap_3 PHY_173 ();
 sky130_as_sc_hs__decap_3 PHY_174 ();
 sky130_as_sc_hs__decap_3 PHY_175 ();
 sky130_as_sc_hs__decap_3 PHY_176 ();
 sky130_as_sc_hs__decap_3 PHY_177 ();
 sky130_as_sc_hs__decap_3 PHY_178 ();
 sky130_as_sc_hs__decap_3 PHY_179 ();
 sky130_as_sc_hs__decap_3 PHY_18 ();
 sky130_as_sc_hs__decap_3 PHY_180 ();
 sky130_as_sc_hs__decap_3 PHY_181 ();
 sky130_as_sc_hs__decap_3 PHY_182 ();
 sky130_as_sc_hs__decap_3 PHY_183 ();
 sky130_as_sc_hs__decap_3 PHY_184 ();
 sky130_as_sc_hs__decap_3 PHY_185 ();
 sky130_as_sc_hs__decap_3 PHY_186 ();
 sky130_as_sc_hs__decap_3 PHY_187 ();
 sky130_as_sc_hs__decap_3 PHY_188 ();
 sky130_as_sc_hs__decap_3 PHY_189 ();
 sky130_as_sc_hs__decap_3 PHY_19 ();
 sky130_as_sc_hs__decap_3 PHY_190 ();
 sky130_as_sc_hs__decap_3 PHY_191 ();
 sky130_as_sc_hs__decap_3 PHY_192 ();
 sky130_as_sc_hs__decap_3 PHY_193 ();
 sky130_as_sc_hs__decap_3 PHY_194 ();
 sky130_as_sc_hs__decap_3 PHY_195 ();
 sky130_as_sc_hs__decap_3 PHY_196 ();
 sky130_as_sc_hs__decap_3 PHY_197 ();
 sky130_as_sc_hs__decap_3 PHY_198 ();
 sky130_as_sc_hs__decap_3 PHY_199 ();
 sky130_as_sc_hs__decap_3 PHY_2 ();
 sky130_as_sc_hs__decap_3 PHY_20 ();
 sky130_as_sc_hs__decap_3 PHY_200 ();
 sky130_as_sc_hs__decap_3 PHY_201 ();
 sky130_as_sc_hs__decap_3 PHY_202 ();
 sky130_as_sc_hs__decap_3 PHY_203 ();
 sky130_as_sc_hs__decap_3 PHY_204 ();
 sky130_as_sc_hs__decap_3 PHY_205 ();
 sky130_as_sc_hs__decap_3 PHY_206 ();
 sky130_as_sc_hs__decap_3 PHY_207 ();
 sky130_as_sc_hs__decap_3 PHY_208 ();
 sky130_as_sc_hs__decap_3 PHY_209 ();
 sky130_as_sc_hs__decap_3 PHY_21 ();
 sky130_as_sc_hs__decap_3 PHY_210 ();
 sky130_as_sc_hs__decap_3 PHY_211 ();
 sky130_as_sc_hs__decap_3 PHY_212 ();
 sky130_as_sc_hs__decap_3 PHY_213 ();
 sky130_as_sc_hs__decap_3 PHY_214 ();
 sky130_as_sc_hs__decap_3 PHY_215 ();
 sky130_as_sc_hs__decap_3 PHY_216 ();
 sky130_as_sc_hs__decap_3 PHY_217 ();
 sky130_as_sc_hs__decap_3 PHY_218 ();
 sky130_as_sc_hs__decap_3 PHY_219 ();
 sky130_as_sc_hs__decap_3 PHY_22 ();
 sky130_as_sc_hs__decap_3 PHY_220 ();
 sky130_as_sc_hs__decap_3 PHY_221 ();
 sky130_as_sc_hs__decap_3 PHY_222 ();
 sky130_as_sc_hs__decap_3 PHY_223 ();
 sky130_as_sc_hs__decap_3 PHY_224 ();
 sky130_as_sc_hs__decap_3 PHY_225 ();
 sky130_as_sc_hs__decap_3 PHY_226 ();
 sky130_as_sc_hs__decap_3 PHY_227 ();
 sky130_as_sc_hs__decap_3 PHY_228 ();
 sky130_as_sc_hs__decap_3 PHY_229 ();
 sky130_as_sc_hs__decap_3 PHY_23 ();
 sky130_as_sc_hs__decap_3 PHY_230 ();
 sky130_as_sc_hs__decap_3 PHY_231 ();
 sky130_as_sc_hs__decap_3 PHY_232 ();
 sky130_as_sc_hs__decap_3 PHY_233 ();
 sky130_as_sc_hs__decap_3 PHY_234 ();
 sky130_as_sc_hs__decap_3 PHY_235 ();
 sky130_as_sc_hs__decap_3 PHY_236 ();
 sky130_as_sc_hs__decap_3 PHY_237 ();
 sky130_as_sc_hs__decap_3 PHY_238 ();
 sky130_as_sc_hs__decap_3 PHY_239 ();
 sky130_as_sc_hs__decap_3 PHY_24 ();
 sky130_as_sc_hs__decap_3 PHY_240 ();
 sky130_as_sc_hs__decap_3 PHY_241 ();
 sky130_as_sc_hs__decap_3 PHY_242 ();
 sky130_as_sc_hs__decap_3 PHY_243 ();
 sky130_as_sc_hs__decap_3 PHY_244 ();
 sky130_as_sc_hs__decap_3 PHY_245 ();
 sky130_as_sc_hs__decap_3 PHY_246 ();
 sky130_as_sc_hs__decap_3 PHY_247 ();
 sky130_as_sc_hs__decap_3 PHY_248 ();
 sky130_as_sc_hs__decap_3 PHY_249 ();
 sky130_as_sc_hs__decap_3 PHY_25 ();
 sky130_as_sc_hs__decap_3 PHY_250 ();
 sky130_as_sc_hs__decap_3 PHY_251 ();
 sky130_as_sc_hs__decap_3 PHY_252 ();
 sky130_as_sc_hs__decap_3 PHY_253 ();
 sky130_as_sc_hs__decap_3 PHY_254 ();
 sky130_as_sc_hs__decap_3 PHY_255 ();
 sky130_as_sc_hs__decap_3 PHY_256 ();
 sky130_as_sc_hs__decap_3 PHY_257 ();
 sky130_as_sc_hs__decap_3 PHY_258 ();
 sky130_as_sc_hs__decap_3 PHY_259 ();
 sky130_as_sc_hs__decap_3 PHY_26 ();
 sky130_as_sc_hs__decap_3 PHY_260 ();
 sky130_as_sc_hs__decap_3 PHY_261 ();
 sky130_as_sc_hs__decap_3 PHY_262 ();
 sky130_as_sc_hs__decap_3 PHY_263 ();
 sky130_as_sc_hs__decap_3 PHY_264 ();
 sky130_as_sc_hs__decap_3 PHY_265 ();
 sky130_as_sc_hs__decap_3 PHY_266 ();
 sky130_as_sc_hs__decap_3 PHY_267 ();
 sky130_as_sc_hs__decap_3 PHY_268 ();
 sky130_as_sc_hs__decap_3 PHY_269 ();
 sky130_as_sc_hs__decap_3 PHY_27 ();
 sky130_as_sc_hs__decap_3 PHY_270 ();
 sky130_as_sc_hs__decap_3 PHY_271 ();
 sky130_as_sc_hs__decap_3 PHY_272 ();
 sky130_as_sc_hs__decap_3 PHY_273 ();
 sky130_as_sc_hs__decap_3 PHY_274 ();
 sky130_as_sc_hs__decap_3 PHY_275 ();
 sky130_as_sc_hs__decap_3 PHY_276 ();
 sky130_as_sc_hs__decap_3 PHY_277 ();
 sky130_as_sc_hs__decap_3 PHY_278 ();
 sky130_as_sc_hs__decap_3 PHY_279 ();
 sky130_as_sc_hs__decap_3 PHY_28 ();
 sky130_as_sc_hs__decap_3 PHY_280 ();
 sky130_as_sc_hs__decap_3 PHY_281 ();
 sky130_as_sc_hs__decap_3 PHY_282 ();
 sky130_as_sc_hs__decap_3 PHY_283 ();
 sky130_as_sc_hs__decap_3 PHY_284 ();
 sky130_as_sc_hs__decap_3 PHY_285 ();
 sky130_as_sc_hs__decap_3 PHY_286 ();
 sky130_as_sc_hs__decap_3 PHY_287 ();
 sky130_as_sc_hs__decap_3 PHY_288 ();
 sky130_as_sc_hs__decap_3 PHY_289 ();
 sky130_as_sc_hs__decap_3 PHY_29 ();
 sky130_as_sc_hs__decap_3 PHY_290 ();
 sky130_as_sc_hs__decap_3 PHY_291 ();
 sky130_as_sc_hs__decap_3 PHY_292 ();
 sky130_as_sc_hs__decap_3 PHY_293 ();
 sky130_as_sc_hs__decap_3 PHY_294 ();
 sky130_as_sc_hs__decap_3 PHY_295 ();
 sky130_as_sc_hs__decap_3 PHY_296 ();
 sky130_as_sc_hs__decap_3 PHY_297 ();
 sky130_as_sc_hs__decap_3 PHY_298 ();
 sky130_as_sc_hs__decap_3 PHY_299 ();
 sky130_as_sc_hs__decap_3 PHY_3 ();
 sky130_as_sc_hs__decap_3 PHY_30 ();
 sky130_as_sc_hs__decap_3 PHY_300 ();
 sky130_as_sc_hs__decap_3 PHY_301 ();
 sky130_as_sc_hs__decap_3 PHY_302 ();
 sky130_as_sc_hs__decap_3 PHY_303 ();
 sky130_as_sc_hs__decap_3 PHY_304 ();
 sky130_as_sc_hs__decap_3 PHY_305 ();
 sky130_as_sc_hs__decap_3 PHY_306 ();
 sky130_as_sc_hs__decap_3 PHY_307 ();
 sky130_as_sc_hs__decap_3 PHY_308 ();
 sky130_as_sc_hs__decap_3 PHY_309 ();
 sky130_as_sc_hs__decap_3 PHY_31 ();
 sky130_as_sc_hs__decap_3 PHY_310 ();
 sky130_as_sc_hs__decap_3 PHY_311 ();
 sky130_as_sc_hs__decap_3 PHY_312 ();
 sky130_as_sc_hs__decap_3 PHY_313 ();
 sky130_as_sc_hs__decap_3 PHY_314 ();
 sky130_as_sc_hs__decap_3 PHY_315 ();
 sky130_as_sc_hs__decap_3 PHY_316 ();
 sky130_as_sc_hs__decap_3 PHY_317 ();
 sky130_as_sc_hs__decap_3 PHY_318 ();
 sky130_as_sc_hs__decap_3 PHY_319 ();
 sky130_as_sc_hs__decap_3 PHY_32 ();
 sky130_as_sc_hs__decap_3 PHY_320 ();
 sky130_as_sc_hs__decap_3 PHY_321 ();
 sky130_as_sc_hs__decap_3 PHY_322 ();
 sky130_as_sc_hs__decap_3 PHY_323 ();
 sky130_as_sc_hs__decap_3 PHY_324 ();
 sky130_as_sc_hs__decap_3 PHY_325 ();
 sky130_as_sc_hs__decap_3 PHY_326 ();
 sky130_as_sc_hs__decap_3 PHY_327 ();
 sky130_as_sc_hs__decap_3 PHY_328 ();
 sky130_as_sc_hs__decap_3 PHY_329 ();
 sky130_as_sc_hs__decap_3 PHY_33 ();
 sky130_as_sc_hs__decap_3 PHY_330 ();
 sky130_as_sc_hs__decap_3 PHY_331 ();
 sky130_as_sc_hs__decap_3 PHY_332 ();
 sky130_as_sc_hs__decap_3 PHY_333 ();
 sky130_as_sc_hs__decap_3 PHY_334 ();
 sky130_as_sc_hs__decap_3 PHY_335 ();
 sky130_as_sc_hs__decap_3 PHY_336 ();
 sky130_as_sc_hs__decap_3 PHY_337 ();
 sky130_as_sc_hs__decap_3 PHY_338 ();
 sky130_as_sc_hs__decap_3 PHY_339 ();
 sky130_as_sc_hs__decap_3 PHY_34 ();
 sky130_as_sc_hs__decap_3 PHY_340 ();
 sky130_as_sc_hs__decap_3 PHY_341 ();
 sky130_as_sc_hs__decap_3 PHY_342 ();
 sky130_as_sc_hs__decap_3 PHY_343 ();
 sky130_as_sc_hs__decap_3 PHY_344 ();
 sky130_as_sc_hs__decap_3 PHY_345 ();
 sky130_as_sc_hs__decap_3 PHY_346 ();
 sky130_as_sc_hs__decap_3 PHY_347 ();
 sky130_as_sc_hs__decap_3 PHY_348 ();
 sky130_as_sc_hs__decap_3 PHY_349 ();
 sky130_as_sc_hs__decap_3 PHY_35 ();
 sky130_as_sc_hs__decap_3 PHY_350 ();
 sky130_as_sc_hs__decap_3 PHY_351 ();
 sky130_as_sc_hs__decap_3 PHY_352 ();
 sky130_as_sc_hs__decap_3 PHY_353 ();
 sky130_as_sc_hs__decap_3 PHY_354 ();
 sky130_as_sc_hs__decap_3 PHY_355 ();
 sky130_as_sc_hs__decap_3 PHY_356 ();
 sky130_as_sc_hs__decap_3 PHY_357 ();
 sky130_as_sc_hs__decap_3 PHY_358 ();
 sky130_as_sc_hs__decap_3 PHY_359 ();
 sky130_as_sc_hs__decap_3 PHY_36 ();
 sky130_as_sc_hs__decap_3 PHY_360 ();
 sky130_as_sc_hs__decap_3 PHY_361 ();
 sky130_as_sc_hs__decap_3 PHY_362 ();
 sky130_as_sc_hs__decap_3 PHY_363 ();
 sky130_as_sc_hs__decap_3 PHY_364 ();
 sky130_as_sc_hs__decap_3 PHY_365 ();
 sky130_as_sc_hs__decap_3 PHY_366 ();
 sky130_as_sc_hs__decap_3 PHY_367 ();
 sky130_as_sc_hs__decap_3 PHY_368 ();
 sky130_as_sc_hs__decap_3 PHY_369 ();
 sky130_as_sc_hs__decap_3 PHY_37 ();
 sky130_as_sc_hs__decap_3 PHY_370 ();
 sky130_as_sc_hs__decap_3 PHY_371 ();
 sky130_as_sc_hs__decap_3 PHY_372 ();
 sky130_as_sc_hs__decap_3 PHY_373 ();
 sky130_as_sc_hs__decap_3 PHY_374 ();
 sky130_as_sc_hs__decap_3 PHY_375 ();
 sky130_as_sc_hs__decap_3 PHY_376 ();
 sky130_as_sc_hs__decap_3 PHY_377 ();
 sky130_as_sc_hs__decap_3 PHY_378 ();
 sky130_as_sc_hs__decap_3 PHY_379 ();
 sky130_as_sc_hs__decap_3 PHY_38 ();
 sky130_as_sc_hs__decap_3 PHY_380 ();
 sky130_as_sc_hs__decap_3 PHY_381 ();
 sky130_as_sc_hs__decap_3 PHY_382 ();
 sky130_as_sc_hs__decap_3 PHY_383 ();
 sky130_as_sc_hs__decap_3 PHY_384 ();
 sky130_as_sc_hs__decap_3 PHY_385 ();
 sky130_as_sc_hs__decap_3 PHY_386 ();
 sky130_as_sc_hs__decap_3 PHY_387 ();
 sky130_as_sc_hs__decap_3 PHY_388 ();
 sky130_as_sc_hs__decap_3 PHY_389 ();
 sky130_as_sc_hs__decap_3 PHY_39 ();
 sky130_as_sc_hs__decap_3 PHY_390 ();
 sky130_as_sc_hs__decap_3 PHY_391 ();
 sky130_as_sc_hs__decap_3 PHY_392 ();
 sky130_as_sc_hs__decap_3 PHY_393 ();
 sky130_as_sc_hs__decap_3 PHY_394 ();
 sky130_as_sc_hs__decap_3 PHY_395 ();
 sky130_as_sc_hs__decap_3 PHY_396 ();
 sky130_as_sc_hs__decap_3 PHY_397 ();
 sky130_as_sc_hs__decap_3 PHY_398 ();
 sky130_as_sc_hs__decap_3 PHY_399 ();
 sky130_as_sc_hs__decap_3 PHY_4 ();
 sky130_as_sc_hs__decap_3 PHY_40 ();
 sky130_as_sc_hs__decap_3 PHY_400 ();
 sky130_as_sc_hs__decap_3 PHY_401 ();
 sky130_as_sc_hs__decap_3 PHY_402 ();
 sky130_as_sc_hs__decap_3 PHY_403 ();
 sky130_as_sc_hs__decap_3 PHY_404 ();
 sky130_as_sc_hs__decap_3 PHY_405 ();
 sky130_as_sc_hs__decap_3 PHY_406 ();
 sky130_as_sc_hs__decap_3 PHY_407 ();
 sky130_as_sc_hs__decap_3 PHY_408 ();
 sky130_as_sc_hs__decap_3 PHY_409 ();
 sky130_as_sc_hs__decap_3 PHY_41 ();
 sky130_as_sc_hs__decap_3 PHY_410 ();
 sky130_as_sc_hs__decap_3 PHY_411 ();
 sky130_as_sc_hs__decap_3 PHY_412 ();
 sky130_as_sc_hs__decap_3 PHY_413 ();
 sky130_as_sc_hs__decap_3 PHY_414 ();
 sky130_as_sc_hs__decap_3 PHY_415 ();
 sky130_as_sc_hs__decap_3 PHY_416 ();
 sky130_as_sc_hs__decap_3 PHY_417 ();
 sky130_as_sc_hs__decap_3 PHY_418 ();
 sky130_as_sc_hs__decap_3 PHY_419 ();
 sky130_as_sc_hs__decap_3 PHY_42 ();
 sky130_as_sc_hs__decap_3 PHY_420 ();
 sky130_as_sc_hs__decap_3 PHY_421 ();
 sky130_as_sc_hs__decap_3 PHY_422 ();
 sky130_as_sc_hs__decap_3 PHY_423 ();
 sky130_as_sc_hs__decap_3 PHY_43 ();
 sky130_as_sc_hs__decap_3 PHY_44 ();
 sky130_as_sc_hs__decap_3 PHY_45 ();
 sky130_as_sc_hs__decap_3 PHY_46 ();
 sky130_as_sc_hs__decap_3 PHY_47 ();
 sky130_as_sc_hs__decap_3 PHY_48 ();
 sky130_as_sc_hs__decap_3 PHY_49 ();
 sky130_as_sc_hs__decap_3 PHY_5 ();
 sky130_as_sc_hs__decap_3 PHY_50 ();
 sky130_as_sc_hs__decap_3 PHY_51 ();
 sky130_as_sc_hs__decap_3 PHY_52 ();
 sky130_as_sc_hs__decap_3 PHY_53 ();
 sky130_as_sc_hs__decap_3 PHY_54 ();
 sky130_as_sc_hs__decap_3 PHY_55 ();
 sky130_as_sc_hs__decap_3 PHY_56 ();
 sky130_as_sc_hs__decap_3 PHY_57 ();
 sky130_as_sc_hs__decap_3 PHY_58 ();
 sky130_as_sc_hs__decap_3 PHY_59 ();
 sky130_as_sc_hs__decap_3 PHY_6 ();
 sky130_as_sc_hs__decap_3 PHY_60 ();
 sky130_as_sc_hs__decap_3 PHY_61 ();
 sky130_as_sc_hs__decap_3 PHY_62 ();
 sky130_as_sc_hs__decap_3 PHY_63 ();
 sky130_as_sc_hs__decap_3 PHY_64 ();
 sky130_as_sc_hs__decap_3 PHY_65 ();
 sky130_as_sc_hs__decap_3 PHY_66 ();
 sky130_as_sc_hs__decap_3 PHY_67 ();
 sky130_as_sc_hs__decap_3 PHY_68 ();
 sky130_as_sc_hs__decap_3 PHY_69 ();
 sky130_as_sc_hs__decap_3 PHY_7 ();
 sky130_as_sc_hs__decap_3 PHY_70 ();
 sky130_as_sc_hs__decap_3 PHY_71 ();
 sky130_as_sc_hs__decap_3 PHY_72 ();
 sky130_as_sc_hs__decap_3 PHY_73 ();
 sky130_as_sc_hs__decap_3 PHY_74 ();
 sky130_as_sc_hs__decap_3 PHY_75 ();
 sky130_as_sc_hs__decap_3 PHY_76 ();
 sky130_as_sc_hs__decap_3 PHY_77 ();
 sky130_as_sc_hs__decap_3 PHY_78 ();
 sky130_as_sc_hs__decap_3 PHY_79 ();
 sky130_as_sc_hs__decap_3 PHY_8 ();
 sky130_as_sc_hs__decap_3 PHY_80 ();
 sky130_as_sc_hs__decap_3 PHY_81 ();
 sky130_as_sc_hs__decap_3 PHY_82 ();
 sky130_as_sc_hs__decap_3 PHY_83 ();
 sky130_as_sc_hs__decap_3 PHY_84 ();
 sky130_as_sc_hs__decap_3 PHY_85 ();
 sky130_as_sc_hs__decap_3 PHY_86 ();
 sky130_as_sc_hs__decap_3 PHY_87 ();
 sky130_as_sc_hs__decap_3 PHY_88 ();
 sky130_as_sc_hs__decap_3 PHY_89 ();
 sky130_as_sc_hs__decap_3 PHY_9 ();
 sky130_as_sc_hs__decap_3 PHY_90 ();
 sky130_as_sc_hs__decap_3 PHY_91 ();
 sky130_as_sc_hs__decap_3 PHY_92 ();
 sky130_as_sc_hs__decap_3 PHY_93 ();
 sky130_as_sc_hs__decap_3 PHY_94 ();
 sky130_as_sc_hs__decap_3 PHY_95 ();
 sky130_as_sc_hs__decap_3 PHY_96 ();
 sky130_as_sc_hs__decap_3 PHY_97 ();
 sky130_as_sc_hs__decap_3 PHY_98 ();
 sky130_as_sc_hs__decap_3 PHY_99 ();
 sky130_as_sc_hs__tap_1 TAP_1000 ();
 sky130_as_sc_hs__tap_1 TAP_1001 ();
 sky130_as_sc_hs__tap_1 TAP_1002 ();
 sky130_as_sc_hs__tap_1 TAP_1003 ();
 sky130_as_sc_hs__tap_1 TAP_1004 ();
 sky130_as_sc_hs__tap_1 TAP_1005 ();
 sky130_as_sc_hs__tap_1 TAP_1006 ();
 sky130_as_sc_hs__tap_1 TAP_1007 ();
 sky130_as_sc_hs__tap_1 TAP_1008 ();
 sky130_as_sc_hs__tap_1 TAP_1009 ();
 sky130_as_sc_hs__tap_1 TAP_1010 ();
 sky130_as_sc_hs__tap_1 TAP_1011 ();
 sky130_as_sc_hs__tap_1 TAP_1012 ();
 sky130_as_sc_hs__tap_1 TAP_1013 ();
 sky130_as_sc_hs__tap_1 TAP_1014 ();
 sky130_as_sc_hs__tap_1 TAP_1015 ();
 sky130_as_sc_hs__tap_1 TAP_1016 ();
 sky130_as_sc_hs__tap_1 TAP_1017 ();
 sky130_as_sc_hs__tap_1 TAP_1018 ();
 sky130_as_sc_hs__tap_1 TAP_1019 ();
 sky130_as_sc_hs__tap_1 TAP_1020 ();
 sky130_as_sc_hs__tap_1 TAP_1021 ();
 sky130_as_sc_hs__tap_1 TAP_1022 ();
 sky130_as_sc_hs__tap_1 TAP_1023 ();
 sky130_as_sc_hs__tap_1 TAP_1024 ();
 sky130_as_sc_hs__tap_1 TAP_1025 ();
 sky130_as_sc_hs__tap_1 TAP_1026 ();
 sky130_as_sc_hs__tap_1 TAP_1027 ();
 sky130_as_sc_hs__tap_1 TAP_1028 ();
 sky130_as_sc_hs__tap_1 TAP_1029 ();
 sky130_as_sc_hs__tap_1 TAP_1030 ();
 sky130_as_sc_hs__tap_1 TAP_1031 ();
 sky130_as_sc_hs__tap_1 TAP_1032 ();
 sky130_as_sc_hs__tap_1 TAP_1033 ();
 sky130_as_sc_hs__tap_1 TAP_1034 ();
 sky130_as_sc_hs__tap_1 TAP_1035 ();
 sky130_as_sc_hs__tap_1 TAP_1036 ();
 sky130_as_sc_hs__tap_1 TAP_1037 ();
 sky130_as_sc_hs__tap_1 TAP_1038 ();
 sky130_as_sc_hs__tap_1 TAP_1039 ();
 sky130_as_sc_hs__tap_1 TAP_1040 ();
 sky130_as_sc_hs__tap_1 TAP_1041 ();
 sky130_as_sc_hs__tap_1 TAP_1042 ();
 sky130_as_sc_hs__tap_1 TAP_1043 ();
 sky130_as_sc_hs__tap_1 TAP_1044 ();
 sky130_as_sc_hs__tap_1 TAP_1045 ();
 sky130_as_sc_hs__tap_1 TAP_1046 ();
 sky130_as_sc_hs__tap_1 TAP_1047 ();
 sky130_as_sc_hs__tap_1 TAP_1048 ();
 sky130_as_sc_hs__tap_1 TAP_1049 ();
 sky130_as_sc_hs__tap_1 TAP_1050 ();
 sky130_as_sc_hs__tap_1 TAP_1051 ();
 sky130_as_sc_hs__tap_1 TAP_1052 ();
 sky130_as_sc_hs__tap_1 TAP_1053 ();
 sky130_as_sc_hs__tap_1 TAP_1054 ();
 sky130_as_sc_hs__tap_1 TAP_1055 ();
 sky130_as_sc_hs__tap_1 TAP_1056 ();
 sky130_as_sc_hs__tap_1 TAP_1057 ();
 sky130_as_sc_hs__tap_1 TAP_1058 ();
 sky130_as_sc_hs__tap_1 TAP_1059 ();
 sky130_as_sc_hs__tap_1 TAP_1060 ();
 sky130_as_sc_hs__tap_1 TAP_1061 ();
 sky130_as_sc_hs__tap_1 TAP_1062 ();
 sky130_as_sc_hs__tap_1 TAP_1063 ();
 sky130_as_sc_hs__tap_1 TAP_1064 ();
 sky130_as_sc_hs__tap_1 TAP_1065 ();
 sky130_as_sc_hs__tap_1 TAP_1066 ();
 sky130_as_sc_hs__tap_1 TAP_1067 ();
 sky130_as_sc_hs__tap_1 TAP_1068 ();
 sky130_as_sc_hs__tap_1 TAP_1069 ();
 sky130_as_sc_hs__tap_1 TAP_1070 ();
 sky130_as_sc_hs__tap_1 TAP_1071 ();
 sky130_as_sc_hs__tap_1 TAP_1072 ();
 sky130_as_sc_hs__tap_1 TAP_1073 ();
 sky130_as_sc_hs__tap_1 TAP_1074 ();
 sky130_as_sc_hs__tap_1 TAP_1075 ();
 sky130_as_sc_hs__tap_1 TAP_1076 ();
 sky130_as_sc_hs__tap_1 TAP_1077 ();
 sky130_as_sc_hs__tap_1 TAP_1078 ();
 sky130_as_sc_hs__tap_1 TAP_1079 ();
 sky130_as_sc_hs__tap_1 TAP_1080 ();
 sky130_as_sc_hs__tap_1 TAP_1081 ();
 sky130_as_sc_hs__tap_1 TAP_1082 ();
 sky130_as_sc_hs__tap_1 TAP_1083 ();
 sky130_as_sc_hs__tap_1 TAP_1084 ();
 sky130_as_sc_hs__tap_1 TAP_1085 ();
 sky130_as_sc_hs__tap_1 TAP_1086 ();
 sky130_as_sc_hs__tap_1 TAP_1087 ();
 sky130_as_sc_hs__tap_1 TAP_1088 ();
 sky130_as_sc_hs__tap_1 TAP_1089 ();
 sky130_as_sc_hs__tap_1 TAP_1090 ();
 sky130_as_sc_hs__tap_1 TAP_1091 ();
 sky130_as_sc_hs__tap_1 TAP_1092 ();
 sky130_as_sc_hs__tap_1 TAP_1093 ();
 sky130_as_sc_hs__tap_1 TAP_1094 ();
 sky130_as_sc_hs__tap_1 TAP_1095 ();
 sky130_as_sc_hs__tap_1 TAP_1096 ();
 sky130_as_sc_hs__tap_1 TAP_1097 ();
 sky130_as_sc_hs__tap_1 TAP_1098 ();
 sky130_as_sc_hs__tap_1 TAP_1099 ();
 sky130_as_sc_hs__tap_1 TAP_1100 ();
 sky130_as_sc_hs__tap_1 TAP_1101 ();
 sky130_as_sc_hs__tap_1 TAP_1102 ();
 sky130_as_sc_hs__tap_1 TAP_1103 ();
 sky130_as_sc_hs__tap_1 TAP_1104 ();
 sky130_as_sc_hs__tap_1 TAP_1105 ();
 sky130_as_sc_hs__tap_1 TAP_1106 ();
 sky130_as_sc_hs__tap_1 TAP_1107 ();
 sky130_as_sc_hs__tap_1 TAP_1108 ();
 sky130_as_sc_hs__tap_1 TAP_1109 ();
 sky130_as_sc_hs__tap_1 TAP_1110 ();
 sky130_as_sc_hs__tap_1 TAP_1111 ();
 sky130_as_sc_hs__tap_1 TAP_1112 ();
 sky130_as_sc_hs__tap_1 TAP_1113 ();
 sky130_as_sc_hs__tap_1 TAP_1114 ();
 sky130_as_sc_hs__tap_1 TAP_1115 ();
 sky130_as_sc_hs__tap_1 TAP_1116 ();
 sky130_as_sc_hs__tap_1 TAP_1117 ();
 sky130_as_sc_hs__tap_1 TAP_1118 ();
 sky130_as_sc_hs__tap_1 TAP_1119 ();
 sky130_as_sc_hs__tap_1 TAP_1120 ();
 sky130_as_sc_hs__tap_1 TAP_1121 ();
 sky130_as_sc_hs__tap_1 TAP_1122 ();
 sky130_as_sc_hs__tap_1 TAP_1123 ();
 sky130_as_sc_hs__tap_1 TAP_1124 ();
 sky130_as_sc_hs__tap_1 TAP_1125 ();
 sky130_as_sc_hs__tap_1 TAP_1126 ();
 sky130_as_sc_hs__tap_1 TAP_1127 ();
 sky130_as_sc_hs__tap_1 TAP_1128 ();
 sky130_as_sc_hs__tap_1 TAP_1129 ();
 sky130_as_sc_hs__tap_1 TAP_1130 ();
 sky130_as_sc_hs__tap_1 TAP_1131 ();
 sky130_as_sc_hs__tap_1 TAP_1132 ();
 sky130_as_sc_hs__tap_1 TAP_1133 ();
 sky130_as_sc_hs__tap_1 TAP_1134 ();
 sky130_as_sc_hs__tap_1 TAP_1135 ();
 sky130_as_sc_hs__tap_1 TAP_1136 ();
 sky130_as_sc_hs__tap_1 TAP_1137 ();
 sky130_as_sc_hs__tap_1 TAP_1138 ();
 sky130_as_sc_hs__tap_1 TAP_1139 ();
 sky130_as_sc_hs__tap_1 TAP_1140 ();
 sky130_as_sc_hs__tap_1 TAP_1141 ();
 sky130_as_sc_hs__tap_1 TAP_1142 ();
 sky130_as_sc_hs__tap_1 TAP_1143 ();
 sky130_as_sc_hs__tap_1 TAP_1144 ();
 sky130_as_sc_hs__tap_1 TAP_1145 ();
 sky130_as_sc_hs__tap_1 TAP_1146 ();
 sky130_as_sc_hs__tap_1 TAP_1147 ();
 sky130_as_sc_hs__tap_1 TAP_1148 ();
 sky130_as_sc_hs__tap_1 TAP_1149 ();
 sky130_as_sc_hs__tap_1 TAP_1150 ();
 sky130_as_sc_hs__tap_1 TAP_1151 ();
 sky130_as_sc_hs__tap_1 TAP_1152 ();
 sky130_as_sc_hs__tap_1 TAP_1153 ();
 sky130_as_sc_hs__tap_1 TAP_1154 ();
 sky130_as_sc_hs__tap_1 TAP_1155 ();
 sky130_as_sc_hs__tap_1 TAP_1156 ();
 sky130_as_sc_hs__tap_1 TAP_1157 ();
 sky130_as_sc_hs__tap_1 TAP_1158 ();
 sky130_as_sc_hs__tap_1 TAP_1159 ();
 sky130_as_sc_hs__tap_1 TAP_1160 ();
 sky130_as_sc_hs__tap_1 TAP_1161 ();
 sky130_as_sc_hs__tap_1 TAP_1162 ();
 sky130_as_sc_hs__tap_1 TAP_1163 ();
 sky130_as_sc_hs__tap_1 TAP_1164 ();
 sky130_as_sc_hs__tap_1 TAP_1165 ();
 sky130_as_sc_hs__tap_1 TAP_1166 ();
 sky130_as_sc_hs__tap_1 TAP_1167 ();
 sky130_as_sc_hs__tap_1 TAP_1168 ();
 sky130_as_sc_hs__tap_1 TAP_1169 ();
 sky130_as_sc_hs__tap_1 TAP_1170 ();
 sky130_as_sc_hs__tap_1 TAP_1171 ();
 sky130_as_sc_hs__tap_1 TAP_1172 ();
 sky130_as_sc_hs__tap_1 TAP_1173 ();
 sky130_as_sc_hs__tap_1 TAP_1174 ();
 sky130_as_sc_hs__tap_1 TAP_1175 ();
 sky130_as_sc_hs__tap_1 TAP_1176 ();
 sky130_as_sc_hs__tap_1 TAP_1177 ();
 sky130_as_sc_hs__tap_1 TAP_1178 ();
 sky130_as_sc_hs__tap_1 TAP_1179 ();
 sky130_as_sc_hs__tap_1 TAP_1180 ();
 sky130_as_sc_hs__tap_1 TAP_1181 ();
 sky130_as_sc_hs__tap_1 TAP_1182 ();
 sky130_as_sc_hs__tap_1 TAP_1183 ();
 sky130_as_sc_hs__tap_1 TAP_1184 ();
 sky130_as_sc_hs__tap_1 TAP_1185 ();
 sky130_as_sc_hs__tap_1 TAP_1186 ();
 sky130_as_sc_hs__tap_1 TAP_1187 ();
 sky130_as_sc_hs__tap_1 TAP_1188 ();
 sky130_as_sc_hs__tap_1 TAP_1189 ();
 sky130_as_sc_hs__tap_1 TAP_1190 ();
 sky130_as_sc_hs__tap_1 TAP_1191 ();
 sky130_as_sc_hs__tap_1 TAP_1192 ();
 sky130_as_sc_hs__tap_1 TAP_1193 ();
 sky130_as_sc_hs__tap_1 TAP_1194 ();
 sky130_as_sc_hs__tap_1 TAP_1195 ();
 sky130_as_sc_hs__tap_1 TAP_1196 ();
 sky130_as_sc_hs__tap_1 TAP_1197 ();
 sky130_as_sc_hs__tap_1 TAP_1198 ();
 sky130_as_sc_hs__tap_1 TAP_1199 ();
 sky130_as_sc_hs__tap_1 TAP_1200 ();
 sky130_as_sc_hs__tap_1 TAP_1201 ();
 sky130_as_sc_hs__tap_1 TAP_1202 ();
 sky130_as_sc_hs__tap_1 TAP_1203 ();
 sky130_as_sc_hs__tap_1 TAP_1204 ();
 sky130_as_sc_hs__tap_1 TAP_1205 ();
 sky130_as_sc_hs__tap_1 TAP_1206 ();
 sky130_as_sc_hs__tap_1 TAP_1207 ();
 sky130_as_sc_hs__tap_1 TAP_1208 ();
 sky130_as_sc_hs__tap_1 TAP_1209 ();
 sky130_as_sc_hs__tap_1 TAP_1210 ();
 sky130_as_sc_hs__tap_1 TAP_1211 ();
 sky130_as_sc_hs__tap_1 TAP_1212 ();
 sky130_as_sc_hs__tap_1 TAP_1213 ();
 sky130_as_sc_hs__tap_1 TAP_1214 ();
 sky130_as_sc_hs__tap_1 TAP_1215 ();
 sky130_as_sc_hs__tap_1 TAP_1216 ();
 sky130_as_sc_hs__tap_1 TAP_1217 ();
 sky130_as_sc_hs__tap_1 TAP_1218 ();
 sky130_as_sc_hs__tap_1 TAP_1219 ();
 sky130_as_sc_hs__tap_1 TAP_1220 ();
 sky130_as_sc_hs__tap_1 TAP_1221 ();
 sky130_as_sc_hs__tap_1 TAP_1222 ();
 sky130_as_sc_hs__tap_1 TAP_1223 ();
 sky130_as_sc_hs__tap_1 TAP_1224 ();
 sky130_as_sc_hs__tap_1 TAP_1225 ();
 sky130_as_sc_hs__tap_1 TAP_1226 ();
 sky130_as_sc_hs__tap_1 TAP_1227 ();
 sky130_as_sc_hs__tap_1 TAP_1228 ();
 sky130_as_sc_hs__tap_1 TAP_1229 ();
 sky130_as_sc_hs__tap_1 TAP_1230 ();
 sky130_as_sc_hs__tap_1 TAP_1231 ();
 sky130_as_sc_hs__tap_1 TAP_1232 ();
 sky130_as_sc_hs__tap_1 TAP_1233 ();
 sky130_as_sc_hs__tap_1 TAP_1234 ();
 sky130_as_sc_hs__tap_1 TAP_1235 ();
 sky130_as_sc_hs__tap_1 TAP_1236 ();
 sky130_as_sc_hs__tap_1 TAP_1237 ();
 sky130_as_sc_hs__tap_1 TAP_1238 ();
 sky130_as_sc_hs__tap_1 TAP_1239 ();
 sky130_as_sc_hs__tap_1 TAP_1240 ();
 sky130_as_sc_hs__tap_1 TAP_1241 ();
 sky130_as_sc_hs__tap_1 TAP_1242 ();
 sky130_as_sc_hs__tap_1 TAP_1243 ();
 sky130_as_sc_hs__tap_1 TAP_1244 ();
 sky130_as_sc_hs__tap_1 TAP_1245 ();
 sky130_as_sc_hs__tap_1 TAP_1246 ();
 sky130_as_sc_hs__tap_1 TAP_1247 ();
 sky130_as_sc_hs__tap_1 TAP_1248 ();
 sky130_as_sc_hs__tap_1 TAP_1249 ();
 sky130_as_sc_hs__tap_1 TAP_1250 ();
 sky130_as_sc_hs__tap_1 TAP_1251 ();
 sky130_as_sc_hs__tap_1 TAP_1252 ();
 sky130_as_sc_hs__tap_1 TAP_1253 ();
 sky130_as_sc_hs__tap_1 TAP_1254 ();
 sky130_as_sc_hs__tap_1 TAP_1255 ();
 sky130_as_sc_hs__tap_1 TAP_1256 ();
 sky130_as_sc_hs__tap_1 TAP_1257 ();
 sky130_as_sc_hs__tap_1 TAP_1258 ();
 sky130_as_sc_hs__tap_1 TAP_1259 ();
 sky130_as_sc_hs__tap_1 TAP_1260 ();
 sky130_as_sc_hs__tap_1 TAP_1261 ();
 sky130_as_sc_hs__tap_1 TAP_1262 ();
 sky130_as_sc_hs__tap_1 TAP_1263 ();
 sky130_as_sc_hs__tap_1 TAP_1264 ();
 sky130_as_sc_hs__tap_1 TAP_1265 ();
 sky130_as_sc_hs__tap_1 TAP_1266 ();
 sky130_as_sc_hs__tap_1 TAP_1267 ();
 sky130_as_sc_hs__tap_1 TAP_1268 ();
 sky130_as_sc_hs__tap_1 TAP_1269 ();
 sky130_as_sc_hs__tap_1 TAP_1270 ();
 sky130_as_sc_hs__tap_1 TAP_1271 ();
 sky130_as_sc_hs__tap_1 TAP_1272 ();
 sky130_as_sc_hs__tap_1 TAP_1273 ();
 sky130_as_sc_hs__tap_1 TAP_1274 ();
 sky130_as_sc_hs__tap_1 TAP_1275 ();
 sky130_as_sc_hs__tap_1 TAP_1276 ();
 sky130_as_sc_hs__tap_1 TAP_1277 ();
 sky130_as_sc_hs__tap_1 TAP_1278 ();
 sky130_as_sc_hs__tap_1 TAP_1279 ();
 sky130_as_sc_hs__tap_1 TAP_1280 ();
 sky130_as_sc_hs__tap_1 TAP_1281 ();
 sky130_as_sc_hs__tap_1 TAP_1282 ();
 sky130_as_sc_hs__tap_1 TAP_1283 ();
 sky130_as_sc_hs__tap_1 TAP_1284 ();
 sky130_as_sc_hs__tap_1 TAP_1285 ();
 sky130_as_sc_hs__tap_1 TAP_1286 ();
 sky130_as_sc_hs__tap_1 TAP_1287 ();
 sky130_as_sc_hs__tap_1 TAP_1288 ();
 sky130_as_sc_hs__tap_1 TAP_1289 ();
 sky130_as_sc_hs__tap_1 TAP_1290 ();
 sky130_as_sc_hs__tap_1 TAP_1291 ();
 sky130_as_sc_hs__tap_1 TAP_1292 ();
 sky130_as_sc_hs__tap_1 TAP_1293 ();
 sky130_as_sc_hs__tap_1 TAP_1294 ();
 sky130_as_sc_hs__tap_1 TAP_1295 ();
 sky130_as_sc_hs__tap_1 TAP_1296 ();
 sky130_as_sc_hs__tap_1 TAP_1297 ();
 sky130_as_sc_hs__tap_1 TAP_1298 ();
 sky130_as_sc_hs__tap_1 TAP_1299 ();
 sky130_as_sc_hs__tap_1 TAP_1300 ();
 sky130_as_sc_hs__tap_1 TAP_1301 ();
 sky130_as_sc_hs__tap_1 TAP_1302 ();
 sky130_as_sc_hs__tap_1 TAP_1303 ();
 sky130_as_sc_hs__tap_1 TAP_1304 ();
 sky130_as_sc_hs__tap_1 TAP_1305 ();
 sky130_as_sc_hs__tap_1 TAP_1306 ();
 sky130_as_sc_hs__tap_1 TAP_1307 ();
 sky130_as_sc_hs__tap_1 TAP_1308 ();
 sky130_as_sc_hs__tap_1 TAP_1309 ();
 sky130_as_sc_hs__tap_1 TAP_1310 ();
 sky130_as_sc_hs__tap_1 TAP_1311 ();
 sky130_as_sc_hs__tap_1 TAP_1312 ();
 sky130_as_sc_hs__tap_1 TAP_1313 ();
 sky130_as_sc_hs__tap_1 TAP_1314 ();
 sky130_as_sc_hs__tap_1 TAP_1315 ();
 sky130_as_sc_hs__tap_1 TAP_1316 ();
 sky130_as_sc_hs__tap_1 TAP_1317 ();
 sky130_as_sc_hs__tap_1 TAP_1318 ();
 sky130_as_sc_hs__tap_1 TAP_1319 ();
 sky130_as_sc_hs__tap_1 TAP_1320 ();
 sky130_as_sc_hs__tap_1 TAP_1321 ();
 sky130_as_sc_hs__tap_1 TAP_1322 ();
 sky130_as_sc_hs__tap_1 TAP_1323 ();
 sky130_as_sc_hs__tap_1 TAP_1324 ();
 sky130_as_sc_hs__tap_1 TAP_1325 ();
 sky130_as_sc_hs__tap_1 TAP_1326 ();
 sky130_as_sc_hs__tap_1 TAP_1327 ();
 sky130_as_sc_hs__tap_1 TAP_1328 ();
 sky130_as_sc_hs__tap_1 TAP_1329 ();
 sky130_as_sc_hs__tap_1 TAP_1330 ();
 sky130_as_sc_hs__tap_1 TAP_1331 ();
 sky130_as_sc_hs__tap_1 TAP_1332 ();
 sky130_as_sc_hs__tap_1 TAP_1333 ();
 sky130_as_sc_hs__tap_1 TAP_1334 ();
 sky130_as_sc_hs__tap_1 TAP_1335 ();
 sky130_as_sc_hs__tap_1 TAP_1336 ();
 sky130_as_sc_hs__tap_1 TAP_1337 ();
 sky130_as_sc_hs__tap_1 TAP_1338 ();
 sky130_as_sc_hs__tap_1 TAP_1339 ();
 sky130_as_sc_hs__tap_1 TAP_1340 ();
 sky130_as_sc_hs__tap_1 TAP_1341 ();
 sky130_as_sc_hs__tap_1 TAP_1342 ();
 sky130_as_sc_hs__tap_1 TAP_1343 ();
 sky130_as_sc_hs__tap_1 TAP_1344 ();
 sky130_as_sc_hs__tap_1 TAP_1345 ();
 sky130_as_sc_hs__tap_1 TAP_1346 ();
 sky130_as_sc_hs__tap_1 TAP_1347 ();
 sky130_as_sc_hs__tap_1 TAP_1348 ();
 sky130_as_sc_hs__tap_1 TAP_1349 ();
 sky130_as_sc_hs__tap_1 TAP_1350 ();
 sky130_as_sc_hs__tap_1 TAP_1351 ();
 sky130_as_sc_hs__tap_1 TAP_1352 ();
 sky130_as_sc_hs__tap_1 TAP_1353 ();
 sky130_as_sc_hs__tap_1 TAP_1354 ();
 sky130_as_sc_hs__tap_1 TAP_1355 ();
 sky130_as_sc_hs__tap_1 TAP_1356 ();
 sky130_as_sc_hs__tap_1 TAP_1357 ();
 sky130_as_sc_hs__tap_1 TAP_1358 ();
 sky130_as_sc_hs__tap_1 TAP_1359 ();
 sky130_as_sc_hs__tap_1 TAP_1360 ();
 sky130_as_sc_hs__tap_1 TAP_1361 ();
 sky130_as_sc_hs__tap_1 TAP_1362 ();
 sky130_as_sc_hs__tap_1 TAP_1363 ();
 sky130_as_sc_hs__tap_1 TAP_1364 ();
 sky130_as_sc_hs__tap_1 TAP_1365 ();
 sky130_as_sc_hs__tap_1 TAP_1366 ();
 sky130_as_sc_hs__tap_1 TAP_1367 ();
 sky130_as_sc_hs__tap_1 TAP_1368 ();
 sky130_as_sc_hs__tap_1 TAP_1369 ();
 sky130_as_sc_hs__tap_1 TAP_1370 ();
 sky130_as_sc_hs__tap_1 TAP_1371 ();
 sky130_as_sc_hs__tap_1 TAP_1372 ();
 sky130_as_sc_hs__tap_1 TAP_1373 ();
 sky130_as_sc_hs__tap_1 TAP_1374 ();
 sky130_as_sc_hs__tap_1 TAP_1375 ();
 sky130_as_sc_hs__tap_1 TAP_1376 ();
 sky130_as_sc_hs__tap_1 TAP_1377 ();
 sky130_as_sc_hs__tap_1 TAP_1378 ();
 sky130_as_sc_hs__tap_1 TAP_1379 ();
 sky130_as_sc_hs__tap_1 TAP_1380 ();
 sky130_as_sc_hs__tap_1 TAP_1381 ();
 sky130_as_sc_hs__tap_1 TAP_1382 ();
 sky130_as_sc_hs__tap_1 TAP_1383 ();
 sky130_as_sc_hs__tap_1 TAP_1384 ();
 sky130_as_sc_hs__tap_1 TAP_1385 ();
 sky130_as_sc_hs__tap_1 TAP_1386 ();
 sky130_as_sc_hs__tap_1 TAP_1387 ();
 sky130_as_sc_hs__tap_1 TAP_1388 ();
 sky130_as_sc_hs__tap_1 TAP_1389 ();
 sky130_as_sc_hs__tap_1 TAP_1390 ();
 sky130_as_sc_hs__tap_1 TAP_1391 ();
 sky130_as_sc_hs__tap_1 TAP_1392 ();
 sky130_as_sc_hs__tap_1 TAP_1393 ();
 sky130_as_sc_hs__tap_1 TAP_1394 ();
 sky130_as_sc_hs__tap_1 TAP_1395 ();
 sky130_as_sc_hs__tap_1 TAP_1396 ();
 sky130_as_sc_hs__tap_1 TAP_1397 ();
 sky130_as_sc_hs__tap_1 TAP_1398 ();
 sky130_as_sc_hs__tap_1 TAP_1399 ();
 sky130_as_sc_hs__tap_1 TAP_1400 ();
 sky130_as_sc_hs__tap_1 TAP_1401 ();
 sky130_as_sc_hs__tap_1 TAP_1402 ();
 sky130_as_sc_hs__tap_1 TAP_1403 ();
 sky130_as_sc_hs__tap_1 TAP_1404 ();
 sky130_as_sc_hs__tap_1 TAP_1405 ();
 sky130_as_sc_hs__tap_1 TAP_1406 ();
 sky130_as_sc_hs__tap_1 TAP_1407 ();
 sky130_as_sc_hs__tap_1 TAP_1408 ();
 sky130_as_sc_hs__tap_1 TAP_1409 ();
 sky130_as_sc_hs__tap_1 TAP_1410 ();
 sky130_as_sc_hs__tap_1 TAP_1411 ();
 sky130_as_sc_hs__tap_1 TAP_1412 ();
 sky130_as_sc_hs__tap_1 TAP_1413 ();
 sky130_as_sc_hs__tap_1 TAP_1414 ();
 sky130_as_sc_hs__tap_1 TAP_1415 ();
 sky130_as_sc_hs__tap_1 TAP_1416 ();
 sky130_as_sc_hs__tap_1 TAP_1417 ();
 sky130_as_sc_hs__tap_1 TAP_1418 ();
 sky130_as_sc_hs__tap_1 TAP_1419 ();
 sky130_as_sc_hs__tap_1 TAP_1420 ();
 sky130_as_sc_hs__tap_1 TAP_1421 ();
 sky130_as_sc_hs__tap_1 TAP_1422 ();
 sky130_as_sc_hs__tap_1 TAP_1423 ();
 sky130_as_sc_hs__tap_1 TAP_1424 ();
 sky130_as_sc_hs__tap_1 TAP_1425 ();
 sky130_as_sc_hs__tap_1 TAP_1426 ();
 sky130_as_sc_hs__tap_1 TAP_1427 ();
 sky130_as_sc_hs__tap_1 TAP_1428 ();
 sky130_as_sc_hs__tap_1 TAP_1429 ();
 sky130_as_sc_hs__tap_1 TAP_1430 ();
 sky130_as_sc_hs__tap_1 TAP_1431 ();
 sky130_as_sc_hs__tap_1 TAP_1432 ();
 sky130_as_sc_hs__tap_1 TAP_1433 ();
 sky130_as_sc_hs__tap_1 TAP_1434 ();
 sky130_as_sc_hs__tap_1 TAP_1435 ();
 sky130_as_sc_hs__tap_1 TAP_1436 ();
 sky130_as_sc_hs__tap_1 TAP_1437 ();
 sky130_as_sc_hs__tap_1 TAP_1438 ();
 sky130_as_sc_hs__tap_1 TAP_1439 ();
 sky130_as_sc_hs__tap_1 TAP_1440 ();
 sky130_as_sc_hs__tap_1 TAP_1441 ();
 sky130_as_sc_hs__tap_1 TAP_1442 ();
 sky130_as_sc_hs__tap_1 TAP_1443 ();
 sky130_as_sc_hs__tap_1 TAP_1444 ();
 sky130_as_sc_hs__tap_1 TAP_1445 ();
 sky130_as_sc_hs__tap_1 TAP_1446 ();
 sky130_as_sc_hs__tap_1 TAP_1447 ();
 sky130_as_sc_hs__tap_1 TAP_1448 ();
 sky130_as_sc_hs__tap_1 TAP_1449 ();
 sky130_as_sc_hs__tap_1 TAP_1450 ();
 sky130_as_sc_hs__tap_1 TAP_1451 ();
 sky130_as_sc_hs__tap_1 TAP_1452 ();
 sky130_as_sc_hs__tap_1 TAP_1453 ();
 sky130_as_sc_hs__tap_1 TAP_1454 ();
 sky130_as_sc_hs__tap_1 TAP_1455 ();
 sky130_as_sc_hs__tap_1 TAP_1456 ();
 sky130_as_sc_hs__tap_1 TAP_1457 ();
 sky130_as_sc_hs__tap_1 TAP_1458 ();
 sky130_as_sc_hs__tap_1 TAP_1459 ();
 sky130_as_sc_hs__tap_1 TAP_1460 ();
 sky130_as_sc_hs__tap_1 TAP_1461 ();
 sky130_as_sc_hs__tap_1 TAP_1462 ();
 sky130_as_sc_hs__tap_1 TAP_1463 ();
 sky130_as_sc_hs__tap_1 TAP_1464 ();
 sky130_as_sc_hs__tap_1 TAP_1465 ();
 sky130_as_sc_hs__tap_1 TAP_1466 ();
 sky130_as_sc_hs__tap_1 TAP_1467 ();
 sky130_as_sc_hs__tap_1 TAP_1468 ();
 sky130_as_sc_hs__tap_1 TAP_1469 ();
 sky130_as_sc_hs__tap_1 TAP_1470 ();
 sky130_as_sc_hs__tap_1 TAP_1471 ();
 sky130_as_sc_hs__tap_1 TAP_1472 ();
 sky130_as_sc_hs__tap_1 TAP_1473 ();
 sky130_as_sc_hs__tap_1 TAP_1474 ();
 sky130_as_sc_hs__tap_1 TAP_1475 ();
 sky130_as_sc_hs__tap_1 TAP_1476 ();
 sky130_as_sc_hs__tap_1 TAP_1477 ();
 sky130_as_sc_hs__tap_1 TAP_1478 ();
 sky130_as_sc_hs__tap_1 TAP_1479 ();
 sky130_as_sc_hs__tap_1 TAP_1480 ();
 sky130_as_sc_hs__tap_1 TAP_1481 ();
 sky130_as_sc_hs__tap_1 TAP_1482 ();
 sky130_as_sc_hs__tap_1 TAP_1483 ();
 sky130_as_sc_hs__tap_1 TAP_1484 ();
 sky130_as_sc_hs__tap_1 TAP_1485 ();
 sky130_as_sc_hs__tap_1 TAP_1486 ();
 sky130_as_sc_hs__tap_1 TAP_1487 ();
 sky130_as_sc_hs__tap_1 TAP_1488 ();
 sky130_as_sc_hs__tap_1 TAP_1489 ();
 sky130_as_sc_hs__tap_1 TAP_1490 ();
 sky130_as_sc_hs__tap_1 TAP_1491 ();
 sky130_as_sc_hs__tap_1 TAP_1492 ();
 sky130_as_sc_hs__tap_1 TAP_1493 ();
 sky130_as_sc_hs__tap_1 TAP_1494 ();
 sky130_as_sc_hs__tap_1 TAP_1495 ();
 sky130_as_sc_hs__tap_1 TAP_1496 ();
 sky130_as_sc_hs__tap_1 TAP_1497 ();
 sky130_as_sc_hs__tap_1 TAP_1498 ();
 sky130_as_sc_hs__tap_1 TAP_1499 ();
 sky130_as_sc_hs__tap_1 TAP_1500 ();
 sky130_as_sc_hs__tap_1 TAP_1501 ();
 sky130_as_sc_hs__tap_1 TAP_1502 ();
 sky130_as_sc_hs__tap_1 TAP_1503 ();
 sky130_as_sc_hs__tap_1 TAP_1504 ();
 sky130_as_sc_hs__tap_1 TAP_1505 ();
 sky130_as_sc_hs__tap_1 TAP_1506 ();
 sky130_as_sc_hs__tap_1 TAP_1507 ();
 sky130_as_sc_hs__tap_1 TAP_1508 ();
 sky130_as_sc_hs__tap_1 TAP_1509 ();
 sky130_as_sc_hs__tap_1 TAP_1510 ();
 sky130_as_sc_hs__tap_1 TAP_1511 ();
 sky130_as_sc_hs__tap_1 TAP_1512 ();
 sky130_as_sc_hs__tap_1 TAP_1513 ();
 sky130_as_sc_hs__tap_1 TAP_1514 ();
 sky130_as_sc_hs__tap_1 TAP_1515 ();
 sky130_as_sc_hs__tap_1 TAP_1516 ();
 sky130_as_sc_hs__tap_1 TAP_1517 ();
 sky130_as_sc_hs__tap_1 TAP_1518 ();
 sky130_as_sc_hs__tap_1 TAP_1519 ();
 sky130_as_sc_hs__tap_1 TAP_1520 ();
 sky130_as_sc_hs__tap_1 TAP_1521 ();
 sky130_as_sc_hs__tap_1 TAP_1522 ();
 sky130_as_sc_hs__tap_1 TAP_1523 ();
 sky130_as_sc_hs__tap_1 TAP_1524 ();
 sky130_as_sc_hs__tap_1 TAP_1525 ();
 sky130_as_sc_hs__tap_1 TAP_1526 ();
 sky130_as_sc_hs__tap_1 TAP_1527 ();
 sky130_as_sc_hs__tap_1 TAP_1528 ();
 sky130_as_sc_hs__tap_1 TAP_1529 ();
 sky130_as_sc_hs__tap_1 TAP_1530 ();
 sky130_as_sc_hs__tap_1 TAP_1531 ();
 sky130_as_sc_hs__tap_1 TAP_1532 ();
 sky130_as_sc_hs__tap_1 TAP_1533 ();
 sky130_as_sc_hs__tap_1 TAP_1534 ();
 sky130_as_sc_hs__tap_1 TAP_1535 ();
 sky130_as_sc_hs__tap_1 TAP_1536 ();
 sky130_as_sc_hs__tap_1 TAP_1537 ();
 sky130_as_sc_hs__tap_1 TAP_1538 ();
 sky130_as_sc_hs__tap_1 TAP_1539 ();
 sky130_as_sc_hs__tap_1 TAP_1540 ();
 sky130_as_sc_hs__tap_1 TAP_1541 ();
 sky130_as_sc_hs__tap_1 TAP_1542 ();
 sky130_as_sc_hs__tap_1 TAP_1543 ();
 sky130_as_sc_hs__tap_1 TAP_1544 ();
 sky130_as_sc_hs__tap_1 TAP_1545 ();
 sky130_as_sc_hs__tap_1 TAP_1546 ();
 sky130_as_sc_hs__tap_1 TAP_1547 ();
 sky130_as_sc_hs__tap_1 TAP_1548 ();
 sky130_as_sc_hs__tap_1 TAP_1549 ();
 sky130_as_sc_hs__tap_1 TAP_1550 ();
 sky130_as_sc_hs__tap_1 TAP_1551 ();
 sky130_as_sc_hs__tap_1 TAP_1552 ();
 sky130_as_sc_hs__tap_1 TAP_1553 ();
 sky130_as_sc_hs__tap_1 TAP_1554 ();
 sky130_as_sc_hs__tap_1 TAP_1555 ();
 sky130_as_sc_hs__tap_1 TAP_1556 ();
 sky130_as_sc_hs__tap_1 TAP_1557 ();
 sky130_as_sc_hs__tap_1 TAP_1558 ();
 sky130_as_sc_hs__tap_1 TAP_1559 ();
 sky130_as_sc_hs__tap_1 TAP_1560 ();
 sky130_as_sc_hs__tap_1 TAP_1561 ();
 sky130_as_sc_hs__tap_1 TAP_1562 ();
 sky130_as_sc_hs__tap_1 TAP_1563 ();
 sky130_as_sc_hs__tap_1 TAP_1564 ();
 sky130_as_sc_hs__tap_1 TAP_1565 ();
 sky130_as_sc_hs__tap_1 TAP_1566 ();
 sky130_as_sc_hs__tap_1 TAP_1567 ();
 sky130_as_sc_hs__tap_1 TAP_1568 ();
 sky130_as_sc_hs__tap_1 TAP_1569 ();
 sky130_as_sc_hs__tap_1 TAP_1570 ();
 sky130_as_sc_hs__tap_1 TAP_1571 ();
 sky130_as_sc_hs__tap_1 TAP_1572 ();
 sky130_as_sc_hs__tap_1 TAP_1573 ();
 sky130_as_sc_hs__tap_1 TAP_1574 ();
 sky130_as_sc_hs__tap_1 TAP_1575 ();
 sky130_as_sc_hs__tap_1 TAP_1576 ();
 sky130_as_sc_hs__tap_1 TAP_1577 ();
 sky130_as_sc_hs__tap_1 TAP_1578 ();
 sky130_as_sc_hs__tap_1 TAP_1579 ();
 sky130_as_sc_hs__tap_1 TAP_1580 ();
 sky130_as_sc_hs__tap_1 TAP_1581 ();
 sky130_as_sc_hs__tap_1 TAP_1582 ();
 sky130_as_sc_hs__tap_1 TAP_1583 ();
 sky130_as_sc_hs__tap_1 TAP_1584 ();
 sky130_as_sc_hs__tap_1 TAP_1585 ();
 sky130_as_sc_hs__tap_1 TAP_1586 ();
 sky130_as_sc_hs__tap_1 TAP_1587 ();
 sky130_as_sc_hs__tap_1 TAP_1588 ();
 sky130_as_sc_hs__tap_1 TAP_1589 ();
 sky130_as_sc_hs__tap_1 TAP_1590 ();
 sky130_as_sc_hs__tap_1 TAP_1591 ();
 sky130_as_sc_hs__tap_1 TAP_1592 ();
 sky130_as_sc_hs__tap_1 TAP_1593 ();
 sky130_as_sc_hs__tap_1 TAP_1594 ();
 sky130_as_sc_hs__tap_1 TAP_1595 ();
 sky130_as_sc_hs__tap_1 TAP_1596 ();
 sky130_as_sc_hs__tap_1 TAP_1597 ();
 sky130_as_sc_hs__tap_1 TAP_1598 ();
 sky130_as_sc_hs__tap_1 TAP_1599 ();
 sky130_as_sc_hs__tap_1 TAP_1600 ();
 sky130_as_sc_hs__tap_1 TAP_1601 ();
 sky130_as_sc_hs__tap_1 TAP_1602 ();
 sky130_as_sc_hs__tap_1 TAP_1603 ();
 sky130_as_sc_hs__tap_1 TAP_1604 ();
 sky130_as_sc_hs__tap_1 TAP_1605 ();
 sky130_as_sc_hs__tap_1 TAP_1606 ();
 sky130_as_sc_hs__tap_1 TAP_1607 ();
 sky130_as_sc_hs__tap_1 TAP_1608 ();
 sky130_as_sc_hs__tap_1 TAP_1609 ();
 sky130_as_sc_hs__tap_1 TAP_1610 ();
 sky130_as_sc_hs__tap_1 TAP_1611 ();
 sky130_as_sc_hs__tap_1 TAP_1612 ();
 sky130_as_sc_hs__tap_1 TAP_1613 ();
 sky130_as_sc_hs__tap_1 TAP_1614 ();
 sky130_as_sc_hs__tap_1 TAP_1615 ();
 sky130_as_sc_hs__tap_1 TAP_1616 ();
 sky130_as_sc_hs__tap_1 TAP_1617 ();
 sky130_as_sc_hs__tap_1 TAP_1618 ();
 sky130_as_sc_hs__tap_1 TAP_1619 ();
 sky130_as_sc_hs__tap_1 TAP_1620 ();
 sky130_as_sc_hs__tap_1 TAP_1621 ();
 sky130_as_sc_hs__tap_1 TAP_1622 ();
 sky130_as_sc_hs__tap_1 TAP_1623 ();
 sky130_as_sc_hs__tap_1 TAP_1624 ();
 sky130_as_sc_hs__tap_1 TAP_1625 ();
 sky130_as_sc_hs__tap_1 TAP_1626 ();
 sky130_as_sc_hs__tap_1 TAP_1627 ();
 sky130_as_sc_hs__tap_1 TAP_1628 ();
 sky130_as_sc_hs__tap_1 TAP_1629 ();
 sky130_as_sc_hs__tap_1 TAP_1630 ();
 sky130_as_sc_hs__tap_1 TAP_1631 ();
 sky130_as_sc_hs__tap_1 TAP_1632 ();
 sky130_as_sc_hs__tap_1 TAP_1633 ();
 sky130_as_sc_hs__tap_1 TAP_1634 ();
 sky130_as_sc_hs__tap_1 TAP_1635 ();
 sky130_as_sc_hs__tap_1 TAP_1636 ();
 sky130_as_sc_hs__tap_1 TAP_1637 ();
 sky130_as_sc_hs__tap_1 TAP_1638 ();
 sky130_as_sc_hs__tap_1 TAP_1639 ();
 sky130_as_sc_hs__tap_1 TAP_1640 ();
 sky130_as_sc_hs__tap_1 TAP_1641 ();
 sky130_as_sc_hs__tap_1 TAP_1642 ();
 sky130_as_sc_hs__tap_1 TAP_1643 ();
 sky130_as_sc_hs__tap_1 TAP_1644 ();
 sky130_as_sc_hs__tap_1 TAP_1645 ();
 sky130_as_sc_hs__tap_1 TAP_1646 ();
 sky130_as_sc_hs__tap_1 TAP_1647 ();
 sky130_as_sc_hs__tap_1 TAP_1648 ();
 sky130_as_sc_hs__tap_1 TAP_1649 ();
 sky130_as_sc_hs__tap_1 TAP_1650 ();
 sky130_as_sc_hs__tap_1 TAP_1651 ();
 sky130_as_sc_hs__tap_1 TAP_1652 ();
 sky130_as_sc_hs__tap_1 TAP_1653 ();
 sky130_as_sc_hs__tap_1 TAP_1654 ();
 sky130_as_sc_hs__tap_1 TAP_1655 ();
 sky130_as_sc_hs__tap_1 TAP_1656 ();
 sky130_as_sc_hs__tap_1 TAP_1657 ();
 sky130_as_sc_hs__tap_1 TAP_1658 ();
 sky130_as_sc_hs__tap_1 TAP_1659 ();
 sky130_as_sc_hs__tap_1 TAP_1660 ();
 sky130_as_sc_hs__tap_1 TAP_1661 ();
 sky130_as_sc_hs__tap_1 TAP_1662 ();
 sky130_as_sc_hs__tap_1 TAP_1663 ();
 sky130_as_sc_hs__tap_1 TAP_1664 ();
 sky130_as_sc_hs__tap_1 TAP_1665 ();
 sky130_as_sc_hs__tap_1 TAP_1666 ();
 sky130_as_sc_hs__tap_1 TAP_1667 ();
 sky130_as_sc_hs__tap_1 TAP_1668 ();
 sky130_as_sc_hs__tap_1 TAP_1669 ();
 sky130_as_sc_hs__tap_1 TAP_1670 ();
 sky130_as_sc_hs__tap_1 TAP_1671 ();
 sky130_as_sc_hs__tap_1 TAP_1672 ();
 sky130_as_sc_hs__tap_1 TAP_1673 ();
 sky130_as_sc_hs__tap_1 TAP_1674 ();
 sky130_as_sc_hs__tap_1 TAP_1675 ();
 sky130_as_sc_hs__tap_1 TAP_1676 ();
 sky130_as_sc_hs__tap_1 TAP_1677 ();
 sky130_as_sc_hs__tap_1 TAP_1678 ();
 sky130_as_sc_hs__tap_1 TAP_1679 ();
 sky130_as_sc_hs__tap_1 TAP_1680 ();
 sky130_as_sc_hs__tap_1 TAP_1681 ();
 sky130_as_sc_hs__tap_1 TAP_1682 ();
 sky130_as_sc_hs__tap_1 TAP_1683 ();
 sky130_as_sc_hs__tap_1 TAP_1684 ();
 sky130_as_sc_hs__tap_1 TAP_1685 ();
 sky130_as_sc_hs__tap_1 TAP_1686 ();
 sky130_as_sc_hs__tap_1 TAP_1687 ();
 sky130_as_sc_hs__tap_1 TAP_1688 ();
 sky130_as_sc_hs__tap_1 TAP_1689 ();
 sky130_as_sc_hs__tap_1 TAP_1690 ();
 sky130_as_sc_hs__tap_1 TAP_1691 ();
 sky130_as_sc_hs__tap_1 TAP_1692 ();
 sky130_as_sc_hs__tap_1 TAP_1693 ();
 sky130_as_sc_hs__tap_1 TAP_1694 ();
 sky130_as_sc_hs__tap_1 TAP_1695 ();
 sky130_as_sc_hs__tap_1 TAP_1696 ();
 sky130_as_sc_hs__tap_1 TAP_1697 ();
 sky130_as_sc_hs__tap_1 TAP_1698 ();
 sky130_as_sc_hs__tap_1 TAP_1699 ();
 sky130_as_sc_hs__tap_1 TAP_1700 ();
 sky130_as_sc_hs__tap_1 TAP_1701 ();
 sky130_as_sc_hs__tap_1 TAP_1702 ();
 sky130_as_sc_hs__tap_1 TAP_1703 ();
 sky130_as_sc_hs__tap_1 TAP_1704 ();
 sky130_as_sc_hs__tap_1 TAP_1705 ();
 sky130_as_sc_hs__tap_1 TAP_1706 ();
 sky130_as_sc_hs__tap_1 TAP_1707 ();
 sky130_as_sc_hs__tap_1 TAP_1708 ();
 sky130_as_sc_hs__tap_1 TAP_1709 ();
 sky130_as_sc_hs__tap_1 TAP_1710 ();
 sky130_as_sc_hs__tap_1 TAP_1711 ();
 sky130_as_sc_hs__tap_1 TAP_1712 ();
 sky130_as_sc_hs__tap_1 TAP_1713 ();
 sky130_as_sc_hs__tap_1 TAP_1714 ();
 sky130_as_sc_hs__tap_1 TAP_1715 ();
 sky130_as_sc_hs__tap_1 TAP_1716 ();
 sky130_as_sc_hs__tap_1 TAP_1717 ();
 sky130_as_sc_hs__tap_1 TAP_1718 ();
 sky130_as_sc_hs__tap_1 TAP_1719 ();
 sky130_as_sc_hs__tap_1 TAP_1720 ();
 sky130_as_sc_hs__tap_1 TAP_1721 ();
 sky130_as_sc_hs__tap_1 TAP_1722 ();
 sky130_as_sc_hs__tap_1 TAP_1723 ();
 sky130_as_sc_hs__tap_1 TAP_1724 ();
 sky130_as_sc_hs__tap_1 TAP_1725 ();
 sky130_as_sc_hs__tap_1 TAP_1726 ();
 sky130_as_sc_hs__tap_1 TAP_1727 ();
 sky130_as_sc_hs__tap_1 TAP_1728 ();
 sky130_as_sc_hs__tap_1 TAP_1729 ();
 sky130_as_sc_hs__tap_1 TAP_1730 ();
 sky130_as_sc_hs__tap_1 TAP_1731 ();
 sky130_as_sc_hs__tap_1 TAP_1732 ();
 sky130_as_sc_hs__tap_1 TAP_1733 ();
 sky130_as_sc_hs__tap_1 TAP_1734 ();
 sky130_as_sc_hs__tap_1 TAP_1735 ();
 sky130_as_sc_hs__tap_1 TAP_1736 ();
 sky130_as_sc_hs__tap_1 TAP_1737 ();
 sky130_as_sc_hs__tap_1 TAP_1738 ();
 sky130_as_sc_hs__tap_1 TAP_1739 ();
 sky130_as_sc_hs__tap_1 TAP_1740 ();
 sky130_as_sc_hs__tap_1 TAP_1741 ();
 sky130_as_sc_hs__tap_1 TAP_1742 ();
 sky130_as_sc_hs__tap_1 TAP_1743 ();
 sky130_as_sc_hs__tap_1 TAP_1744 ();
 sky130_as_sc_hs__tap_1 TAP_1745 ();
 sky130_as_sc_hs__tap_1 TAP_1746 ();
 sky130_as_sc_hs__tap_1 TAP_1747 ();
 sky130_as_sc_hs__tap_1 TAP_1748 ();
 sky130_as_sc_hs__tap_1 TAP_1749 ();
 sky130_as_sc_hs__tap_1 TAP_1750 ();
 sky130_as_sc_hs__tap_1 TAP_1751 ();
 sky130_as_sc_hs__tap_1 TAP_1752 ();
 sky130_as_sc_hs__tap_1 TAP_1753 ();
 sky130_as_sc_hs__tap_1 TAP_1754 ();
 sky130_as_sc_hs__tap_1 TAP_1755 ();
 sky130_as_sc_hs__tap_1 TAP_1756 ();
 sky130_as_sc_hs__tap_1 TAP_1757 ();
 sky130_as_sc_hs__tap_1 TAP_1758 ();
 sky130_as_sc_hs__tap_1 TAP_1759 ();
 sky130_as_sc_hs__tap_1 TAP_1760 ();
 sky130_as_sc_hs__tap_1 TAP_1761 ();
 sky130_as_sc_hs__tap_1 TAP_1762 ();
 sky130_as_sc_hs__tap_1 TAP_1763 ();
 sky130_as_sc_hs__tap_1 TAP_1764 ();
 sky130_as_sc_hs__tap_1 TAP_1765 ();
 sky130_as_sc_hs__tap_1 TAP_1766 ();
 sky130_as_sc_hs__tap_1 TAP_1767 ();
 sky130_as_sc_hs__tap_1 TAP_1768 ();
 sky130_as_sc_hs__tap_1 TAP_1769 ();
 sky130_as_sc_hs__tap_1 TAP_1770 ();
 sky130_as_sc_hs__tap_1 TAP_1771 ();
 sky130_as_sc_hs__tap_1 TAP_1772 ();
 sky130_as_sc_hs__tap_1 TAP_1773 ();
 sky130_as_sc_hs__tap_1 TAP_1774 ();
 sky130_as_sc_hs__tap_1 TAP_1775 ();
 sky130_as_sc_hs__tap_1 TAP_1776 ();
 sky130_as_sc_hs__tap_1 TAP_1777 ();
 sky130_as_sc_hs__tap_1 TAP_1778 ();
 sky130_as_sc_hs__tap_1 TAP_1779 ();
 sky130_as_sc_hs__tap_1 TAP_1780 ();
 sky130_as_sc_hs__tap_1 TAP_1781 ();
 sky130_as_sc_hs__tap_1 TAP_1782 ();
 sky130_as_sc_hs__tap_1 TAP_1783 ();
 sky130_as_sc_hs__tap_1 TAP_1784 ();
 sky130_as_sc_hs__tap_1 TAP_1785 ();
 sky130_as_sc_hs__tap_1 TAP_1786 ();
 sky130_as_sc_hs__tap_1 TAP_1787 ();
 sky130_as_sc_hs__tap_1 TAP_1788 ();
 sky130_as_sc_hs__tap_1 TAP_1789 ();
 sky130_as_sc_hs__tap_1 TAP_1790 ();
 sky130_as_sc_hs__tap_1 TAP_1791 ();
 sky130_as_sc_hs__tap_1 TAP_1792 ();
 sky130_as_sc_hs__tap_1 TAP_1793 ();
 sky130_as_sc_hs__tap_1 TAP_1794 ();
 sky130_as_sc_hs__tap_1 TAP_1795 ();
 sky130_as_sc_hs__tap_1 TAP_1796 ();
 sky130_as_sc_hs__tap_1 TAP_1797 ();
 sky130_as_sc_hs__tap_1 TAP_1798 ();
 sky130_as_sc_hs__tap_1 TAP_1799 ();
 sky130_as_sc_hs__tap_1 TAP_1800 ();
 sky130_as_sc_hs__tap_1 TAP_1801 ();
 sky130_as_sc_hs__tap_1 TAP_1802 ();
 sky130_as_sc_hs__tap_1 TAP_1803 ();
 sky130_as_sc_hs__tap_1 TAP_1804 ();
 sky130_as_sc_hs__tap_1 TAP_1805 ();
 sky130_as_sc_hs__tap_1 TAP_1806 ();
 sky130_as_sc_hs__tap_1 TAP_1807 ();
 sky130_as_sc_hs__tap_1 TAP_1808 ();
 sky130_as_sc_hs__tap_1 TAP_1809 ();
 sky130_as_sc_hs__tap_1 TAP_1810 ();
 sky130_as_sc_hs__tap_1 TAP_1811 ();
 sky130_as_sc_hs__tap_1 TAP_1812 ();
 sky130_as_sc_hs__tap_1 TAP_1813 ();
 sky130_as_sc_hs__tap_1 TAP_1814 ();
 sky130_as_sc_hs__tap_1 TAP_1815 ();
 sky130_as_sc_hs__tap_1 TAP_1816 ();
 sky130_as_sc_hs__tap_1 TAP_1817 ();
 sky130_as_sc_hs__tap_1 TAP_1818 ();
 sky130_as_sc_hs__tap_1 TAP_1819 ();
 sky130_as_sc_hs__tap_1 TAP_1820 ();
 sky130_as_sc_hs__tap_1 TAP_1821 ();
 sky130_as_sc_hs__tap_1 TAP_1822 ();
 sky130_as_sc_hs__tap_1 TAP_1823 ();
 sky130_as_sc_hs__tap_1 TAP_1824 ();
 sky130_as_sc_hs__tap_1 TAP_1825 ();
 sky130_as_sc_hs__tap_1 TAP_1826 ();
 sky130_as_sc_hs__tap_1 TAP_1827 ();
 sky130_as_sc_hs__tap_1 TAP_1828 ();
 sky130_as_sc_hs__tap_1 TAP_1829 ();
 sky130_as_sc_hs__tap_1 TAP_1830 ();
 sky130_as_sc_hs__tap_1 TAP_1831 ();
 sky130_as_sc_hs__tap_1 TAP_1832 ();
 sky130_as_sc_hs__tap_1 TAP_1833 ();
 sky130_as_sc_hs__tap_1 TAP_1834 ();
 sky130_as_sc_hs__tap_1 TAP_1835 ();
 sky130_as_sc_hs__tap_1 TAP_1836 ();
 sky130_as_sc_hs__tap_1 TAP_1837 ();
 sky130_as_sc_hs__tap_1 TAP_1838 ();
 sky130_as_sc_hs__tap_1 TAP_1839 ();
 sky130_as_sc_hs__tap_1 TAP_1840 ();
 sky130_as_sc_hs__tap_1 TAP_1841 ();
 sky130_as_sc_hs__tap_1 TAP_1842 ();
 sky130_as_sc_hs__tap_1 TAP_1843 ();
 sky130_as_sc_hs__tap_1 TAP_1844 ();
 sky130_as_sc_hs__tap_1 TAP_1845 ();
 sky130_as_sc_hs__tap_1 TAP_1846 ();
 sky130_as_sc_hs__tap_1 TAP_1847 ();
 sky130_as_sc_hs__tap_1 TAP_1848 ();
 sky130_as_sc_hs__tap_1 TAP_1849 ();
 sky130_as_sc_hs__tap_1 TAP_1850 ();
 sky130_as_sc_hs__tap_1 TAP_1851 ();
 sky130_as_sc_hs__tap_1 TAP_1852 ();
 sky130_as_sc_hs__tap_1 TAP_1853 ();
 sky130_as_sc_hs__tap_1 TAP_1854 ();
 sky130_as_sc_hs__tap_1 TAP_1855 ();
 sky130_as_sc_hs__tap_1 TAP_1856 ();
 sky130_as_sc_hs__tap_1 TAP_1857 ();
 sky130_as_sc_hs__tap_1 TAP_1858 ();
 sky130_as_sc_hs__tap_1 TAP_1859 ();
 sky130_as_sc_hs__tap_1 TAP_1860 ();
 sky130_as_sc_hs__tap_1 TAP_1861 ();
 sky130_as_sc_hs__tap_1 TAP_1862 ();
 sky130_as_sc_hs__tap_1 TAP_1863 ();
 sky130_as_sc_hs__tap_1 TAP_1864 ();
 sky130_as_sc_hs__tap_1 TAP_1865 ();
 sky130_as_sc_hs__tap_1 TAP_1866 ();
 sky130_as_sc_hs__tap_1 TAP_1867 ();
 sky130_as_sc_hs__tap_1 TAP_1868 ();
 sky130_as_sc_hs__tap_1 TAP_1869 ();
 sky130_as_sc_hs__tap_1 TAP_1870 ();
 sky130_as_sc_hs__tap_1 TAP_1871 ();
 sky130_as_sc_hs__tap_1 TAP_1872 ();
 sky130_as_sc_hs__tap_1 TAP_1873 ();
 sky130_as_sc_hs__tap_1 TAP_1874 ();
 sky130_as_sc_hs__tap_1 TAP_1875 ();
 sky130_as_sc_hs__tap_1 TAP_1876 ();
 sky130_as_sc_hs__tap_1 TAP_1877 ();
 sky130_as_sc_hs__tap_1 TAP_1878 ();
 sky130_as_sc_hs__tap_1 TAP_1879 ();
 sky130_as_sc_hs__tap_1 TAP_1880 ();
 sky130_as_sc_hs__tap_1 TAP_1881 ();
 sky130_as_sc_hs__tap_1 TAP_1882 ();
 sky130_as_sc_hs__tap_1 TAP_1883 ();
 sky130_as_sc_hs__tap_1 TAP_1884 ();
 sky130_as_sc_hs__tap_1 TAP_1885 ();
 sky130_as_sc_hs__tap_1 TAP_1886 ();
 sky130_as_sc_hs__tap_1 TAP_1887 ();
 sky130_as_sc_hs__tap_1 TAP_1888 ();
 sky130_as_sc_hs__tap_1 TAP_1889 ();
 sky130_as_sc_hs__tap_1 TAP_1890 ();
 sky130_as_sc_hs__tap_1 TAP_1891 ();
 sky130_as_sc_hs__tap_1 TAP_1892 ();
 sky130_as_sc_hs__tap_1 TAP_1893 ();
 sky130_as_sc_hs__tap_1 TAP_1894 ();
 sky130_as_sc_hs__tap_1 TAP_1895 ();
 sky130_as_sc_hs__tap_1 TAP_1896 ();
 sky130_as_sc_hs__tap_1 TAP_1897 ();
 sky130_as_sc_hs__tap_1 TAP_1898 ();
 sky130_as_sc_hs__tap_1 TAP_1899 ();
 sky130_as_sc_hs__tap_1 TAP_1900 ();
 sky130_as_sc_hs__tap_1 TAP_1901 ();
 sky130_as_sc_hs__tap_1 TAP_1902 ();
 sky130_as_sc_hs__tap_1 TAP_1903 ();
 sky130_as_sc_hs__tap_1 TAP_1904 ();
 sky130_as_sc_hs__tap_1 TAP_1905 ();
 sky130_as_sc_hs__tap_1 TAP_1906 ();
 sky130_as_sc_hs__tap_1 TAP_1907 ();
 sky130_as_sc_hs__tap_1 TAP_1908 ();
 sky130_as_sc_hs__tap_1 TAP_1909 ();
 sky130_as_sc_hs__tap_1 TAP_1910 ();
 sky130_as_sc_hs__tap_1 TAP_1911 ();
 sky130_as_sc_hs__tap_1 TAP_1912 ();
 sky130_as_sc_hs__tap_1 TAP_1913 ();
 sky130_as_sc_hs__tap_1 TAP_1914 ();
 sky130_as_sc_hs__tap_1 TAP_1915 ();
 sky130_as_sc_hs__tap_1 TAP_1916 ();
 sky130_as_sc_hs__tap_1 TAP_1917 ();
 sky130_as_sc_hs__tap_1 TAP_1918 ();
 sky130_as_sc_hs__tap_1 TAP_1919 ();
 sky130_as_sc_hs__tap_1 TAP_1920 ();
 sky130_as_sc_hs__tap_1 TAP_1921 ();
 sky130_as_sc_hs__tap_1 TAP_1922 ();
 sky130_as_sc_hs__tap_1 TAP_1923 ();
 sky130_as_sc_hs__tap_1 TAP_1924 ();
 sky130_as_sc_hs__tap_1 TAP_1925 ();
 sky130_as_sc_hs__tap_1 TAP_1926 ();
 sky130_as_sc_hs__tap_1 TAP_1927 ();
 sky130_as_sc_hs__tap_1 TAP_1928 ();
 sky130_as_sc_hs__tap_1 TAP_1929 ();
 sky130_as_sc_hs__tap_1 TAP_1930 ();
 sky130_as_sc_hs__tap_1 TAP_1931 ();
 sky130_as_sc_hs__tap_1 TAP_1932 ();
 sky130_as_sc_hs__tap_1 TAP_1933 ();
 sky130_as_sc_hs__tap_1 TAP_1934 ();
 sky130_as_sc_hs__tap_1 TAP_1935 ();
 sky130_as_sc_hs__tap_1 TAP_1936 ();
 sky130_as_sc_hs__tap_1 TAP_1937 ();
 sky130_as_sc_hs__tap_1 TAP_1938 ();
 sky130_as_sc_hs__tap_1 TAP_1939 ();
 sky130_as_sc_hs__tap_1 TAP_1940 ();
 sky130_as_sc_hs__tap_1 TAP_1941 ();
 sky130_as_sc_hs__tap_1 TAP_1942 ();
 sky130_as_sc_hs__tap_1 TAP_1943 ();
 sky130_as_sc_hs__tap_1 TAP_1944 ();
 sky130_as_sc_hs__tap_1 TAP_1945 ();
 sky130_as_sc_hs__tap_1 TAP_1946 ();
 sky130_as_sc_hs__tap_1 TAP_1947 ();
 sky130_as_sc_hs__tap_1 TAP_1948 ();
 sky130_as_sc_hs__tap_1 TAP_1949 ();
 sky130_as_sc_hs__tap_1 TAP_1950 ();
 sky130_as_sc_hs__tap_1 TAP_1951 ();
 sky130_as_sc_hs__tap_1 TAP_1952 ();
 sky130_as_sc_hs__tap_1 TAP_1953 ();
 sky130_as_sc_hs__tap_1 TAP_1954 ();
 sky130_as_sc_hs__tap_1 TAP_1955 ();
 sky130_as_sc_hs__tap_1 TAP_1956 ();
 sky130_as_sc_hs__tap_1 TAP_1957 ();
 sky130_as_sc_hs__tap_1 TAP_1958 ();
 sky130_as_sc_hs__tap_1 TAP_1959 ();
 sky130_as_sc_hs__tap_1 TAP_1960 ();
 sky130_as_sc_hs__tap_1 TAP_1961 ();
 sky130_as_sc_hs__tap_1 TAP_1962 ();
 sky130_as_sc_hs__tap_1 TAP_1963 ();
 sky130_as_sc_hs__tap_1 TAP_1964 ();
 sky130_as_sc_hs__tap_1 TAP_1965 ();
 sky130_as_sc_hs__tap_1 TAP_1966 ();
 sky130_as_sc_hs__tap_1 TAP_1967 ();
 sky130_as_sc_hs__tap_1 TAP_1968 ();
 sky130_as_sc_hs__tap_1 TAP_1969 ();
 sky130_as_sc_hs__tap_1 TAP_1970 ();
 sky130_as_sc_hs__tap_1 TAP_1971 ();
 sky130_as_sc_hs__tap_1 TAP_1972 ();
 sky130_as_sc_hs__tap_1 TAP_1973 ();
 sky130_as_sc_hs__tap_1 TAP_1974 ();
 sky130_as_sc_hs__tap_1 TAP_1975 ();
 sky130_as_sc_hs__tap_1 TAP_1976 ();
 sky130_as_sc_hs__tap_1 TAP_1977 ();
 sky130_as_sc_hs__tap_1 TAP_1978 ();
 sky130_as_sc_hs__tap_1 TAP_1979 ();
 sky130_as_sc_hs__tap_1 TAP_1980 ();
 sky130_as_sc_hs__tap_1 TAP_1981 ();
 sky130_as_sc_hs__tap_1 TAP_1982 ();
 sky130_as_sc_hs__tap_1 TAP_1983 ();
 sky130_as_sc_hs__tap_1 TAP_1984 ();
 sky130_as_sc_hs__tap_1 TAP_1985 ();
 sky130_as_sc_hs__tap_1 TAP_1986 ();
 sky130_as_sc_hs__tap_1 TAP_1987 ();
 sky130_as_sc_hs__tap_1 TAP_1988 ();
 sky130_as_sc_hs__tap_1 TAP_1989 ();
 sky130_as_sc_hs__tap_1 TAP_1990 ();
 sky130_as_sc_hs__tap_1 TAP_1991 ();
 sky130_as_sc_hs__tap_1 TAP_1992 ();
 sky130_as_sc_hs__tap_1 TAP_1993 ();
 sky130_as_sc_hs__tap_1 TAP_1994 ();
 sky130_as_sc_hs__tap_1 TAP_1995 ();
 sky130_as_sc_hs__tap_1 TAP_1996 ();
 sky130_as_sc_hs__tap_1 TAP_1997 ();
 sky130_as_sc_hs__tap_1 TAP_1998 ();
 sky130_as_sc_hs__tap_1 TAP_1999 ();
 sky130_as_sc_hs__tap_1 TAP_2000 ();
 sky130_as_sc_hs__tap_1 TAP_2001 ();
 sky130_as_sc_hs__tap_1 TAP_2002 ();
 sky130_as_sc_hs__tap_1 TAP_2003 ();
 sky130_as_sc_hs__tap_1 TAP_2004 ();
 sky130_as_sc_hs__tap_1 TAP_2005 ();
 sky130_as_sc_hs__tap_1 TAP_2006 ();
 sky130_as_sc_hs__tap_1 TAP_2007 ();
 sky130_as_sc_hs__tap_1 TAP_2008 ();
 sky130_as_sc_hs__tap_1 TAP_2009 ();
 sky130_as_sc_hs__tap_1 TAP_2010 ();
 sky130_as_sc_hs__tap_1 TAP_2011 ();
 sky130_as_sc_hs__tap_1 TAP_2012 ();
 sky130_as_sc_hs__tap_1 TAP_2013 ();
 sky130_as_sc_hs__tap_1 TAP_2014 ();
 sky130_as_sc_hs__tap_1 TAP_2015 ();
 sky130_as_sc_hs__tap_1 TAP_2016 ();
 sky130_as_sc_hs__tap_1 TAP_2017 ();
 sky130_as_sc_hs__tap_1 TAP_2018 ();
 sky130_as_sc_hs__tap_1 TAP_2019 ();
 sky130_as_sc_hs__tap_1 TAP_2020 ();
 sky130_as_sc_hs__tap_1 TAP_2021 ();
 sky130_as_sc_hs__tap_1 TAP_2022 ();
 sky130_as_sc_hs__tap_1 TAP_2023 ();
 sky130_as_sc_hs__tap_1 TAP_2024 ();
 sky130_as_sc_hs__tap_1 TAP_2025 ();
 sky130_as_sc_hs__tap_1 TAP_2026 ();
 sky130_as_sc_hs__tap_1 TAP_2027 ();
 sky130_as_sc_hs__tap_1 TAP_2028 ();
 sky130_as_sc_hs__tap_1 TAP_2029 ();
 sky130_as_sc_hs__tap_1 TAP_2030 ();
 sky130_as_sc_hs__tap_1 TAP_2031 ();
 sky130_as_sc_hs__tap_1 TAP_2032 ();
 sky130_as_sc_hs__tap_1 TAP_2033 ();
 sky130_as_sc_hs__tap_1 TAP_2034 ();
 sky130_as_sc_hs__tap_1 TAP_2035 ();
 sky130_as_sc_hs__tap_1 TAP_2036 ();
 sky130_as_sc_hs__tap_1 TAP_2037 ();
 sky130_as_sc_hs__tap_1 TAP_2038 ();
 sky130_as_sc_hs__tap_1 TAP_2039 ();
 sky130_as_sc_hs__tap_1 TAP_2040 ();
 sky130_as_sc_hs__tap_1 TAP_2041 ();
 sky130_as_sc_hs__tap_1 TAP_2042 ();
 sky130_as_sc_hs__tap_1 TAP_2043 ();
 sky130_as_sc_hs__tap_1 TAP_2044 ();
 sky130_as_sc_hs__tap_1 TAP_2045 ();
 sky130_as_sc_hs__tap_1 TAP_2046 ();
 sky130_as_sc_hs__tap_1 TAP_2047 ();
 sky130_as_sc_hs__tap_1 TAP_2048 ();
 sky130_as_sc_hs__tap_1 TAP_2049 ();
 sky130_as_sc_hs__tap_1 TAP_2050 ();
 sky130_as_sc_hs__tap_1 TAP_2051 ();
 sky130_as_sc_hs__tap_1 TAP_2052 ();
 sky130_as_sc_hs__tap_1 TAP_2053 ();
 sky130_as_sc_hs__tap_1 TAP_2054 ();
 sky130_as_sc_hs__tap_1 TAP_2055 ();
 sky130_as_sc_hs__tap_1 TAP_2056 ();
 sky130_as_sc_hs__tap_1 TAP_2057 ();
 sky130_as_sc_hs__tap_1 TAP_2058 ();
 sky130_as_sc_hs__tap_1 TAP_2059 ();
 sky130_as_sc_hs__tap_1 TAP_2060 ();
 sky130_as_sc_hs__tap_1 TAP_2061 ();
 sky130_as_sc_hs__tap_1 TAP_2062 ();
 sky130_as_sc_hs__tap_1 TAP_2063 ();
 sky130_as_sc_hs__tap_1 TAP_2064 ();
 sky130_as_sc_hs__tap_1 TAP_2065 ();
 sky130_as_sc_hs__tap_1 TAP_2066 ();
 sky130_as_sc_hs__tap_1 TAP_2067 ();
 sky130_as_sc_hs__tap_1 TAP_2068 ();
 sky130_as_sc_hs__tap_1 TAP_2069 ();
 sky130_as_sc_hs__tap_1 TAP_2070 ();
 sky130_as_sc_hs__tap_1 TAP_2071 ();
 sky130_as_sc_hs__tap_1 TAP_2072 ();
 sky130_as_sc_hs__tap_1 TAP_2073 ();
 sky130_as_sc_hs__tap_1 TAP_2074 ();
 sky130_as_sc_hs__tap_1 TAP_2075 ();
 sky130_as_sc_hs__tap_1 TAP_2076 ();
 sky130_as_sc_hs__tap_1 TAP_2077 ();
 sky130_as_sc_hs__tap_1 TAP_2078 ();
 sky130_as_sc_hs__tap_1 TAP_2079 ();
 sky130_as_sc_hs__tap_1 TAP_2080 ();
 sky130_as_sc_hs__tap_1 TAP_2081 ();
 sky130_as_sc_hs__tap_1 TAP_2082 ();
 sky130_as_sc_hs__tap_1 TAP_2083 ();
 sky130_as_sc_hs__tap_1 TAP_2084 ();
 sky130_as_sc_hs__tap_1 TAP_2085 ();
 sky130_as_sc_hs__tap_1 TAP_2086 ();
 sky130_as_sc_hs__tap_1 TAP_2087 ();
 sky130_as_sc_hs__tap_1 TAP_2088 ();
 sky130_as_sc_hs__tap_1 TAP_2089 ();
 sky130_as_sc_hs__tap_1 TAP_2090 ();
 sky130_as_sc_hs__tap_1 TAP_2091 ();
 sky130_as_sc_hs__tap_1 TAP_2092 ();
 sky130_as_sc_hs__tap_1 TAP_2093 ();
 sky130_as_sc_hs__tap_1 TAP_2094 ();
 sky130_as_sc_hs__tap_1 TAP_2095 ();
 sky130_as_sc_hs__tap_1 TAP_2096 ();
 sky130_as_sc_hs__tap_1 TAP_2097 ();
 sky130_as_sc_hs__tap_1 TAP_2098 ();
 sky130_as_sc_hs__tap_1 TAP_2099 ();
 sky130_as_sc_hs__tap_1 TAP_2100 ();
 sky130_as_sc_hs__tap_1 TAP_2101 ();
 sky130_as_sc_hs__tap_1 TAP_2102 ();
 sky130_as_sc_hs__tap_1 TAP_2103 ();
 sky130_as_sc_hs__tap_1 TAP_2104 ();
 sky130_as_sc_hs__tap_1 TAP_2105 ();
 sky130_as_sc_hs__tap_1 TAP_2106 ();
 sky130_as_sc_hs__tap_1 TAP_2107 ();
 sky130_as_sc_hs__tap_1 TAP_2108 ();
 sky130_as_sc_hs__tap_1 TAP_2109 ();
 sky130_as_sc_hs__tap_1 TAP_2110 ();
 sky130_as_sc_hs__tap_1 TAP_2111 ();
 sky130_as_sc_hs__tap_1 TAP_2112 ();
 sky130_as_sc_hs__tap_1 TAP_2113 ();
 sky130_as_sc_hs__tap_1 TAP_2114 ();
 sky130_as_sc_hs__tap_1 TAP_2115 ();
 sky130_as_sc_hs__tap_1 TAP_2116 ();
 sky130_as_sc_hs__tap_1 TAP_2117 ();
 sky130_as_sc_hs__tap_1 TAP_2118 ();
 sky130_as_sc_hs__tap_1 TAP_2119 ();
 sky130_as_sc_hs__tap_1 TAP_2120 ();
 sky130_as_sc_hs__tap_1 TAP_2121 ();
 sky130_as_sc_hs__tap_1 TAP_2122 ();
 sky130_as_sc_hs__tap_1 TAP_2123 ();
 sky130_as_sc_hs__tap_1 TAP_2124 ();
 sky130_as_sc_hs__tap_1 TAP_2125 ();
 sky130_as_sc_hs__tap_1 TAP_2126 ();
 sky130_as_sc_hs__tap_1 TAP_2127 ();
 sky130_as_sc_hs__tap_1 TAP_2128 ();
 sky130_as_sc_hs__tap_1 TAP_2129 ();
 sky130_as_sc_hs__tap_1 TAP_2130 ();
 sky130_as_sc_hs__tap_1 TAP_2131 ();
 sky130_as_sc_hs__tap_1 TAP_2132 ();
 sky130_as_sc_hs__tap_1 TAP_2133 ();
 sky130_as_sc_hs__tap_1 TAP_2134 ();
 sky130_as_sc_hs__tap_1 TAP_2135 ();
 sky130_as_sc_hs__tap_1 TAP_2136 ();
 sky130_as_sc_hs__tap_1 TAP_2137 ();
 sky130_as_sc_hs__tap_1 TAP_2138 ();
 sky130_as_sc_hs__tap_1 TAP_2139 ();
 sky130_as_sc_hs__tap_1 TAP_2140 ();
 sky130_as_sc_hs__tap_1 TAP_2141 ();
 sky130_as_sc_hs__tap_1 TAP_2142 ();
 sky130_as_sc_hs__tap_1 TAP_2143 ();
 sky130_as_sc_hs__tap_1 TAP_2144 ();
 sky130_as_sc_hs__tap_1 TAP_2145 ();
 sky130_as_sc_hs__tap_1 TAP_2146 ();
 sky130_as_sc_hs__tap_1 TAP_2147 ();
 sky130_as_sc_hs__tap_1 TAP_2148 ();
 sky130_as_sc_hs__tap_1 TAP_2149 ();
 sky130_as_sc_hs__tap_1 TAP_2150 ();
 sky130_as_sc_hs__tap_1 TAP_2151 ();
 sky130_as_sc_hs__tap_1 TAP_2152 ();
 sky130_as_sc_hs__tap_1 TAP_2153 ();
 sky130_as_sc_hs__tap_1 TAP_2154 ();
 sky130_as_sc_hs__tap_1 TAP_2155 ();
 sky130_as_sc_hs__tap_1 TAP_2156 ();
 sky130_as_sc_hs__tap_1 TAP_2157 ();
 sky130_as_sc_hs__tap_1 TAP_2158 ();
 sky130_as_sc_hs__tap_1 TAP_2159 ();
 sky130_as_sc_hs__tap_1 TAP_2160 ();
 sky130_as_sc_hs__tap_1 TAP_2161 ();
 sky130_as_sc_hs__tap_1 TAP_2162 ();
 sky130_as_sc_hs__tap_1 TAP_2163 ();
 sky130_as_sc_hs__tap_1 TAP_2164 ();
 sky130_as_sc_hs__tap_1 TAP_2165 ();
 sky130_as_sc_hs__tap_1 TAP_2166 ();
 sky130_as_sc_hs__tap_1 TAP_2167 ();
 sky130_as_sc_hs__tap_1 TAP_2168 ();
 sky130_as_sc_hs__tap_1 TAP_2169 ();
 sky130_as_sc_hs__tap_1 TAP_2170 ();
 sky130_as_sc_hs__tap_1 TAP_2171 ();
 sky130_as_sc_hs__tap_1 TAP_2172 ();
 sky130_as_sc_hs__tap_1 TAP_2173 ();
 sky130_as_sc_hs__tap_1 TAP_2174 ();
 sky130_as_sc_hs__tap_1 TAP_2175 ();
 sky130_as_sc_hs__tap_1 TAP_2176 ();
 sky130_as_sc_hs__tap_1 TAP_2177 ();
 sky130_as_sc_hs__tap_1 TAP_2178 ();
 sky130_as_sc_hs__tap_1 TAP_2179 ();
 sky130_as_sc_hs__tap_1 TAP_2180 ();
 sky130_as_sc_hs__tap_1 TAP_2181 ();
 sky130_as_sc_hs__tap_1 TAP_2182 ();
 sky130_as_sc_hs__tap_1 TAP_2183 ();
 sky130_as_sc_hs__tap_1 TAP_2184 ();
 sky130_as_sc_hs__tap_1 TAP_2185 ();
 sky130_as_sc_hs__tap_1 TAP_2186 ();
 sky130_as_sc_hs__tap_1 TAP_2187 ();
 sky130_as_sc_hs__tap_1 TAP_2188 ();
 sky130_as_sc_hs__tap_1 TAP_2189 ();
 sky130_as_sc_hs__tap_1 TAP_2190 ();
 sky130_as_sc_hs__tap_1 TAP_2191 ();
 sky130_as_sc_hs__tap_1 TAP_2192 ();
 sky130_as_sc_hs__tap_1 TAP_2193 ();
 sky130_as_sc_hs__tap_1 TAP_2194 ();
 sky130_as_sc_hs__tap_1 TAP_2195 ();
 sky130_as_sc_hs__tap_1 TAP_2196 ();
 sky130_as_sc_hs__tap_1 TAP_2197 ();
 sky130_as_sc_hs__tap_1 TAP_2198 ();
 sky130_as_sc_hs__tap_1 TAP_2199 ();
 sky130_as_sc_hs__tap_1 TAP_2200 ();
 sky130_as_sc_hs__tap_1 TAP_2201 ();
 sky130_as_sc_hs__tap_1 TAP_2202 ();
 sky130_as_sc_hs__tap_1 TAP_2203 ();
 sky130_as_sc_hs__tap_1 TAP_2204 ();
 sky130_as_sc_hs__tap_1 TAP_2205 ();
 sky130_as_sc_hs__tap_1 TAP_2206 ();
 sky130_as_sc_hs__tap_1 TAP_2207 ();
 sky130_as_sc_hs__tap_1 TAP_2208 ();
 sky130_as_sc_hs__tap_1 TAP_2209 ();
 sky130_as_sc_hs__tap_1 TAP_2210 ();
 sky130_as_sc_hs__tap_1 TAP_2211 ();
 sky130_as_sc_hs__tap_1 TAP_2212 ();
 sky130_as_sc_hs__tap_1 TAP_2213 ();
 sky130_as_sc_hs__tap_1 TAP_2214 ();
 sky130_as_sc_hs__tap_1 TAP_2215 ();
 sky130_as_sc_hs__tap_1 TAP_2216 ();
 sky130_as_sc_hs__tap_1 TAP_2217 ();
 sky130_as_sc_hs__tap_1 TAP_2218 ();
 sky130_as_sc_hs__tap_1 TAP_2219 ();
 sky130_as_sc_hs__tap_1 TAP_2220 ();
 sky130_as_sc_hs__tap_1 TAP_2221 ();
 sky130_as_sc_hs__tap_1 TAP_2222 ();
 sky130_as_sc_hs__tap_1 TAP_2223 ();
 sky130_as_sc_hs__tap_1 TAP_2224 ();
 sky130_as_sc_hs__tap_1 TAP_2225 ();
 sky130_as_sc_hs__tap_1 TAP_2226 ();
 sky130_as_sc_hs__tap_1 TAP_2227 ();
 sky130_as_sc_hs__tap_1 TAP_2228 ();
 sky130_as_sc_hs__tap_1 TAP_2229 ();
 sky130_as_sc_hs__tap_1 TAP_2230 ();
 sky130_as_sc_hs__tap_1 TAP_2231 ();
 sky130_as_sc_hs__tap_1 TAP_2232 ();
 sky130_as_sc_hs__tap_1 TAP_2233 ();
 sky130_as_sc_hs__tap_1 TAP_2234 ();
 sky130_as_sc_hs__tap_1 TAP_2235 ();
 sky130_as_sc_hs__tap_1 TAP_2236 ();
 sky130_as_sc_hs__tap_1 TAP_2237 ();
 sky130_as_sc_hs__tap_1 TAP_2238 ();
 sky130_as_sc_hs__tap_1 TAP_2239 ();
 sky130_as_sc_hs__tap_1 TAP_2240 ();
 sky130_as_sc_hs__tap_1 TAP_2241 ();
 sky130_as_sc_hs__tap_1 TAP_2242 ();
 sky130_as_sc_hs__tap_1 TAP_2243 ();
 sky130_as_sc_hs__tap_1 TAP_2244 ();
 sky130_as_sc_hs__tap_1 TAP_2245 ();
 sky130_as_sc_hs__tap_1 TAP_2246 ();
 sky130_as_sc_hs__tap_1 TAP_2247 ();
 sky130_as_sc_hs__tap_1 TAP_2248 ();
 sky130_as_sc_hs__tap_1 TAP_2249 ();
 sky130_as_sc_hs__tap_1 TAP_2250 ();
 sky130_as_sc_hs__tap_1 TAP_2251 ();
 sky130_as_sc_hs__tap_1 TAP_2252 ();
 sky130_as_sc_hs__tap_1 TAP_2253 ();
 sky130_as_sc_hs__tap_1 TAP_2254 ();
 sky130_as_sc_hs__tap_1 TAP_2255 ();
 sky130_as_sc_hs__tap_1 TAP_2256 ();
 sky130_as_sc_hs__tap_1 TAP_2257 ();
 sky130_as_sc_hs__tap_1 TAP_2258 ();
 sky130_as_sc_hs__tap_1 TAP_2259 ();
 sky130_as_sc_hs__tap_1 TAP_2260 ();
 sky130_as_sc_hs__tap_1 TAP_2261 ();
 sky130_as_sc_hs__tap_1 TAP_2262 ();
 sky130_as_sc_hs__tap_1 TAP_2263 ();
 sky130_as_sc_hs__tap_1 TAP_2264 ();
 sky130_as_sc_hs__tap_1 TAP_2265 ();
 sky130_as_sc_hs__tap_1 TAP_2266 ();
 sky130_as_sc_hs__tap_1 TAP_2267 ();
 sky130_as_sc_hs__tap_1 TAP_2268 ();
 sky130_as_sc_hs__tap_1 TAP_2269 ();
 sky130_as_sc_hs__tap_1 TAP_2270 ();
 sky130_as_sc_hs__tap_1 TAP_2271 ();
 sky130_as_sc_hs__tap_1 TAP_2272 ();
 sky130_as_sc_hs__tap_1 TAP_2273 ();
 sky130_as_sc_hs__tap_1 TAP_2274 ();
 sky130_as_sc_hs__tap_1 TAP_2275 ();
 sky130_as_sc_hs__tap_1 TAP_2276 ();
 sky130_as_sc_hs__tap_1 TAP_2277 ();
 sky130_as_sc_hs__tap_1 TAP_2278 ();
 sky130_as_sc_hs__tap_1 TAP_2279 ();
 sky130_as_sc_hs__tap_1 TAP_2280 ();
 sky130_as_sc_hs__tap_1 TAP_2281 ();
 sky130_as_sc_hs__tap_1 TAP_2282 ();
 sky130_as_sc_hs__tap_1 TAP_2283 ();
 sky130_as_sc_hs__tap_1 TAP_2284 ();
 sky130_as_sc_hs__tap_1 TAP_2285 ();
 sky130_as_sc_hs__tap_1 TAP_2286 ();
 sky130_as_sc_hs__tap_1 TAP_2287 ();
 sky130_as_sc_hs__tap_1 TAP_2288 ();
 sky130_as_sc_hs__tap_1 TAP_2289 ();
 sky130_as_sc_hs__tap_1 TAP_2290 ();
 sky130_as_sc_hs__tap_1 TAP_2291 ();
 sky130_as_sc_hs__tap_1 TAP_2292 ();
 sky130_as_sc_hs__tap_1 TAP_2293 ();
 sky130_as_sc_hs__tap_1 TAP_2294 ();
 sky130_as_sc_hs__tap_1 TAP_2295 ();
 sky130_as_sc_hs__tap_1 TAP_2296 ();
 sky130_as_sc_hs__tap_1 TAP_2297 ();
 sky130_as_sc_hs__tap_1 TAP_2298 ();
 sky130_as_sc_hs__tap_1 TAP_2299 ();
 sky130_as_sc_hs__tap_1 TAP_2300 ();
 sky130_as_sc_hs__tap_1 TAP_2301 ();
 sky130_as_sc_hs__tap_1 TAP_2302 ();
 sky130_as_sc_hs__tap_1 TAP_2303 ();
 sky130_as_sc_hs__tap_1 TAP_2304 ();
 sky130_as_sc_hs__tap_1 TAP_2305 ();
 sky130_as_sc_hs__tap_1 TAP_2306 ();
 sky130_as_sc_hs__tap_1 TAP_2307 ();
 sky130_as_sc_hs__tap_1 TAP_2308 ();
 sky130_as_sc_hs__tap_1 TAP_2309 ();
 sky130_as_sc_hs__tap_1 TAP_2310 ();
 sky130_as_sc_hs__tap_1 TAP_2311 ();
 sky130_as_sc_hs__tap_1 TAP_2312 ();
 sky130_as_sc_hs__tap_1 TAP_2313 ();
 sky130_as_sc_hs__tap_1 TAP_2314 ();
 sky130_as_sc_hs__tap_1 TAP_2315 ();
 sky130_as_sc_hs__tap_1 TAP_2316 ();
 sky130_as_sc_hs__tap_1 TAP_2317 ();
 sky130_as_sc_hs__tap_1 TAP_2318 ();
 sky130_as_sc_hs__tap_1 TAP_2319 ();
 sky130_as_sc_hs__tap_1 TAP_2320 ();
 sky130_as_sc_hs__tap_1 TAP_2321 ();
 sky130_as_sc_hs__tap_1 TAP_2322 ();
 sky130_as_sc_hs__tap_1 TAP_2323 ();
 sky130_as_sc_hs__tap_1 TAP_2324 ();
 sky130_as_sc_hs__tap_1 TAP_2325 ();
 sky130_as_sc_hs__tap_1 TAP_2326 ();
 sky130_as_sc_hs__tap_1 TAP_2327 ();
 sky130_as_sc_hs__tap_1 TAP_2328 ();
 sky130_as_sc_hs__tap_1 TAP_2329 ();
 sky130_as_sc_hs__tap_1 TAP_2330 ();
 sky130_as_sc_hs__tap_1 TAP_2331 ();
 sky130_as_sc_hs__tap_1 TAP_2332 ();
 sky130_as_sc_hs__tap_1 TAP_2333 ();
 sky130_as_sc_hs__tap_1 TAP_2334 ();
 sky130_as_sc_hs__tap_1 TAP_2335 ();
 sky130_as_sc_hs__tap_1 TAP_2336 ();
 sky130_as_sc_hs__tap_1 TAP_2337 ();
 sky130_as_sc_hs__tap_1 TAP_2338 ();
 sky130_as_sc_hs__tap_1 TAP_2339 ();
 sky130_as_sc_hs__tap_1 TAP_2340 ();
 sky130_as_sc_hs__tap_1 TAP_2341 ();
 sky130_as_sc_hs__tap_1 TAP_2342 ();
 sky130_as_sc_hs__tap_1 TAP_2343 ();
 sky130_as_sc_hs__tap_1 TAP_2344 ();
 sky130_as_sc_hs__tap_1 TAP_2345 ();
 sky130_as_sc_hs__tap_1 TAP_2346 ();
 sky130_as_sc_hs__tap_1 TAP_2347 ();
 sky130_as_sc_hs__tap_1 TAP_2348 ();
 sky130_as_sc_hs__tap_1 TAP_2349 ();
 sky130_as_sc_hs__tap_1 TAP_2350 ();
 sky130_as_sc_hs__tap_1 TAP_2351 ();
 sky130_as_sc_hs__tap_1 TAP_2352 ();
 sky130_as_sc_hs__tap_1 TAP_2353 ();
 sky130_as_sc_hs__tap_1 TAP_2354 ();
 sky130_as_sc_hs__tap_1 TAP_2355 ();
 sky130_as_sc_hs__tap_1 TAP_2356 ();
 sky130_as_sc_hs__tap_1 TAP_2357 ();
 sky130_as_sc_hs__tap_1 TAP_2358 ();
 sky130_as_sc_hs__tap_1 TAP_2359 ();
 sky130_as_sc_hs__tap_1 TAP_2360 ();
 sky130_as_sc_hs__tap_1 TAP_2361 ();
 sky130_as_sc_hs__tap_1 TAP_2362 ();
 sky130_as_sc_hs__tap_1 TAP_2363 ();
 sky130_as_sc_hs__tap_1 TAP_2364 ();
 sky130_as_sc_hs__tap_1 TAP_2365 ();
 sky130_as_sc_hs__tap_1 TAP_2366 ();
 sky130_as_sc_hs__tap_1 TAP_2367 ();
 sky130_as_sc_hs__tap_1 TAP_2368 ();
 sky130_as_sc_hs__tap_1 TAP_2369 ();
 sky130_as_sc_hs__tap_1 TAP_2370 ();
 sky130_as_sc_hs__tap_1 TAP_2371 ();
 sky130_as_sc_hs__tap_1 TAP_2372 ();
 sky130_as_sc_hs__tap_1 TAP_2373 ();
 sky130_as_sc_hs__tap_1 TAP_2374 ();
 sky130_as_sc_hs__tap_1 TAP_2375 ();
 sky130_as_sc_hs__tap_1 TAP_2376 ();
 sky130_as_sc_hs__tap_1 TAP_2377 ();
 sky130_as_sc_hs__tap_1 TAP_2378 ();
 sky130_as_sc_hs__tap_1 TAP_2379 ();
 sky130_as_sc_hs__tap_1 TAP_2380 ();
 sky130_as_sc_hs__tap_1 TAP_2381 ();
 sky130_as_sc_hs__tap_1 TAP_2382 ();
 sky130_as_sc_hs__tap_1 TAP_2383 ();
 sky130_as_sc_hs__tap_1 TAP_2384 ();
 sky130_as_sc_hs__tap_1 TAP_2385 ();
 sky130_as_sc_hs__tap_1 TAP_2386 ();
 sky130_as_sc_hs__tap_1 TAP_2387 ();
 sky130_as_sc_hs__tap_1 TAP_2388 ();
 sky130_as_sc_hs__tap_1 TAP_2389 ();
 sky130_as_sc_hs__tap_1 TAP_2390 ();
 sky130_as_sc_hs__tap_1 TAP_2391 ();
 sky130_as_sc_hs__tap_1 TAP_2392 ();
 sky130_as_sc_hs__tap_1 TAP_2393 ();
 sky130_as_sc_hs__tap_1 TAP_2394 ();
 sky130_as_sc_hs__tap_1 TAP_2395 ();
 sky130_as_sc_hs__tap_1 TAP_2396 ();
 sky130_as_sc_hs__tap_1 TAP_2397 ();
 sky130_as_sc_hs__tap_1 TAP_2398 ();
 sky130_as_sc_hs__tap_1 TAP_2399 ();
 sky130_as_sc_hs__tap_1 TAP_2400 ();
 sky130_as_sc_hs__tap_1 TAP_2401 ();
 sky130_as_sc_hs__tap_1 TAP_2402 ();
 sky130_as_sc_hs__tap_1 TAP_2403 ();
 sky130_as_sc_hs__tap_1 TAP_2404 ();
 sky130_as_sc_hs__tap_1 TAP_2405 ();
 sky130_as_sc_hs__tap_1 TAP_2406 ();
 sky130_as_sc_hs__tap_1 TAP_2407 ();
 sky130_as_sc_hs__tap_1 TAP_2408 ();
 sky130_as_sc_hs__tap_1 TAP_2409 ();
 sky130_as_sc_hs__tap_1 TAP_2410 ();
 sky130_as_sc_hs__tap_1 TAP_2411 ();
 sky130_as_sc_hs__tap_1 TAP_2412 ();
 sky130_as_sc_hs__tap_1 TAP_2413 ();
 sky130_as_sc_hs__tap_1 TAP_2414 ();
 sky130_as_sc_hs__tap_1 TAP_2415 ();
 sky130_as_sc_hs__tap_1 TAP_2416 ();
 sky130_as_sc_hs__tap_1 TAP_2417 ();
 sky130_as_sc_hs__tap_1 TAP_2418 ();
 sky130_as_sc_hs__tap_1 TAP_2419 ();
 sky130_as_sc_hs__tap_1 TAP_2420 ();
 sky130_as_sc_hs__tap_1 TAP_2421 ();
 sky130_as_sc_hs__tap_1 TAP_2422 ();
 sky130_as_sc_hs__tap_1 TAP_2423 ();
 sky130_as_sc_hs__tap_1 TAP_2424 ();
 sky130_as_sc_hs__tap_1 TAP_2425 ();
 sky130_as_sc_hs__tap_1 TAP_2426 ();
 sky130_as_sc_hs__tap_1 TAP_2427 ();
 sky130_as_sc_hs__tap_1 TAP_2428 ();
 sky130_as_sc_hs__tap_1 TAP_2429 ();
 sky130_as_sc_hs__tap_1 TAP_2430 ();
 sky130_as_sc_hs__tap_1 TAP_2431 ();
 sky130_as_sc_hs__tap_1 TAP_2432 ();
 sky130_as_sc_hs__tap_1 TAP_2433 ();
 sky130_as_sc_hs__tap_1 TAP_2434 ();
 sky130_as_sc_hs__tap_1 TAP_2435 ();
 sky130_as_sc_hs__tap_1 TAP_2436 ();
 sky130_as_sc_hs__tap_1 TAP_2437 ();
 sky130_as_sc_hs__tap_1 TAP_2438 ();
 sky130_as_sc_hs__tap_1 TAP_2439 ();
 sky130_as_sc_hs__tap_1 TAP_2440 ();
 sky130_as_sc_hs__tap_1 TAP_2441 ();
 sky130_as_sc_hs__tap_1 TAP_2442 ();
 sky130_as_sc_hs__tap_1 TAP_2443 ();
 sky130_as_sc_hs__tap_1 TAP_2444 ();
 sky130_as_sc_hs__tap_1 TAP_2445 ();
 sky130_as_sc_hs__tap_1 TAP_2446 ();
 sky130_as_sc_hs__tap_1 TAP_2447 ();
 sky130_as_sc_hs__tap_1 TAP_2448 ();
 sky130_as_sc_hs__tap_1 TAP_2449 ();
 sky130_as_sc_hs__tap_1 TAP_2450 ();
 sky130_as_sc_hs__tap_1 TAP_2451 ();
 sky130_as_sc_hs__tap_1 TAP_2452 ();
 sky130_as_sc_hs__tap_1 TAP_2453 ();
 sky130_as_sc_hs__tap_1 TAP_2454 ();
 sky130_as_sc_hs__tap_1 TAP_2455 ();
 sky130_as_sc_hs__tap_1 TAP_2456 ();
 sky130_as_sc_hs__tap_1 TAP_2457 ();
 sky130_as_sc_hs__tap_1 TAP_2458 ();
 sky130_as_sc_hs__tap_1 TAP_2459 ();
 sky130_as_sc_hs__tap_1 TAP_2460 ();
 sky130_as_sc_hs__tap_1 TAP_2461 ();
 sky130_as_sc_hs__tap_1 TAP_2462 ();
 sky130_as_sc_hs__tap_1 TAP_2463 ();
 sky130_as_sc_hs__tap_1 TAP_2464 ();
 sky130_as_sc_hs__tap_1 TAP_2465 ();
 sky130_as_sc_hs__tap_1 TAP_2466 ();
 sky130_as_sc_hs__tap_1 TAP_2467 ();
 sky130_as_sc_hs__tap_1 TAP_2468 ();
 sky130_as_sc_hs__tap_1 TAP_2469 ();
 sky130_as_sc_hs__tap_1 TAP_2470 ();
 sky130_as_sc_hs__tap_1 TAP_2471 ();
 sky130_as_sc_hs__tap_1 TAP_2472 ();
 sky130_as_sc_hs__tap_1 TAP_2473 ();
 sky130_as_sc_hs__tap_1 TAP_2474 ();
 sky130_as_sc_hs__tap_1 TAP_2475 ();
 sky130_as_sc_hs__tap_1 TAP_2476 ();
 sky130_as_sc_hs__tap_1 TAP_2477 ();
 sky130_as_sc_hs__tap_1 TAP_2478 ();
 sky130_as_sc_hs__tap_1 TAP_2479 ();
 sky130_as_sc_hs__tap_1 TAP_2480 ();
 sky130_as_sc_hs__tap_1 TAP_2481 ();
 sky130_as_sc_hs__tap_1 TAP_2482 ();
 sky130_as_sc_hs__tap_1 TAP_2483 ();
 sky130_as_sc_hs__tap_1 TAP_2484 ();
 sky130_as_sc_hs__tap_1 TAP_2485 ();
 sky130_as_sc_hs__tap_1 TAP_2486 ();
 sky130_as_sc_hs__tap_1 TAP_2487 ();
 sky130_as_sc_hs__tap_1 TAP_2488 ();
 sky130_as_sc_hs__tap_1 TAP_2489 ();
 sky130_as_sc_hs__tap_1 TAP_2490 ();
 sky130_as_sc_hs__tap_1 TAP_2491 ();
 sky130_as_sc_hs__tap_1 TAP_2492 ();
 sky130_as_sc_hs__tap_1 TAP_2493 ();
 sky130_as_sc_hs__tap_1 TAP_2494 ();
 sky130_as_sc_hs__tap_1 TAP_2495 ();
 sky130_as_sc_hs__tap_1 TAP_2496 ();
 sky130_as_sc_hs__tap_1 TAP_2497 ();
 sky130_as_sc_hs__tap_1 TAP_2498 ();
 sky130_as_sc_hs__tap_1 TAP_2499 ();
 sky130_as_sc_hs__tap_1 TAP_2500 ();
 sky130_as_sc_hs__tap_1 TAP_2501 ();
 sky130_as_sc_hs__tap_1 TAP_2502 ();
 sky130_as_sc_hs__tap_1 TAP_2503 ();
 sky130_as_sc_hs__tap_1 TAP_2504 ();
 sky130_as_sc_hs__tap_1 TAP_2505 ();
 sky130_as_sc_hs__tap_1 TAP_2506 ();
 sky130_as_sc_hs__tap_1 TAP_2507 ();
 sky130_as_sc_hs__tap_1 TAP_2508 ();
 sky130_as_sc_hs__tap_1 TAP_2509 ();
 sky130_as_sc_hs__tap_1 TAP_2510 ();
 sky130_as_sc_hs__tap_1 TAP_2511 ();
 sky130_as_sc_hs__tap_1 TAP_2512 ();
 sky130_as_sc_hs__tap_1 TAP_2513 ();
 sky130_as_sc_hs__tap_1 TAP_2514 ();
 sky130_as_sc_hs__tap_1 TAP_2515 ();
 sky130_as_sc_hs__tap_1 TAP_2516 ();
 sky130_as_sc_hs__tap_1 TAP_2517 ();
 sky130_as_sc_hs__tap_1 TAP_2518 ();
 sky130_as_sc_hs__tap_1 TAP_2519 ();
 sky130_as_sc_hs__tap_1 TAP_2520 ();
 sky130_as_sc_hs__tap_1 TAP_2521 ();
 sky130_as_sc_hs__tap_1 TAP_2522 ();
 sky130_as_sc_hs__tap_1 TAP_2523 ();
 sky130_as_sc_hs__tap_1 TAP_2524 ();
 sky130_as_sc_hs__tap_1 TAP_2525 ();
 sky130_as_sc_hs__tap_1 TAP_2526 ();
 sky130_as_sc_hs__tap_1 TAP_2527 ();
 sky130_as_sc_hs__tap_1 TAP_2528 ();
 sky130_as_sc_hs__tap_1 TAP_2529 ();
 sky130_as_sc_hs__tap_1 TAP_2530 ();
 sky130_as_sc_hs__tap_1 TAP_2531 ();
 sky130_as_sc_hs__tap_1 TAP_2532 ();
 sky130_as_sc_hs__tap_1 TAP_2533 ();
 sky130_as_sc_hs__tap_1 TAP_2534 ();
 sky130_as_sc_hs__tap_1 TAP_2535 ();
 sky130_as_sc_hs__tap_1 TAP_2536 ();
 sky130_as_sc_hs__tap_1 TAP_2537 ();
 sky130_as_sc_hs__tap_1 TAP_2538 ();
 sky130_as_sc_hs__tap_1 TAP_2539 ();
 sky130_as_sc_hs__tap_1 TAP_2540 ();
 sky130_as_sc_hs__tap_1 TAP_2541 ();
 sky130_as_sc_hs__tap_1 TAP_2542 ();
 sky130_as_sc_hs__tap_1 TAP_2543 ();
 sky130_as_sc_hs__tap_1 TAP_2544 ();
 sky130_as_sc_hs__tap_1 TAP_2545 ();
 sky130_as_sc_hs__tap_1 TAP_2546 ();
 sky130_as_sc_hs__tap_1 TAP_2547 ();
 sky130_as_sc_hs__tap_1 TAP_2548 ();
 sky130_as_sc_hs__tap_1 TAP_2549 ();
 sky130_as_sc_hs__tap_1 TAP_2550 ();
 sky130_as_sc_hs__tap_1 TAP_2551 ();
 sky130_as_sc_hs__tap_1 TAP_2552 ();
 sky130_as_sc_hs__tap_1 TAP_2553 ();
 sky130_as_sc_hs__tap_1 TAP_2554 ();
 sky130_as_sc_hs__tap_1 TAP_2555 ();
 sky130_as_sc_hs__tap_1 TAP_2556 ();
 sky130_as_sc_hs__tap_1 TAP_2557 ();
 sky130_as_sc_hs__tap_1 TAP_2558 ();
 sky130_as_sc_hs__tap_1 TAP_2559 ();
 sky130_as_sc_hs__tap_1 TAP_2560 ();
 sky130_as_sc_hs__tap_1 TAP_2561 ();
 sky130_as_sc_hs__tap_1 TAP_2562 ();
 sky130_as_sc_hs__tap_1 TAP_2563 ();
 sky130_as_sc_hs__tap_1 TAP_2564 ();
 sky130_as_sc_hs__tap_1 TAP_2565 ();
 sky130_as_sc_hs__tap_1 TAP_2566 ();
 sky130_as_sc_hs__tap_1 TAP_2567 ();
 sky130_as_sc_hs__tap_1 TAP_2568 ();
 sky130_as_sc_hs__tap_1 TAP_2569 ();
 sky130_as_sc_hs__tap_1 TAP_2570 ();
 sky130_as_sc_hs__tap_1 TAP_2571 ();
 sky130_as_sc_hs__tap_1 TAP_2572 ();
 sky130_as_sc_hs__tap_1 TAP_2573 ();
 sky130_as_sc_hs__tap_1 TAP_2574 ();
 sky130_as_sc_hs__tap_1 TAP_2575 ();
 sky130_as_sc_hs__tap_1 TAP_2576 ();
 sky130_as_sc_hs__tap_1 TAP_2577 ();
 sky130_as_sc_hs__tap_1 TAP_2578 ();
 sky130_as_sc_hs__tap_1 TAP_2579 ();
 sky130_as_sc_hs__tap_1 TAP_2580 ();
 sky130_as_sc_hs__tap_1 TAP_2581 ();
 sky130_as_sc_hs__tap_1 TAP_2582 ();
 sky130_as_sc_hs__tap_1 TAP_2583 ();
 sky130_as_sc_hs__tap_1 TAP_2584 ();
 sky130_as_sc_hs__tap_1 TAP_2585 ();
 sky130_as_sc_hs__tap_1 TAP_2586 ();
 sky130_as_sc_hs__tap_1 TAP_2587 ();
 sky130_as_sc_hs__tap_1 TAP_2588 ();
 sky130_as_sc_hs__tap_1 TAP_2589 ();
 sky130_as_sc_hs__tap_1 TAP_2590 ();
 sky130_as_sc_hs__tap_1 TAP_2591 ();
 sky130_as_sc_hs__tap_1 TAP_2592 ();
 sky130_as_sc_hs__tap_1 TAP_2593 ();
 sky130_as_sc_hs__tap_1 TAP_2594 ();
 sky130_as_sc_hs__tap_1 TAP_2595 ();
 sky130_as_sc_hs__tap_1 TAP_2596 ();
 sky130_as_sc_hs__tap_1 TAP_2597 ();
 sky130_as_sc_hs__tap_1 TAP_2598 ();
 sky130_as_sc_hs__tap_1 TAP_2599 ();
 sky130_as_sc_hs__tap_1 TAP_2600 ();
 sky130_as_sc_hs__tap_1 TAP_2601 ();
 sky130_as_sc_hs__tap_1 TAP_2602 ();
 sky130_as_sc_hs__tap_1 TAP_2603 ();
 sky130_as_sc_hs__tap_1 TAP_2604 ();
 sky130_as_sc_hs__tap_1 TAP_2605 ();
 sky130_as_sc_hs__tap_1 TAP_2606 ();
 sky130_as_sc_hs__tap_1 TAP_2607 ();
 sky130_as_sc_hs__tap_1 TAP_2608 ();
 sky130_as_sc_hs__tap_1 TAP_2609 ();
 sky130_as_sc_hs__tap_1 TAP_2610 ();
 sky130_as_sc_hs__tap_1 TAP_2611 ();
 sky130_as_sc_hs__tap_1 TAP_2612 ();
 sky130_as_sc_hs__tap_1 TAP_2613 ();
 sky130_as_sc_hs__tap_1 TAP_2614 ();
 sky130_as_sc_hs__tap_1 TAP_2615 ();
 sky130_as_sc_hs__tap_1 TAP_2616 ();
 sky130_as_sc_hs__tap_1 TAP_2617 ();
 sky130_as_sc_hs__tap_1 TAP_2618 ();
 sky130_as_sc_hs__tap_1 TAP_2619 ();
 sky130_as_sc_hs__tap_1 TAP_2620 ();
 sky130_as_sc_hs__tap_1 TAP_2621 ();
 sky130_as_sc_hs__tap_1 TAP_2622 ();
 sky130_as_sc_hs__tap_1 TAP_2623 ();
 sky130_as_sc_hs__tap_1 TAP_2624 ();
 sky130_as_sc_hs__tap_1 TAP_2625 ();
 sky130_as_sc_hs__tap_1 TAP_2626 ();
 sky130_as_sc_hs__tap_1 TAP_2627 ();
 sky130_as_sc_hs__tap_1 TAP_2628 ();
 sky130_as_sc_hs__tap_1 TAP_2629 ();
 sky130_as_sc_hs__tap_1 TAP_2630 ();
 sky130_as_sc_hs__tap_1 TAP_2631 ();
 sky130_as_sc_hs__tap_1 TAP_2632 ();
 sky130_as_sc_hs__tap_1 TAP_2633 ();
 sky130_as_sc_hs__tap_1 TAP_2634 ();
 sky130_as_sc_hs__tap_1 TAP_2635 ();
 sky130_as_sc_hs__tap_1 TAP_2636 ();
 sky130_as_sc_hs__tap_1 TAP_2637 ();
 sky130_as_sc_hs__tap_1 TAP_2638 ();
 sky130_as_sc_hs__tap_1 TAP_2639 ();
 sky130_as_sc_hs__tap_1 TAP_2640 ();
 sky130_as_sc_hs__tap_1 TAP_2641 ();
 sky130_as_sc_hs__tap_1 TAP_2642 ();
 sky130_as_sc_hs__tap_1 TAP_2643 ();
 sky130_as_sc_hs__tap_1 TAP_2644 ();
 sky130_as_sc_hs__tap_1 TAP_2645 ();
 sky130_as_sc_hs__tap_1 TAP_2646 ();
 sky130_as_sc_hs__tap_1 TAP_2647 ();
 sky130_as_sc_hs__tap_1 TAP_2648 ();
 sky130_as_sc_hs__tap_1 TAP_2649 ();
 sky130_as_sc_hs__tap_1 TAP_2650 ();
 sky130_as_sc_hs__tap_1 TAP_2651 ();
 sky130_as_sc_hs__tap_1 TAP_2652 ();
 sky130_as_sc_hs__tap_1 TAP_2653 ();
 sky130_as_sc_hs__tap_1 TAP_2654 ();
 sky130_as_sc_hs__tap_1 TAP_2655 ();
 sky130_as_sc_hs__tap_1 TAP_2656 ();
 sky130_as_sc_hs__tap_1 TAP_2657 ();
 sky130_as_sc_hs__tap_1 TAP_2658 ();
 sky130_as_sc_hs__tap_1 TAP_2659 ();
 sky130_as_sc_hs__tap_1 TAP_2660 ();
 sky130_as_sc_hs__tap_1 TAP_2661 ();
 sky130_as_sc_hs__tap_1 TAP_2662 ();
 sky130_as_sc_hs__tap_1 TAP_2663 ();
 sky130_as_sc_hs__tap_1 TAP_2664 ();
 sky130_as_sc_hs__tap_1 TAP_2665 ();
 sky130_as_sc_hs__tap_1 TAP_2666 ();
 sky130_as_sc_hs__tap_1 TAP_2667 ();
 sky130_as_sc_hs__tap_1 TAP_2668 ();
 sky130_as_sc_hs__tap_1 TAP_2669 ();
 sky130_as_sc_hs__tap_1 TAP_2670 ();
 sky130_as_sc_hs__tap_1 TAP_2671 ();
 sky130_as_sc_hs__tap_1 TAP_2672 ();
 sky130_as_sc_hs__tap_1 TAP_2673 ();
 sky130_as_sc_hs__tap_1 TAP_2674 ();
 sky130_as_sc_hs__tap_1 TAP_2675 ();
 sky130_as_sc_hs__tap_1 TAP_2676 ();
 sky130_as_sc_hs__tap_1 TAP_2677 ();
 sky130_as_sc_hs__tap_1 TAP_2678 ();
 sky130_as_sc_hs__tap_1 TAP_2679 ();
 sky130_as_sc_hs__tap_1 TAP_2680 ();
 sky130_as_sc_hs__tap_1 TAP_2681 ();
 sky130_as_sc_hs__tap_1 TAP_2682 ();
 sky130_as_sc_hs__tap_1 TAP_2683 ();
 sky130_as_sc_hs__tap_1 TAP_2684 ();
 sky130_as_sc_hs__tap_1 TAP_2685 ();
 sky130_as_sc_hs__tap_1 TAP_2686 ();
 sky130_as_sc_hs__tap_1 TAP_2687 ();
 sky130_as_sc_hs__tap_1 TAP_2688 ();
 sky130_as_sc_hs__tap_1 TAP_2689 ();
 sky130_as_sc_hs__tap_1 TAP_2690 ();
 sky130_as_sc_hs__tap_1 TAP_2691 ();
 sky130_as_sc_hs__tap_1 TAP_2692 ();
 sky130_as_sc_hs__tap_1 TAP_2693 ();
 sky130_as_sc_hs__tap_1 TAP_2694 ();
 sky130_as_sc_hs__tap_1 TAP_2695 ();
 sky130_as_sc_hs__tap_1 TAP_2696 ();
 sky130_as_sc_hs__tap_1 TAP_2697 ();
 sky130_as_sc_hs__tap_1 TAP_2698 ();
 sky130_as_sc_hs__tap_1 TAP_2699 ();
 sky130_as_sc_hs__tap_1 TAP_2700 ();
 sky130_as_sc_hs__tap_1 TAP_2701 ();
 sky130_as_sc_hs__tap_1 TAP_2702 ();
 sky130_as_sc_hs__tap_1 TAP_2703 ();
 sky130_as_sc_hs__tap_1 TAP_2704 ();
 sky130_as_sc_hs__tap_1 TAP_2705 ();
 sky130_as_sc_hs__tap_1 TAP_2706 ();
 sky130_as_sc_hs__tap_1 TAP_2707 ();
 sky130_as_sc_hs__tap_1 TAP_2708 ();
 sky130_as_sc_hs__tap_1 TAP_2709 ();
 sky130_as_sc_hs__tap_1 TAP_2710 ();
 sky130_as_sc_hs__tap_1 TAP_2711 ();
 sky130_as_sc_hs__tap_1 TAP_2712 ();
 sky130_as_sc_hs__tap_1 TAP_2713 ();
 sky130_as_sc_hs__tap_1 TAP_2714 ();
 sky130_as_sc_hs__tap_1 TAP_2715 ();
 sky130_as_sc_hs__tap_1 TAP_2716 ();
 sky130_as_sc_hs__tap_1 TAP_2717 ();
 sky130_as_sc_hs__tap_1 TAP_2718 ();
 sky130_as_sc_hs__tap_1 TAP_2719 ();
 sky130_as_sc_hs__tap_1 TAP_2720 ();
 sky130_as_sc_hs__tap_1 TAP_2721 ();
 sky130_as_sc_hs__tap_1 TAP_2722 ();
 sky130_as_sc_hs__tap_1 TAP_2723 ();
 sky130_as_sc_hs__tap_1 TAP_2724 ();
 sky130_as_sc_hs__tap_1 TAP_2725 ();
 sky130_as_sc_hs__tap_1 TAP_2726 ();
 sky130_as_sc_hs__tap_1 TAP_2727 ();
 sky130_as_sc_hs__tap_1 TAP_2728 ();
 sky130_as_sc_hs__tap_1 TAP_2729 ();
 sky130_as_sc_hs__tap_1 TAP_2730 ();
 sky130_as_sc_hs__tap_1 TAP_2731 ();
 sky130_as_sc_hs__tap_1 TAP_2732 ();
 sky130_as_sc_hs__tap_1 TAP_2733 ();
 sky130_as_sc_hs__tap_1 TAP_2734 ();
 sky130_as_sc_hs__tap_1 TAP_2735 ();
 sky130_as_sc_hs__tap_1 TAP_2736 ();
 sky130_as_sc_hs__tap_1 TAP_2737 ();
 sky130_as_sc_hs__tap_1 TAP_2738 ();
 sky130_as_sc_hs__tap_1 TAP_2739 ();
 sky130_as_sc_hs__tap_1 TAP_2740 ();
 sky130_as_sc_hs__tap_1 TAP_2741 ();
 sky130_as_sc_hs__tap_1 TAP_2742 ();
 sky130_as_sc_hs__tap_1 TAP_2743 ();
 sky130_as_sc_hs__tap_1 TAP_2744 ();
 sky130_as_sc_hs__tap_1 TAP_2745 ();
 sky130_as_sc_hs__tap_1 TAP_2746 ();
 sky130_as_sc_hs__tap_1 TAP_2747 ();
 sky130_as_sc_hs__tap_1 TAP_2748 ();
 sky130_as_sc_hs__tap_1 TAP_2749 ();
 sky130_as_sc_hs__tap_1 TAP_2750 ();
 sky130_as_sc_hs__tap_1 TAP_2751 ();
 sky130_as_sc_hs__tap_1 TAP_2752 ();
 sky130_as_sc_hs__tap_1 TAP_2753 ();
 sky130_as_sc_hs__tap_1 TAP_2754 ();
 sky130_as_sc_hs__tap_1 TAP_2755 ();
 sky130_as_sc_hs__tap_1 TAP_2756 ();
 sky130_as_sc_hs__tap_1 TAP_2757 ();
 sky130_as_sc_hs__tap_1 TAP_2758 ();
 sky130_as_sc_hs__tap_1 TAP_2759 ();
 sky130_as_sc_hs__tap_1 TAP_2760 ();
 sky130_as_sc_hs__tap_1 TAP_2761 ();
 sky130_as_sc_hs__tap_1 TAP_2762 ();
 sky130_as_sc_hs__tap_1 TAP_2763 ();
 sky130_as_sc_hs__tap_1 TAP_2764 ();
 sky130_as_sc_hs__tap_1 TAP_2765 ();
 sky130_as_sc_hs__tap_1 TAP_2766 ();
 sky130_as_sc_hs__tap_1 TAP_2767 ();
 sky130_as_sc_hs__tap_1 TAP_2768 ();
 sky130_as_sc_hs__tap_1 TAP_2769 ();
 sky130_as_sc_hs__tap_1 TAP_2770 ();
 sky130_as_sc_hs__tap_1 TAP_2771 ();
 sky130_as_sc_hs__tap_1 TAP_2772 ();
 sky130_as_sc_hs__tap_1 TAP_2773 ();
 sky130_as_sc_hs__tap_1 TAP_2774 ();
 sky130_as_sc_hs__tap_1 TAP_2775 ();
 sky130_as_sc_hs__tap_1 TAP_2776 ();
 sky130_as_sc_hs__tap_1 TAP_2777 ();
 sky130_as_sc_hs__tap_1 TAP_2778 ();
 sky130_as_sc_hs__tap_1 TAP_2779 ();
 sky130_as_sc_hs__tap_1 TAP_2780 ();
 sky130_as_sc_hs__tap_1 TAP_2781 ();
 sky130_as_sc_hs__tap_1 TAP_2782 ();
 sky130_as_sc_hs__tap_1 TAP_2783 ();
 sky130_as_sc_hs__tap_1 TAP_2784 ();
 sky130_as_sc_hs__tap_1 TAP_2785 ();
 sky130_as_sc_hs__tap_1 TAP_2786 ();
 sky130_as_sc_hs__tap_1 TAP_2787 ();
 sky130_as_sc_hs__tap_1 TAP_2788 ();
 sky130_as_sc_hs__tap_1 TAP_2789 ();
 sky130_as_sc_hs__tap_1 TAP_2790 ();
 sky130_as_sc_hs__tap_1 TAP_2791 ();
 sky130_as_sc_hs__tap_1 TAP_2792 ();
 sky130_as_sc_hs__tap_1 TAP_2793 ();
 sky130_as_sc_hs__tap_1 TAP_2794 ();
 sky130_as_sc_hs__tap_1 TAP_2795 ();
 sky130_as_sc_hs__tap_1 TAP_2796 ();
 sky130_as_sc_hs__tap_1 TAP_2797 ();
 sky130_as_sc_hs__tap_1 TAP_2798 ();
 sky130_as_sc_hs__tap_1 TAP_2799 ();
 sky130_as_sc_hs__tap_1 TAP_2800 ();
 sky130_as_sc_hs__tap_1 TAP_2801 ();
 sky130_as_sc_hs__tap_1 TAP_2802 ();
 sky130_as_sc_hs__tap_1 TAP_2803 ();
 sky130_as_sc_hs__tap_1 TAP_2804 ();
 sky130_as_sc_hs__tap_1 TAP_2805 ();
 sky130_as_sc_hs__tap_1 TAP_2806 ();
 sky130_as_sc_hs__tap_1 TAP_2807 ();
 sky130_as_sc_hs__tap_1 TAP_2808 ();
 sky130_as_sc_hs__tap_1 TAP_2809 ();
 sky130_as_sc_hs__tap_1 TAP_2810 ();
 sky130_as_sc_hs__tap_1 TAP_2811 ();
 sky130_as_sc_hs__tap_1 TAP_2812 ();
 sky130_as_sc_hs__tap_1 TAP_2813 ();
 sky130_as_sc_hs__tap_1 TAP_2814 ();
 sky130_as_sc_hs__tap_1 TAP_2815 ();
 sky130_as_sc_hs__tap_1 TAP_2816 ();
 sky130_as_sc_hs__tap_1 TAP_2817 ();
 sky130_as_sc_hs__tap_1 TAP_2818 ();
 sky130_as_sc_hs__tap_1 TAP_2819 ();
 sky130_as_sc_hs__tap_1 TAP_2820 ();
 sky130_as_sc_hs__tap_1 TAP_2821 ();
 sky130_as_sc_hs__tap_1 TAP_2822 ();
 sky130_as_sc_hs__tap_1 TAP_2823 ();
 sky130_as_sc_hs__tap_1 TAP_2824 ();
 sky130_as_sc_hs__tap_1 TAP_2825 ();
 sky130_as_sc_hs__tap_1 TAP_2826 ();
 sky130_as_sc_hs__tap_1 TAP_2827 ();
 sky130_as_sc_hs__tap_1 TAP_2828 ();
 sky130_as_sc_hs__tap_1 TAP_2829 ();
 sky130_as_sc_hs__tap_1 TAP_2830 ();
 sky130_as_sc_hs__tap_1 TAP_2831 ();
 sky130_as_sc_hs__tap_1 TAP_2832 ();
 sky130_as_sc_hs__tap_1 TAP_2833 ();
 sky130_as_sc_hs__tap_1 TAP_2834 ();
 sky130_as_sc_hs__tap_1 TAP_2835 ();
 sky130_as_sc_hs__tap_1 TAP_2836 ();
 sky130_as_sc_hs__tap_1 TAP_2837 ();
 sky130_as_sc_hs__tap_1 TAP_2838 ();
 sky130_as_sc_hs__tap_1 TAP_2839 ();
 sky130_as_sc_hs__tap_1 TAP_2840 ();
 sky130_as_sc_hs__tap_1 TAP_2841 ();
 sky130_as_sc_hs__tap_1 TAP_2842 ();
 sky130_as_sc_hs__tap_1 TAP_2843 ();
 sky130_as_sc_hs__tap_1 TAP_2844 ();
 sky130_as_sc_hs__tap_1 TAP_2845 ();
 sky130_as_sc_hs__tap_1 TAP_2846 ();
 sky130_as_sc_hs__tap_1 TAP_2847 ();
 sky130_as_sc_hs__tap_1 TAP_2848 ();
 sky130_as_sc_hs__tap_1 TAP_2849 ();
 sky130_as_sc_hs__tap_1 TAP_2850 ();
 sky130_as_sc_hs__tap_1 TAP_2851 ();
 sky130_as_sc_hs__tap_1 TAP_2852 ();
 sky130_as_sc_hs__tap_1 TAP_2853 ();
 sky130_as_sc_hs__tap_1 TAP_2854 ();
 sky130_as_sc_hs__tap_1 TAP_2855 ();
 sky130_as_sc_hs__tap_1 TAP_2856 ();
 sky130_as_sc_hs__tap_1 TAP_2857 ();
 sky130_as_sc_hs__tap_1 TAP_2858 ();
 sky130_as_sc_hs__tap_1 TAP_2859 ();
 sky130_as_sc_hs__tap_1 TAP_2860 ();
 sky130_as_sc_hs__tap_1 TAP_2861 ();
 sky130_as_sc_hs__tap_1 TAP_2862 ();
 sky130_as_sc_hs__tap_1 TAP_2863 ();
 sky130_as_sc_hs__tap_1 TAP_2864 ();
 sky130_as_sc_hs__tap_1 TAP_2865 ();
 sky130_as_sc_hs__tap_1 TAP_2866 ();
 sky130_as_sc_hs__tap_1 TAP_2867 ();
 sky130_as_sc_hs__tap_1 TAP_2868 ();
 sky130_as_sc_hs__tap_1 TAP_2869 ();
 sky130_as_sc_hs__tap_1 TAP_2870 ();
 sky130_as_sc_hs__tap_1 TAP_2871 ();
 sky130_as_sc_hs__tap_1 TAP_2872 ();
 sky130_as_sc_hs__tap_1 TAP_2873 ();
 sky130_as_sc_hs__tap_1 TAP_2874 ();
 sky130_as_sc_hs__tap_1 TAP_2875 ();
 sky130_as_sc_hs__tap_1 TAP_2876 ();
 sky130_as_sc_hs__tap_1 TAP_2877 ();
 sky130_as_sc_hs__tap_1 TAP_2878 ();
 sky130_as_sc_hs__tap_1 TAP_2879 ();
 sky130_as_sc_hs__tap_1 TAP_2880 ();
 sky130_as_sc_hs__tap_1 TAP_2881 ();
 sky130_as_sc_hs__tap_1 TAP_2882 ();
 sky130_as_sc_hs__tap_1 TAP_2883 ();
 sky130_as_sc_hs__tap_1 TAP_2884 ();
 sky130_as_sc_hs__tap_1 TAP_2885 ();
 sky130_as_sc_hs__tap_1 TAP_2886 ();
 sky130_as_sc_hs__tap_1 TAP_2887 ();
 sky130_as_sc_hs__tap_1 TAP_2888 ();
 sky130_as_sc_hs__tap_1 TAP_2889 ();
 sky130_as_sc_hs__tap_1 TAP_2890 ();
 sky130_as_sc_hs__tap_1 TAP_2891 ();
 sky130_as_sc_hs__tap_1 TAP_2892 ();
 sky130_as_sc_hs__tap_1 TAP_2893 ();
 sky130_as_sc_hs__tap_1 TAP_2894 ();
 sky130_as_sc_hs__tap_1 TAP_2895 ();
 sky130_as_sc_hs__tap_1 TAP_2896 ();
 sky130_as_sc_hs__tap_1 TAP_2897 ();
 sky130_as_sc_hs__tap_1 TAP_2898 ();
 sky130_as_sc_hs__tap_1 TAP_2899 ();
 sky130_as_sc_hs__tap_1 TAP_2900 ();
 sky130_as_sc_hs__tap_1 TAP_2901 ();
 sky130_as_sc_hs__tap_1 TAP_2902 ();
 sky130_as_sc_hs__tap_1 TAP_2903 ();
 sky130_as_sc_hs__tap_1 TAP_2904 ();
 sky130_as_sc_hs__tap_1 TAP_2905 ();
 sky130_as_sc_hs__tap_1 TAP_2906 ();
 sky130_as_sc_hs__tap_1 TAP_2907 ();
 sky130_as_sc_hs__tap_1 TAP_2908 ();
 sky130_as_sc_hs__tap_1 TAP_2909 ();
 sky130_as_sc_hs__tap_1 TAP_2910 ();
 sky130_as_sc_hs__tap_1 TAP_2911 ();
 sky130_as_sc_hs__tap_1 TAP_2912 ();
 sky130_as_sc_hs__tap_1 TAP_2913 ();
 sky130_as_sc_hs__tap_1 TAP_2914 ();
 sky130_as_sc_hs__tap_1 TAP_2915 ();
 sky130_as_sc_hs__tap_1 TAP_2916 ();
 sky130_as_sc_hs__tap_1 TAP_2917 ();
 sky130_as_sc_hs__tap_1 TAP_2918 ();
 sky130_as_sc_hs__tap_1 TAP_2919 ();
 sky130_as_sc_hs__tap_1 TAP_2920 ();
 sky130_as_sc_hs__tap_1 TAP_2921 ();
 sky130_as_sc_hs__tap_1 TAP_2922 ();
 sky130_as_sc_hs__tap_1 TAP_2923 ();
 sky130_as_sc_hs__tap_1 TAP_2924 ();
 sky130_as_sc_hs__tap_1 TAP_2925 ();
 sky130_as_sc_hs__tap_1 TAP_2926 ();
 sky130_as_sc_hs__tap_1 TAP_2927 ();
 sky130_as_sc_hs__tap_1 TAP_2928 ();
 sky130_as_sc_hs__tap_1 TAP_2929 ();
 sky130_as_sc_hs__tap_1 TAP_2930 ();
 sky130_as_sc_hs__tap_1 TAP_2931 ();
 sky130_as_sc_hs__tap_1 TAP_2932 ();
 sky130_as_sc_hs__tap_1 TAP_2933 ();
 sky130_as_sc_hs__tap_1 TAP_2934 ();
 sky130_as_sc_hs__tap_1 TAP_2935 ();
 sky130_as_sc_hs__tap_1 TAP_2936 ();
 sky130_as_sc_hs__tap_1 TAP_2937 ();
 sky130_as_sc_hs__tap_1 TAP_2938 ();
 sky130_as_sc_hs__tap_1 TAP_2939 ();
 sky130_as_sc_hs__tap_1 TAP_2940 ();
 sky130_as_sc_hs__tap_1 TAP_2941 ();
 sky130_as_sc_hs__tap_1 TAP_2942 ();
 sky130_as_sc_hs__tap_1 TAP_2943 ();
 sky130_as_sc_hs__tap_1 TAP_2944 ();
 sky130_as_sc_hs__tap_1 TAP_2945 ();
 sky130_as_sc_hs__tap_1 TAP_2946 ();
 sky130_as_sc_hs__tap_1 TAP_2947 ();
 sky130_as_sc_hs__tap_1 TAP_2948 ();
 sky130_as_sc_hs__tap_1 TAP_2949 ();
 sky130_as_sc_hs__tap_1 TAP_2950 ();
 sky130_as_sc_hs__tap_1 TAP_2951 ();
 sky130_as_sc_hs__tap_1 TAP_2952 ();
 sky130_as_sc_hs__tap_1 TAP_2953 ();
 sky130_as_sc_hs__tap_1 TAP_2954 ();
 sky130_as_sc_hs__tap_1 TAP_2955 ();
 sky130_as_sc_hs__tap_1 TAP_2956 ();
 sky130_as_sc_hs__tap_1 TAP_2957 ();
 sky130_as_sc_hs__tap_1 TAP_2958 ();
 sky130_as_sc_hs__tap_1 TAP_2959 ();
 sky130_as_sc_hs__tap_1 TAP_2960 ();
 sky130_as_sc_hs__tap_1 TAP_2961 ();
 sky130_as_sc_hs__tap_1 TAP_2962 ();
 sky130_as_sc_hs__tap_1 TAP_2963 ();
 sky130_as_sc_hs__tap_1 TAP_2964 ();
 sky130_as_sc_hs__tap_1 TAP_2965 ();
 sky130_as_sc_hs__tap_1 TAP_2966 ();
 sky130_as_sc_hs__tap_1 TAP_2967 ();
 sky130_as_sc_hs__tap_1 TAP_2968 ();
 sky130_as_sc_hs__tap_1 TAP_2969 ();
 sky130_as_sc_hs__tap_1 TAP_2970 ();
 sky130_as_sc_hs__tap_1 TAP_2971 ();
 sky130_as_sc_hs__tap_1 TAP_2972 ();
 sky130_as_sc_hs__tap_1 TAP_2973 ();
 sky130_as_sc_hs__tap_1 TAP_2974 ();
 sky130_as_sc_hs__tap_1 TAP_2975 ();
 sky130_as_sc_hs__tap_1 TAP_2976 ();
 sky130_as_sc_hs__tap_1 TAP_2977 ();
 sky130_as_sc_hs__tap_1 TAP_2978 ();
 sky130_as_sc_hs__tap_1 TAP_2979 ();
 sky130_as_sc_hs__tap_1 TAP_2980 ();
 sky130_as_sc_hs__tap_1 TAP_2981 ();
 sky130_as_sc_hs__tap_1 TAP_2982 ();
 sky130_as_sc_hs__tap_1 TAP_2983 ();
 sky130_as_sc_hs__tap_1 TAP_2984 ();
 sky130_as_sc_hs__tap_1 TAP_2985 ();
 sky130_as_sc_hs__tap_1 TAP_2986 ();
 sky130_as_sc_hs__tap_1 TAP_2987 ();
 sky130_as_sc_hs__tap_1 TAP_2988 ();
 sky130_as_sc_hs__tap_1 TAP_2989 ();
 sky130_as_sc_hs__tap_1 TAP_2990 ();
 sky130_as_sc_hs__tap_1 TAP_2991 ();
 sky130_as_sc_hs__tap_1 TAP_2992 ();
 sky130_as_sc_hs__tap_1 TAP_2993 ();
 sky130_as_sc_hs__tap_1 TAP_2994 ();
 sky130_as_sc_hs__tap_1 TAP_2995 ();
 sky130_as_sc_hs__tap_1 TAP_2996 ();
 sky130_as_sc_hs__tap_1 TAP_2997 ();
 sky130_as_sc_hs__tap_1 TAP_2998 ();
 sky130_as_sc_hs__tap_1 TAP_2999 ();
 sky130_as_sc_hs__tap_1 TAP_3000 ();
 sky130_as_sc_hs__tap_1 TAP_3001 ();
 sky130_as_sc_hs__tap_1 TAP_3002 ();
 sky130_as_sc_hs__tap_1 TAP_3003 ();
 sky130_as_sc_hs__tap_1 TAP_3004 ();
 sky130_as_sc_hs__tap_1 TAP_3005 ();
 sky130_as_sc_hs__tap_1 TAP_3006 ();
 sky130_as_sc_hs__tap_1 TAP_3007 ();
 sky130_as_sc_hs__tap_1 TAP_3008 ();
 sky130_as_sc_hs__tap_1 TAP_3009 ();
 sky130_as_sc_hs__tap_1 TAP_3010 ();
 sky130_as_sc_hs__tap_1 TAP_3011 ();
 sky130_as_sc_hs__tap_1 TAP_3012 ();
 sky130_as_sc_hs__tap_1 TAP_3013 ();
 sky130_as_sc_hs__tap_1 TAP_3014 ();
 sky130_as_sc_hs__tap_1 TAP_3015 ();
 sky130_as_sc_hs__tap_1 TAP_3016 ();
 sky130_as_sc_hs__tap_1 TAP_3017 ();
 sky130_as_sc_hs__tap_1 TAP_3018 ();
 sky130_as_sc_hs__tap_1 TAP_3019 ();
 sky130_as_sc_hs__tap_1 TAP_3020 ();
 sky130_as_sc_hs__tap_1 TAP_3021 ();
 sky130_as_sc_hs__tap_1 TAP_3022 ();
 sky130_as_sc_hs__tap_1 TAP_3023 ();
 sky130_as_sc_hs__tap_1 TAP_3024 ();
 sky130_as_sc_hs__tap_1 TAP_3025 ();
 sky130_as_sc_hs__tap_1 TAP_3026 ();
 sky130_as_sc_hs__tap_1 TAP_3027 ();
 sky130_as_sc_hs__tap_1 TAP_3028 ();
 sky130_as_sc_hs__tap_1 TAP_3029 ();
 sky130_as_sc_hs__tap_1 TAP_3030 ();
 sky130_as_sc_hs__tap_1 TAP_3031 ();
 sky130_as_sc_hs__tap_1 TAP_3032 ();
 sky130_as_sc_hs__tap_1 TAP_3033 ();
 sky130_as_sc_hs__tap_1 TAP_3034 ();
 sky130_as_sc_hs__tap_1 TAP_3035 ();
 sky130_as_sc_hs__tap_1 TAP_3036 ();
 sky130_as_sc_hs__tap_1 TAP_3037 ();
 sky130_as_sc_hs__tap_1 TAP_3038 ();
 sky130_as_sc_hs__tap_1 TAP_3039 ();
 sky130_as_sc_hs__tap_1 TAP_3040 ();
 sky130_as_sc_hs__tap_1 TAP_3041 ();
 sky130_as_sc_hs__tap_1 TAP_3042 ();
 sky130_as_sc_hs__tap_1 TAP_3043 ();
 sky130_as_sc_hs__tap_1 TAP_3044 ();
 sky130_as_sc_hs__tap_1 TAP_3045 ();
 sky130_as_sc_hs__tap_1 TAP_3046 ();
 sky130_as_sc_hs__tap_1 TAP_3047 ();
 sky130_as_sc_hs__tap_1 TAP_3048 ();
 sky130_as_sc_hs__tap_1 TAP_3049 ();
 sky130_as_sc_hs__tap_1 TAP_3050 ();
 sky130_as_sc_hs__tap_1 TAP_3051 ();
 sky130_as_sc_hs__tap_1 TAP_3052 ();
 sky130_as_sc_hs__tap_1 TAP_3053 ();
 sky130_as_sc_hs__tap_1 TAP_3054 ();
 sky130_as_sc_hs__tap_1 TAP_3055 ();
 sky130_as_sc_hs__tap_1 TAP_3056 ();
 sky130_as_sc_hs__tap_1 TAP_3057 ();
 sky130_as_sc_hs__tap_1 TAP_3058 ();
 sky130_as_sc_hs__tap_1 TAP_3059 ();
 sky130_as_sc_hs__tap_1 TAP_3060 ();
 sky130_as_sc_hs__tap_1 TAP_3061 ();
 sky130_as_sc_hs__tap_1 TAP_3062 ();
 sky130_as_sc_hs__tap_1 TAP_3063 ();
 sky130_as_sc_hs__tap_1 TAP_3064 ();
 sky130_as_sc_hs__tap_1 TAP_3065 ();
 sky130_as_sc_hs__tap_1 TAP_3066 ();
 sky130_as_sc_hs__tap_1 TAP_3067 ();
 sky130_as_sc_hs__tap_1 TAP_3068 ();
 sky130_as_sc_hs__tap_1 TAP_3069 ();
 sky130_as_sc_hs__tap_1 TAP_3070 ();
 sky130_as_sc_hs__tap_1 TAP_3071 ();
 sky130_as_sc_hs__tap_1 TAP_3072 ();
 sky130_as_sc_hs__tap_1 TAP_3073 ();
 sky130_as_sc_hs__tap_1 TAP_3074 ();
 sky130_as_sc_hs__tap_1 TAP_3075 ();
 sky130_as_sc_hs__tap_1 TAP_3076 ();
 sky130_as_sc_hs__tap_1 TAP_3077 ();
 sky130_as_sc_hs__tap_1 TAP_3078 ();
 sky130_as_sc_hs__tap_1 TAP_3079 ();
 sky130_as_sc_hs__tap_1 TAP_3080 ();
 sky130_as_sc_hs__tap_1 TAP_3081 ();
 sky130_as_sc_hs__tap_1 TAP_3082 ();
 sky130_as_sc_hs__tap_1 TAP_3083 ();
 sky130_as_sc_hs__tap_1 TAP_3084 ();
 sky130_as_sc_hs__tap_1 TAP_3085 ();
 sky130_as_sc_hs__tap_1 TAP_3086 ();
 sky130_as_sc_hs__tap_1 TAP_3087 ();
 sky130_as_sc_hs__tap_1 TAP_3088 ();
 sky130_as_sc_hs__tap_1 TAP_3089 ();
 sky130_as_sc_hs__tap_1 TAP_3090 ();
 sky130_as_sc_hs__tap_1 TAP_3091 ();
 sky130_as_sc_hs__tap_1 TAP_3092 ();
 sky130_as_sc_hs__tap_1 TAP_3093 ();
 sky130_as_sc_hs__tap_1 TAP_3094 ();
 sky130_as_sc_hs__tap_1 TAP_3095 ();
 sky130_as_sc_hs__tap_1 TAP_3096 ();
 sky130_as_sc_hs__tap_1 TAP_3097 ();
 sky130_as_sc_hs__tap_1 TAP_3098 ();
 sky130_as_sc_hs__tap_1 TAP_3099 ();
 sky130_as_sc_hs__tap_1 TAP_3100 ();
 sky130_as_sc_hs__tap_1 TAP_3101 ();
 sky130_as_sc_hs__tap_1 TAP_3102 ();
 sky130_as_sc_hs__tap_1 TAP_3103 ();
 sky130_as_sc_hs__tap_1 TAP_3104 ();
 sky130_as_sc_hs__tap_1 TAP_3105 ();
 sky130_as_sc_hs__tap_1 TAP_3106 ();
 sky130_as_sc_hs__tap_1 TAP_3107 ();
 sky130_as_sc_hs__tap_1 TAP_3108 ();
 sky130_as_sc_hs__tap_1 TAP_3109 ();
 sky130_as_sc_hs__tap_1 TAP_3110 ();
 sky130_as_sc_hs__tap_1 TAP_3111 ();
 sky130_as_sc_hs__tap_1 TAP_3112 ();
 sky130_as_sc_hs__tap_1 TAP_3113 ();
 sky130_as_sc_hs__tap_1 TAP_3114 ();
 sky130_as_sc_hs__tap_1 TAP_3115 ();
 sky130_as_sc_hs__tap_1 TAP_3116 ();
 sky130_as_sc_hs__tap_1 TAP_3117 ();
 sky130_as_sc_hs__tap_1 TAP_3118 ();
 sky130_as_sc_hs__tap_1 TAP_3119 ();
 sky130_as_sc_hs__tap_1 TAP_3120 ();
 sky130_as_sc_hs__tap_1 TAP_3121 ();
 sky130_as_sc_hs__tap_1 TAP_3122 ();
 sky130_as_sc_hs__tap_1 TAP_3123 ();
 sky130_as_sc_hs__tap_1 TAP_3124 ();
 sky130_as_sc_hs__tap_1 TAP_3125 ();
 sky130_as_sc_hs__tap_1 TAP_3126 ();
 sky130_as_sc_hs__tap_1 TAP_3127 ();
 sky130_as_sc_hs__tap_1 TAP_3128 ();
 sky130_as_sc_hs__tap_1 TAP_3129 ();
 sky130_as_sc_hs__tap_1 TAP_3130 ();
 sky130_as_sc_hs__tap_1 TAP_3131 ();
 sky130_as_sc_hs__tap_1 TAP_3132 ();
 sky130_as_sc_hs__tap_1 TAP_3133 ();
 sky130_as_sc_hs__tap_1 TAP_3134 ();
 sky130_as_sc_hs__tap_1 TAP_3135 ();
 sky130_as_sc_hs__tap_1 TAP_3136 ();
 sky130_as_sc_hs__tap_1 TAP_3137 ();
 sky130_as_sc_hs__tap_1 TAP_3138 ();
 sky130_as_sc_hs__tap_1 TAP_3139 ();
 sky130_as_sc_hs__tap_1 TAP_3140 ();
 sky130_as_sc_hs__tap_1 TAP_3141 ();
 sky130_as_sc_hs__tap_1 TAP_3142 ();
 sky130_as_sc_hs__tap_1 TAP_3143 ();
 sky130_as_sc_hs__tap_1 TAP_3144 ();
 sky130_as_sc_hs__tap_1 TAP_3145 ();
 sky130_as_sc_hs__tap_1 TAP_3146 ();
 sky130_as_sc_hs__tap_1 TAP_3147 ();
 sky130_as_sc_hs__tap_1 TAP_3148 ();
 sky130_as_sc_hs__tap_1 TAP_3149 ();
 sky130_as_sc_hs__tap_1 TAP_3150 ();
 sky130_as_sc_hs__tap_1 TAP_3151 ();
 sky130_as_sc_hs__tap_1 TAP_3152 ();
 sky130_as_sc_hs__tap_1 TAP_3153 ();
 sky130_as_sc_hs__tap_1 TAP_3154 ();
 sky130_as_sc_hs__tap_1 TAP_3155 ();
 sky130_as_sc_hs__tap_1 TAP_3156 ();
 sky130_as_sc_hs__tap_1 TAP_3157 ();
 sky130_as_sc_hs__tap_1 TAP_3158 ();
 sky130_as_sc_hs__tap_1 TAP_3159 ();
 sky130_as_sc_hs__tap_1 TAP_3160 ();
 sky130_as_sc_hs__tap_1 TAP_3161 ();
 sky130_as_sc_hs__tap_1 TAP_3162 ();
 sky130_as_sc_hs__tap_1 TAP_3163 ();
 sky130_as_sc_hs__tap_1 TAP_3164 ();
 sky130_as_sc_hs__tap_1 TAP_3165 ();
 sky130_as_sc_hs__tap_1 TAP_3166 ();
 sky130_as_sc_hs__tap_1 TAP_3167 ();
 sky130_as_sc_hs__tap_1 TAP_3168 ();
 sky130_as_sc_hs__tap_1 TAP_3169 ();
 sky130_as_sc_hs__tap_1 TAP_3170 ();
 sky130_as_sc_hs__tap_1 TAP_3171 ();
 sky130_as_sc_hs__tap_1 TAP_3172 ();
 sky130_as_sc_hs__tap_1 TAP_3173 ();
 sky130_as_sc_hs__tap_1 TAP_3174 ();
 sky130_as_sc_hs__tap_1 TAP_3175 ();
 sky130_as_sc_hs__tap_1 TAP_3176 ();
 sky130_as_sc_hs__tap_1 TAP_3177 ();
 sky130_as_sc_hs__tap_1 TAP_3178 ();
 sky130_as_sc_hs__tap_1 TAP_3179 ();
 sky130_as_sc_hs__tap_1 TAP_3180 ();
 sky130_as_sc_hs__tap_1 TAP_3181 ();
 sky130_as_sc_hs__tap_1 TAP_3182 ();
 sky130_as_sc_hs__tap_1 TAP_3183 ();
 sky130_as_sc_hs__tap_1 TAP_3184 ();
 sky130_as_sc_hs__tap_1 TAP_3185 ();
 sky130_as_sc_hs__tap_1 TAP_3186 ();
 sky130_as_sc_hs__tap_1 TAP_3187 ();
 sky130_as_sc_hs__tap_1 TAP_3188 ();
 sky130_as_sc_hs__tap_1 TAP_3189 ();
 sky130_as_sc_hs__tap_1 TAP_3190 ();
 sky130_as_sc_hs__tap_1 TAP_3191 ();
 sky130_as_sc_hs__tap_1 TAP_3192 ();
 sky130_as_sc_hs__tap_1 TAP_3193 ();
 sky130_as_sc_hs__tap_1 TAP_3194 ();
 sky130_as_sc_hs__tap_1 TAP_3195 ();
 sky130_as_sc_hs__tap_1 TAP_3196 ();
 sky130_as_sc_hs__tap_1 TAP_3197 ();
 sky130_as_sc_hs__tap_1 TAP_3198 ();
 sky130_as_sc_hs__tap_1 TAP_3199 ();
 sky130_as_sc_hs__tap_1 TAP_3200 ();
 sky130_as_sc_hs__tap_1 TAP_3201 ();
 sky130_as_sc_hs__tap_1 TAP_3202 ();
 sky130_as_sc_hs__tap_1 TAP_3203 ();
 sky130_as_sc_hs__tap_1 TAP_3204 ();
 sky130_as_sc_hs__tap_1 TAP_3205 ();
 sky130_as_sc_hs__tap_1 TAP_3206 ();
 sky130_as_sc_hs__tap_1 TAP_3207 ();
 sky130_as_sc_hs__tap_1 TAP_3208 ();
 sky130_as_sc_hs__tap_1 TAP_3209 ();
 sky130_as_sc_hs__tap_1 TAP_3210 ();
 sky130_as_sc_hs__tap_1 TAP_3211 ();
 sky130_as_sc_hs__tap_1 TAP_3212 ();
 sky130_as_sc_hs__tap_1 TAP_3213 ();
 sky130_as_sc_hs__tap_1 TAP_3214 ();
 sky130_as_sc_hs__tap_1 TAP_3215 ();
 sky130_as_sc_hs__tap_1 TAP_3216 ();
 sky130_as_sc_hs__tap_1 TAP_3217 ();
 sky130_as_sc_hs__tap_1 TAP_3218 ();
 sky130_as_sc_hs__tap_1 TAP_3219 ();
 sky130_as_sc_hs__tap_1 TAP_3220 ();
 sky130_as_sc_hs__tap_1 TAP_3221 ();
 sky130_as_sc_hs__tap_1 TAP_3222 ();
 sky130_as_sc_hs__tap_1 TAP_3223 ();
 sky130_as_sc_hs__tap_1 TAP_3224 ();
 sky130_as_sc_hs__tap_1 TAP_3225 ();
 sky130_as_sc_hs__tap_1 TAP_3226 ();
 sky130_as_sc_hs__tap_1 TAP_3227 ();
 sky130_as_sc_hs__tap_1 TAP_3228 ();
 sky130_as_sc_hs__tap_1 TAP_3229 ();
 sky130_as_sc_hs__tap_1 TAP_3230 ();
 sky130_as_sc_hs__tap_1 TAP_3231 ();
 sky130_as_sc_hs__tap_1 TAP_3232 ();
 sky130_as_sc_hs__tap_1 TAP_3233 ();
 sky130_as_sc_hs__tap_1 TAP_3234 ();
 sky130_as_sc_hs__tap_1 TAP_3235 ();
 sky130_as_sc_hs__tap_1 TAP_3236 ();
 sky130_as_sc_hs__tap_1 TAP_3237 ();
 sky130_as_sc_hs__tap_1 TAP_3238 ();
 sky130_as_sc_hs__tap_1 TAP_3239 ();
 sky130_as_sc_hs__tap_1 TAP_3240 ();
 sky130_as_sc_hs__tap_1 TAP_3241 ();
 sky130_as_sc_hs__tap_1 TAP_3242 ();
 sky130_as_sc_hs__tap_1 TAP_3243 ();
 sky130_as_sc_hs__tap_1 TAP_3244 ();
 sky130_as_sc_hs__tap_1 TAP_3245 ();
 sky130_as_sc_hs__tap_1 TAP_3246 ();
 sky130_as_sc_hs__tap_1 TAP_3247 ();
 sky130_as_sc_hs__tap_1 TAP_3248 ();
 sky130_as_sc_hs__tap_1 TAP_3249 ();
 sky130_as_sc_hs__tap_1 TAP_3250 ();
 sky130_as_sc_hs__tap_1 TAP_3251 ();
 sky130_as_sc_hs__tap_1 TAP_3252 ();
 sky130_as_sc_hs__tap_1 TAP_3253 ();
 sky130_as_sc_hs__tap_1 TAP_3254 ();
 sky130_as_sc_hs__tap_1 TAP_3255 ();
 sky130_as_sc_hs__tap_1 TAP_3256 ();
 sky130_as_sc_hs__tap_1 TAP_3257 ();
 sky130_as_sc_hs__tap_1 TAP_3258 ();
 sky130_as_sc_hs__tap_1 TAP_3259 ();
 sky130_as_sc_hs__tap_1 TAP_3260 ();
 sky130_as_sc_hs__tap_1 TAP_3261 ();
 sky130_as_sc_hs__tap_1 TAP_3262 ();
 sky130_as_sc_hs__tap_1 TAP_3263 ();
 sky130_as_sc_hs__tap_1 TAP_3264 ();
 sky130_as_sc_hs__tap_1 TAP_3265 ();
 sky130_as_sc_hs__tap_1 TAP_3266 ();
 sky130_as_sc_hs__tap_1 TAP_3267 ();
 sky130_as_sc_hs__tap_1 TAP_3268 ();
 sky130_as_sc_hs__tap_1 TAP_3269 ();
 sky130_as_sc_hs__tap_1 TAP_3270 ();
 sky130_as_sc_hs__tap_1 TAP_3271 ();
 sky130_as_sc_hs__tap_1 TAP_3272 ();
 sky130_as_sc_hs__tap_1 TAP_3273 ();
 sky130_as_sc_hs__tap_1 TAP_3274 ();
 sky130_as_sc_hs__tap_1 TAP_3275 ();
 sky130_as_sc_hs__tap_1 TAP_3276 ();
 sky130_as_sc_hs__tap_1 TAP_3277 ();
 sky130_as_sc_hs__tap_1 TAP_3278 ();
 sky130_as_sc_hs__tap_1 TAP_3279 ();
 sky130_as_sc_hs__tap_1 TAP_3280 ();
 sky130_as_sc_hs__tap_1 TAP_3281 ();
 sky130_as_sc_hs__tap_1 TAP_3282 ();
 sky130_as_sc_hs__tap_1 TAP_3283 ();
 sky130_as_sc_hs__tap_1 TAP_3284 ();
 sky130_as_sc_hs__tap_1 TAP_3285 ();
 sky130_as_sc_hs__tap_1 TAP_3286 ();
 sky130_as_sc_hs__tap_1 TAP_3287 ();
 sky130_as_sc_hs__tap_1 TAP_3288 ();
 sky130_as_sc_hs__tap_1 TAP_3289 ();
 sky130_as_sc_hs__tap_1 TAP_3290 ();
 sky130_as_sc_hs__tap_1 TAP_3291 ();
 sky130_as_sc_hs__tap_1 TAP_3292 ();
 sky130_as_sc_hs__tap_1 TAP_3293 ();
 sky130_as_sc_hs__tap_1 TAP_3294 ();
 sky130_as_sc_hs__tap_1 TAP_3295 ();
 sky130_as_sc_hs__tap_1 TAP_3296 ();
 sky130_as_sc_hs__tap_1 TAP_3297 ();
 sky130_as_sc_hs__tap_1 TAP_3298 ();
 sky130_as_sc_hs__tap_1 TAP_3299 ();
 sky130_as_sc_hs__tap_1 TAP_3300 ();
 sky130_as_sc_hs__tap_1 TAP_3301 ();
 sky130_as_sc_hs__tap_1 TAP_3302 ();
 sky130_as_sc_hs__tap_1 TAP_3303 ();
 sky130_as_sc_hs__tap_1 TAP_3304 ();
 sky130_as_sc_hs__tap_1 TAP_3305 ();
 sky130_as_sc_hs__tap_1 TAP_3306 ();
 sky130_as_sc_hs__tap_1 TAP_3307 ();
 sky130_as_sc_hs__tap_1 TAP_3308 ();
 sky130_as_sc_hs__tap_1 TAP_3309 ();
 sky130_as_sc_hs__tap_1 TAP_3310 ();
 sky130_as_sc_hs__tap_1 TAP_3311 ();
 sky130_as_sc_hs__tap_1 TAP_3312 ();
 sky130_as_sc_hs__tap_1 TAP_3313 ();
 sky130_as_sc_hs__tap_1 TAP_3314 ();
 sky130_as_sc_hs__tap_1 TAP_3315 ();
 sky130_as_sc_hs__tap_1 TAP_3316 ();
 sky130_as_sc_hs__tap_1 TAP_3317 ();
 sky130_as_sc_hs__tap_1 TAP_3318 ();
 sky130_as_sc_hs__tap_1 TAP_3319 ();
 sky130_as_sc_hs__tap_1 TAP_3320 ();
 sky130_as_sc_hs__tap_1 TAP_3321 ();
 sky130_as_sc_hs__tap_1 TAP_3322 ();
 sky130_as_sc_hs__tap_1 TAP_3323 ();
 sky130_as_sc_hs__tap_1 TAP_3324 ();
 sky130_as_sc_hs__tap_1 TAP_3325 ();
 sky130_as_sc_hs__tap_1 TAP_3326 ();
 sky130_as_sc_hs__tap_1 TAP_3327 ();
 sky130_as_sc_hs__tap_1 TAP_3328 ();
 sky130_as_sc_hs__tap_1 TAP_3329 ();
 sky130_as_sc_hs__tap_1 TAP_3330 ();
 sky130_as_sc_hs__tap_1 TAP_3331 ();
 sky130_as_sc_hs__tap_1 TAP_3332 ();
 sky130_as_sc_hs__tap_1 TAP_3333 ();
 sky130_as_sc_hs__tap_1 TAP_3334 ();
 sky130_as_sc_hs__tap_1 TAP_3335 ();
 sky130_as_sc_hs__tap_1 TAP_3336 ();
 sky130_as_sc_hs__tap_1 TAP_3337 ();
 sky130_as_sc_hs__tap_1 TAP_3338 ();
 sky130_as_sc_hs__tap_1 TAP_3339 ();
 sky130_as_sc_hs__tap_1 TAP_3340 ();
 sky130_as_sc_hs__tap_1 TAP_3341 ();
 sky130_as_sc_hs__tap_1 TAP_3342 ();
 sky130_as_sc_hs__tap_1 TAP_3343 ();
 sky130_as_sc_hs__tap_1 TAP_3344 ();
 sky130_as_sc_hs__tap_1 TAP_3345 ();
 sky130_as_sc_hs__tap_1 TAP_3346 ();
 sky130_as_sc_hs__tap_1 TAP_3347 ();
 sky130_as_sc_hs__tap_1 TAP_3348 ();
 sky130_as_sc_hs__tap_1 TAP_3349 ();
 sky130_as_sc_hs__tap_1 TAP_3350 ();
 sky130_as_sc_hs__tap_1 TAP_3351 ();
 sky130_as_sc_hs__tap_1 TAP_3352 ();
 sky130_as_sc_hs__tap_1 TAP_3353 ();
 sky130_as_sc_hs__tap_1 TAP_3354 ();
 sky130_as_sc_hs__tap_1 TAP_3355 ();
 sky130_as_sc_hs__tap_1 TAP_3356 ();
 sky130_as_sc_hs__tap_1 TAP_3357 ();
 sky130_as_sc_hs__tap_1 TAP_3358 ();
 sky130_as_sc_hs__tap_1 TAP_3359 ();
 sky130_as_sc_hs__tap_1 TAP_3360 ();
 sky130_as_sc_hs__tap_1 TAP_3361 ();
 sky130_as_sc_hs__tap_1 TAP_3362 ();
 sky130_as_sc_hs__tap_1 TAP_3363 ();
 sky130_as_sc_hs__tap_1 TAP_3364 ();
 sky130_as_sc_hs__tap_1 TAP_3365 ();
 sky130_as_sc_hs__tap_1 TAP_3366 ();
 sky130_as_sc_hs__tap_1 TAP_3367 ();
 sky130_as_sc_hs__tap_1 TAP_3368 ();
 sky130_as_sc_hs__tap_1 TAP_3369 ();
 sky130_as_sc_hs__tap_1 TAP_3370 ();
 sky130_as_sc_hs__tap_1 TAP_3371 ();
 sky130_as_sc_hs__tap_1 TAP_3372 ();
 sky130_as_sc_hs__tap_1 TAP_3373 ();
 sky130_as_sc_hs__tap_1 TAP_3374 ();
 sky130_as_sc_hs__tap_1 TAP_3375 ();
 sky130_as_sc_hs__tap_1 TAP_3376 ();
 sky130_as_sc_hs__tap_1 TAP_3377 ();
 sky130_as_sc_hs__tap_1 TAP_3378 ();
 sky130_as_sc_hs__tap_1 TAP_3379 ();
 sky130_as_sc_hs__tap_1 TAP_3380 ();
 sky130_as_sc_hs__tap_1 TAP_3381 ();
 sky130_as_sc_hs__tap_1 TAP_3382 ();
 sky130_as_sc_hs__tap_1 TAP_3383 ();
 sky130_as_sc_hs__tap_1 TAP_3384 ();
 sky130_as_sc_hs__tap_1 TAP_3385 ();
 sky130_as_sc_hs__tap_1 TAP_3386 ();
 sky130_as_sc_hs__tap_1 TAP_3387 ();
 sky130_as_sc_hs__tap_1 TAP_3388 ();
 sky130_as_sc_hs__tap_1 TAP_3389 ();
 sky130_as_sc_hs__tap_1 TAP_3390 ();
 sky130_as_sc_hs__tap_1 TAP_3391 ();
 sky130_as_sc_hs__tap_1 TAP_3392 ();
 sky130_as_sc_hs__tap_1 TAP_3393 ();
 sky130_as_sc_hs__tap_1 TAP_3394 ();
 sky130_as_sc_hs__tap_1 TAP_3395 ();
 sky130_as_sc_hs__tap_1 TAP_3396 ();
 sky130_as_sc_hs__tap_1 TAP_3397 ();
 sky130_as_sc_hs__tap_1 TAP_3398 ();
 sky130_as_sc_hs__tap_1 TAP_3399 ();
 sky130_as_sc_hs__tap_1 TAP_3400 ();
 sky130_as_sc_hs__tap_1 TAP_3401 ();
 sky130_as_sc_hs__tap_1 TAP_3402 ();
 sky130_as_sc_hs__tap_1 TAP_3403 ();
 sky130_as_sc_hs__tap_1 TAP_3404 ();
 sky130_as_sc_hs__tap_1 TAP_3405 ();
 sky130_as_sc_hs__tap_1 TAP_3406 ();
 sky130_as_sc_hs__tap_1 TAP_3407 ();
 sky130_as_sc_hs__tap_1 TAP_3408 ();
 sky130_as_sc_hs__tap_1 TAP_3409 ();
 sky130_as_sc_hs__tap_1 TAP_3410 ();
 sky130_as_sc_hs__tap_1 TAP_3411 ();
 sky130_as_sc_hs__tap_1 TAP_3412 ();
 sky130_as_sc_hs__tap_1 TAP_3413 ();
 sky130_as_sc_hs__tap_1 TAP_3414 ();
 sky130_as_sc_hs__tap_1 TAP_3415 ();
 sky130_as_sc_hs__tap_1 TAP_3416 ();
 sky130_as_sc_hs__tap_1 TAP_3417 ();
 sky130_as_sc_hs__tap_1 TAP_3418 ();
 sky130_as_sc_hs__tap_1 TAP_3419 ();
 sky130_as_sc_hs__tap_1 TAP_3420 ();
 sky130_as_sc_hs__tap_1 TAP_3421 ();
 sky130_as_sc_hs__tap_1 TAP_3422 ();
 sky130_as_sc_hs__tap_1 TAP_3423 ();
 sky130_as_sc_hs__tap_1 TAP_3424 ();
 sky130_as_sc_hs__tap_1 TAP_3425 ();
 sky130_as_sc_hs__tap_1 TAP_3426 ();
 sky130_as_sc_hs__tap_1 TAP_3427 ();
 sky130_as_sc_hs__tap_1 TAP_3428 ();
 sky130_as_sc_hs__tap_1 TAP_3429 ();
 sky130_as_sc_hs__tap_1 TAP_3430 ();
 sky130_as_sc_hs__tap_1 TAP_3431 ();
 sky130_as_sc_hs__tap_1 TAP_3432 ();
 sky130_as_sc_hs__tap_1 TAP_3433 ();
 sky130_as_sc_hs__tap_1 TAP_3434 ();
 sky130_as_sc_hs__tap_1 TAP_3435 ();
 sky130_as_sc_hs__tap_1 TAP_3436 ();
 sky130_as_sc_hs__tap_1 TAP_3437 ();
 sky130_as_sc_hs__tap_1 TAP_3438 ();
 sky130_as_sc_hs__tap_1 TAP_3439 ();
 sky130_as_sc_hs__tap_1 TAP_3440 ();
 sky130_as_sc_hs__tap_1 TAP_3441 ();
 sky130_as_sc_hs__tap_1 TAP_3442 ();
 sky130_as_sc_hs__tap_1 TAP_3443 ();
 sky130_as_sc_hs__tap_1 TAP_3444 ();
 sky130_as_sc_hs__tap_1 TAP_3445 ();
 sky130_as_sc_hs__tap_1 TAP_3446 ();
 sky130_as_sc_hs__tap_1 TAP_3447 ();
 sky130_as_sc_hs__tap_1 TAP_3448 ();
 sky130_as_sc_hs__tap_1 TAP_3449 ();
 sky130_as_sc_hs__tap_1 TAP_3450 ();
 sky130_as_sc_hs__tap_1 TAP_3451 ();
 sky130_as_sc_hs__tap_1 TAP_3452 ();
 sky130_as_sc_hs__tap_1 TAP_3453 ();
 sky130_as_sc_hs__tap_1 TAP_3454 ();
 sky130_as_sc_hs__tap_1 TAP_3455 ();
 sky130_as_sc_hs__tap_1 TAP_3456 ();
 sky130_as_sc_hs__tap_1 TAP_3457 ();
 sky130_as_sc_hs__tap_1 TAP_3458 ();
 sky130_as_sc_hs__tap_1 TAP_3459 ();
 sky130_as_sc_hs__tap_1 TAP_3460 ();
 sky130_as_sc_hs__tap_1 TAP_3461 ();
 sky130_as_sc_hs__tap_1 TAP_3462 ();
 sky130_as_sc_hs__tap_1 TAP_3463 ();
 sky130_as_sc_hs__tap_1 TAP_3464 ();
 sky130_as_sc_hs__tap_1 TAP_3465 ();
 sky130_as_sc_hs__tap_1 TAP_3466 ();
 sky130_as_sc_hs__tap_1 TAP_3467 ();
 sky130_as_sc_hs__tap_1 TAP_3468 ();
 sky130_as_sc_hs__tap_1 TAP_3469 ();
 sky130_as_sc_hs__tap_1 TAP_3470 ();
 sky130_as_sc_hs__tap_1 TAP_3471 ();
 sky130_as_sc_hs__tap_1 TAP_3472 ();
 sky130_as_sc_hs__tap_1 TAP_3473 ();
 sky130_as_sc_hs__tap_1 TAP_3474 ();
 sky130_as_sc_hs__tap_1 TAP_3475 ();
 sky130_as_sc_hs__tap_1 TAP_3476 ();
 sky130_as_sc_hs__tap_1 TAP_3477 ();
 sky130_as_sc_hs__tap_1 TAP_3478 ();
 sky130_as_sc_hs__tap_1 TAP_3479 ();
 sky130_as_sc_hs__tap_1 TAP_3480 ();
 sky130_as_sc_hs__tap_1 TAP_3481 ();
 sky130_as_sc_hs__tap_1 TAP_3482 ();
 sky130_as_sc_hs__tap_1 TAP_3483 ();
 sky130_as_sc_hs__tap_1 TAP_3484 ();
 sky130_as_sc_hs__tap_1 TAP_3485 ();
 sky130_as_sc_hs__tap_1 TAP_3486 ();
 sky130_as_sc_hs__tap_1 TAP_3487 ();
 sky130_as_sc_hs__tap_1 TAP_3488 ();
 sky130_as_sc_hs__tap_1 TAP_3489 ();
 sky130_as_sc_hs__tap_1 TAP_3490 ();
 sky130_as_sc_hs__tap_1 TAP_3491 ();
 sky130_as_sc_hs__tap_1 TAP_3492 ();
 sky130_as_sc_hs__tap_1 TAP_3493 ();
 sky130_as_sc_hs__tap_1 TAP_3494 ();
 sky130_as_sc_hs__tap_1 TAP_3495 ();
 sky130_as_sc_hs__tap_1 TAP_3496 ();
 sky130_as_sc_hs__tap_1 TAP_3497 ();
 sky130_as_sc_hs__tap_1 TAP_3498 ();
 sky130_as_sc_hs__tap_1 TAP_3499 ();
 sky130_as_sc_hs__tap_1 TAP_3500 ();
 sky130_as_sc_hs__tap_1 TAP_3501 ();
 sky130_as_sc_hs__tap_1 TAP_3502 ();
 sky130_as_sc_hs__tap_1 TAP_3503 ();
 sky130_as_sc_hs__tap_1 TAP_3504 ();
 sky130_as_sc_hs__tap_1 TAP_3505 ();
 sky130_as_sc_hs__tap_1 TAP_3506 ();
 sky130_as_sc_hs__tap_1 TAP_3507 ();
 sky130_as_sc_hs__tap_1 TAP_3508 ();
 sky130_as_sc_hs__tap_1 TAP_3509 ();
 sky130_as_sc_hs__tap_1 TAP_3510 ();
 sky130_as_sc_hs__tap_1 TAP_3511 ();
 sky130_as_sc_hs__tap_1 TAP_3512 ();
 sky130_as_sc_hs__tap_1 TAP_3513 ();
 sky130_as_sc_hs__tap_1 TAP_3514 ();
 sky130_as_sc_hs__tap_1 TAP_3515 ();
 sky130_as_sc_hs__tap_1 TAP_3516 ();
 sky130_as_sc_hs__tap_1 TAP_3517 ();
 sky130_as_sc_hs__tap_1 TAP_3518 ();
 sky130_as_sc_hs__tap_1 TAP_3519 ();
 sky130_as_sc_hs__tap_1 TAP_3520 ();
 sky130_as_sc_hs__tap_1 TAP_3521 ();
 sky130_as_sc_hs__tap_1 TAP_3522 ();
 sky130_as_sc_hs__tap_1 TAP_3523 ();
 sky130_as_sc_hs__tap_1 TAP_3524 ();
 sky130_as_sc_hs__tap_1 TAP_3525 ();
 sky130_as_sc_hs__tap_1 TAP_3526 ();
 sky130_as_sc_hs__tap_1 TAP_3527 ();
 sky130_as_sc_hs__tap_1 TAP_3528 ();
 sky130_as_sc_hs__tap_1 TAP_3529 ();
 sky130_as_sc_hs__tap_1 TAP_3530 ();
 sky130_as_sc_hs__tap_1 TAP_3531 ();
 sky130_as_sc_hs__tap_1 TAP_3532 ();
 sky130_as_sc_hs__tap_1 TAP_3533 ();
 sky130_as_sc_hs__tap_1 TAP_3534 ();
 sky130_as_sc_hs__tap_1 TAP_3535 ();
 sky130_as_sc_hs__tap_1 TAP_3536 ();
 sky130_as_sc_hs__tap_1 TAP_3537 ();
 sky130_as_sc_hs__tap_1 TAP_3538 ();
 sky130_as_sc_hs__tap_1 TAP_3539 ();
 sky130_as_sc_hs__tap_1 TAP_3540 ();
 sky130_as_sc_hs__tap_1 TAP_3541 ();
 sky130_as_sc_hs__tap_1 TAP_3542 ();
 sky130_as_sc_hs__tap_1 TAP_3543 ();
 sky130_as_sc_hs__tap_1 TAP_3544 ();
 sky130_as_sc_hs__tap_1 TAP_3545 ();
 sky130_as_sc_hs__tap_1 TAP_3546 ();
 sky130_as_sc_hs__tap_1 TAP_3547 ();
 sky130_as_sc_hs__tap_1 TAP_3548 ();
 sky130_as_sc_hs__tap_1 TAP_3549 ();
 sky130_as_sc_hs__tap_1 TAP_3550 ();
 sky130_as_sc_hs__tap_1 TAP_3551 ();
 sky130_as_sc_hs__tap_1 TAP_3552 ();
 sky130_as_sc_hs__tap_1 TAP_3553 ();
 sky130_as_sc_hs__tap_1 TAP_3554 ();
 sky130_as_sc_hs__tap_1 TAP_3555 ();
 sky130_as_sc_hs__tap_1 TAP_3556 ();
 sky130_as_sc_hs__tap_1 TAP_3557 ();
 sky130_as_sc_hs__tap_1 TAP_3558 ();
 sky130_as_sc_hs__tap_1 TAP_3559 ();
 sky130_as_sc_hs__tap_1 TAP_3560 ();
 sky130_as_sc_hs__tap_1 TAP_3561 ();
 sky130_as_sc_hs__tap_1 TAP_3562 ();
 sky130_as_sc_hs__tap_1 TAP_3563 ();
 sky130_as_sc_hs__tap_1 TAP_3564 ();
 sky130_as_sc_hs__tap_1 TAP_3565 ();
 sky130_as_sc_hs__tap_1 TAP_3566 ();
 sky130_as_sc_hs__tap_1 TAP_3567 ();
 sky130_as_sc_hs__tap_1 TAP_3568 ();
 sky130_as_sc_hs__tap_1 TAP_3569 ();
 sky130_as_sc_hs__tap_1 TAP_3570 ();
 sky130_as_sc_hs__tap_1 TAP_3571 ();
 sky130_as_sc_hs__tap_1 TAP_3572 ();
 sky130_as_sc_hs__tap_1 TAP_3573 ();
 sky130_as_sc_hs__tap_1 TAP_3574 ();
 sky130_as_sc_hs__tap_1 TAP_3575 ();
 sky130_as_sc_hs__tap_1 TAP_3576 ();
 sky130_as_sc_hs__tap_1 TAP_3577 ();
 sky130_as_sc_hs__tap_1 TAP_3578 ();
 sky130_as_sc_hs__tap_1 TAP_3579 ();
 sky130_as_sc_hs__tap_1 TAP_3580 ();
 sky130_as_sc_hs__tap_1 TAP_3581 ();
 sky130_as_sc_hs__tap_1 TAP_3582 ();
 sky130_as_sc_hs__tap_1 TAP_3583 ();
 sky130_as_sc_hs__tap_1 TAP_3584 ();
 sky130_as_sc_hs__tap_1 TAP_3585 ();
 sky130_as_sc_hs__tap_1 TAP_3586 ();
 sky130_as_sc_hs__tap_1 TAP_3587 ();
 sky130_as_sc_hs__tap_1 TAP_3588 ();
 sky130_as_sc_hs__tap_1 TAP_3589 ();
 sky130_as_sc_hs__tap_1 TAP_3590 ();
 sky130_as_sc_hs__tap_1 TAP_3591 ();
 sky130_as_sc_hs__tap_1 TAP_3592 ();
 sky130_as_sc_hs__tap_1 TAP_3593 ();
 sky130_as_sc_hs__tap_1 TAP_3594 ();
 sky130_as_sc_hs__tap_1 TAP_3595 ();
 sky130_as_sc_hs__tap_1 TAP_3596 ();
 sky130_as_sc_hs__tap_1 TAP_3597 ();
 sky130_as_sc_hs__tap_1 TAP_3598 ();
 sky130_as_sc_hs__tap_1 TAP_3599 ();
 sky130_as_sc_hs__tap_1 TAP_3600 ();
 sky130_as_sc_hs__tap_1 TAP_3601 ();
 sky130_as_sc_hs__tap_1 TAP_3602 ();
 sky130_as_sc_hs__tap_1 TAP_3603 ();
 sky130_as_sc_hs__tap_1 TAP_3604 ();
 sky130_as_sc_hs__tap_1 TAP_3605 ();
 sky130_as_sc_hs__tap_1 TAP_3606 ();
 sky130_as_sc_hs__tap_1 TAP_3607 ();
 sky130_as_sc_hs__tap_1 TAP_3608 ();
 sky130_as_sc_hs__tap_1 TAP_3609 ();
 sky130_as_sc_hs__tap_1 TAP_3610 ();
 sky130_as_sc_hs__tap_1 TAP_3611 ();
 sky130_as_sc_hs__tap_1 TAP_3612 ();
 sky130_as_sc_hs__tap_1 TAP_3613 ();
 sky130_as_sc_hs__tap_1 TAP_3614 ();
 sky130_as_sc_hs__tap_1 TAP_3615 ();
 sky130_as_sc_hs__tap_1 TAP_3616 ();
 sky130_as_sc_hs__tap_1 TAP_3617 ();
 sky130_as_sc_hs__tap_1 TAP_3618 ();
 sky130_as_sc_hs__tap_1 TAP_3619 ();
 sky130_as_sc_hs__tap_1 TAP_3620 ();
 sky130_as_sc_hs__tap_1 TAP_3621 ();
 sky130_as_sc_hs__tap_1 TAP_3622 ();
 sky130_as_sc_hs__tap_1 TAP_3623 ();
 sky130_as_sc_hs__tap_1 TAP_3624 ();
 sky130_as_sc_hs__tap_1 TAP_3625 ();
 sky130_as_sc_hs__tap_1 TAP_3626 ();
 sky130_as_sc_hs__tap_1 TAP_3627 ();
 sky130_as_sc_hs__tap_1 TAP_3628 ();
 sky130_as_sc_hs__tap_1 TAP_3629 ();
 sky130_as_sc_hs__tap_1 TAP_3630 ();
 sky130_as_sc_hs__tap_1 TAP_3631 ();
 sky130_as_sc_hs__tap_1 TAP_3632 ();
 sky130_as_sc_hs__tap_1 TAP_3633 ();
 sky130_as_sc_hs__tap_1 TAP_3634 ();
 sky130_as_sc_hs__tap_1 TAP_3635 ();
 sky130_as_sc_hs__tap_1 TAP_3636 ();
 sky130_as_sc_hs__tap_1 TAP_3637 ();
 sky130_as_sc_hs__tap_1 TAP_3638 ();
 sky130_as_sc_hs__tap_1 TAP_3639 ();
 sky130_as_sc_hs__tap_1 TAP_3640 ();
 sky130_as_sc_hs__tap_1 TAP_3641 ();
 sky130_as_sc_hs__tap_1 TAP_3642 ();
 sky130_as_sc_hs__tap_1 TAP_3643 ();
 sky130_as_sc_hs__tap_1 TAP_3644 ();
 sky130_as_sc_hs__tap_1 TAP_3645 ();
 sky130_as_sc_hs__tap_1 TAP_3646 ();
 sky130_as_sc_hs__tap_1 TAP_3647 ();
 sky130_as_sc_hs__tap_1 TAP_3648 ();
 sky130_as_sc_hs__tap_1 TAP_3649 ();
 sky130_as_sc_hs__tap_1 TAP_3650 ();
 sky130_as_sc_hs__tap_1 TAP_3651 ();
 sky130_as_sc_hs__tap_1 TAP_3652 ();
 sky130_as_sc_hs__tap_1 TAP_3653 ();
 sky130_as_sc_hs__tap_1 TAP_3654 ();
 sky130_as_sc_hs__tap_1 TAP_3655 ();
 sky130_as_sc_hs__tap_1 TAP_3656 ();
 sky130_as_sc_hs__tap_1 TAP_3657 ();
 sky130_as_sc_hs__tap_1 TAP_3658 ();
 sky130_as_sc_hs__tap_1 TAP_3659 ();
 sky130_as_sc_hs__tap_1 TAP_3660 ();
 sky130_as_sc_hs__tap_1 TAP_3661 ();
 sky130_as_sc_hs__tap_1 TAP_3662 ();
 sky130_as_sc_hs__tap_1 TAP_3663 ();
 sky130_as_sc_hs__tap_1 TAP_3664 ();
 sky130_as_sc_hs__tap_1 TAP_3665 ();
 sky130_as_sc_hs__tap_1 TAP_3666 ();
 sky130_as_sc_hs__tap_1 TAP_3667 ();
 sky130_as_sc_hs__tap_1 TAP_3668 ();
 sky130_as_sc_hs__tap_1 TAP_3669 ();
 sky130_as_sc_hs__tap_1 TAP_3670 ();
 sky130_as_sc_hs__tap_1 TAP_3671 ();
 sky130_as_sc_hs__tap_1 TAP_3672 ();
 sky130_as_sc_hs__tap_1 TAP_3673 ();
 sky130_as_sc_hs__tap_1 TAP_3674 ();
 sky130_as_sc_hs__tap_1 TAP_3675 ();
 sky130_as_sc_hs__tap_1 TAP_3676 ();
 sky130_as_sc_hs__tap_1 TAP_3677 ();
 sky130_as_sc_hs__tap_1 TAP_3678 ();
 sky130_as_sc_hs__tap_1 TAP_3679 ();
 sky130_as_sc_hs__tap_1 TAP_3680 ();
 sky130_as_sc_hs__tap_1 TAP_3681 ();
 sky130_as_sc_hs__tap_1 TAP_3682 ();
 sky130_as_sc_hs__tap_1 TAP_3683 ();
 sky130_as_sc_hs__tap_1 TAP_3684 ();
 sky130_as_sc_hs__tap_1 TAP_3685 ();
 sky130_as_sc_hs__tap_1 TAP_3686 ();
 sky130_as_sc_hs__tap_1 TAP_3687 ();
 sky130_as_sc_hs__tap_1 TAP_3688 ();
 sky130_as_sc_hs__tap_1 TAP_3689 ();
 sky130_as_sc_hs__tap_1 TAP_3690 ();
 sky130_as_sc_hs__tap_1 TAP_3691 ();
 sky130_as_sc_hs__tap_1 TAP_3692 ();
 sky130_as_sc_hs__tap_1 TAP_3693 ();
 sky130_as_sc_hs__tap_1 TAP_3694 ();
 sky130_as_sc_hs__tap_1 TAP_3695 ();
 sky130_as_sc_hs__tap_1 TAP_3696 ();
 sky130_as_sc_hs__tap_1 TAP_3697 ();
 sky130_as_sc_hs__tap_1 TAP_3698 ();
 sky130_as_sc_hs__tap_1 TAP_3699 ();
 sky130_as_sc_hs__tap_1 TAP_3700 ();
 sky130_as_sc_hs__tap_1 TAP_3701 ();
 sky130_as_sc_hs__tap_1 TAP_3702 ();
 sky130_as_sc_hs__tap_1 TAP_3703 ();
 sky130_as_sc_hs__tap_1 TAP_3704 ();
 sky130_as_sc_hs__tap_1 TAP_3705 ();
 sky130_as_sc_hs__tap_1 TAP_3706 ();
 sky130_as_sc_hs__tap_1 TAP_3707 ();
 sky130_as_sc_hs__tap_1 TAP_3708 ();
 sky130_as_sc_hs__tap_1 TAP_3709 ();
 sky130_as_sc_hs__tap_1 TAP_3710 ();
 sky130_as_sc_hs__tap_1 TAP_3711 ();
 sky130_as_sc_hs__tap_1 TAP_3712 ();
 sky130_as_sc_hs__tap_1 TAP_3713 ();
 sky130_as_sc_hs__tap_1 TAP_3714 ();
 sky130_as_sc_hs__tap_1 TAP_3715 ();
 sky130_as_sc_hs__tap_1 TAP_3716 ();
 sky130_as_sc_hs__tap_1 TAP_3717 ();
 sky130_as_sc_hs__tap_1 TAP_3718 ();
 sky130_as_sc_hs__tap_1 TAP_3719 ();
 sky130_as_sc_hs__tap_1 TAP_3720 ();
 sky130_as_sc_hs__tap_1 TAP_3721 ();
 sky130_as_sc_hs__tap_1 TAP_3722 ();
 sky130_as_sc_hs__tap_1 TAP_3723 ();
 sky130_as_sc_hs__tap_1 TAP_3724 ();
 sky130_as_sc_hs__tap_1 TAP_3725 ();
 sky130_as_sc_hs__tap_1 TAP_3726 ();
 sky130_as_sc_hs__tap_1 TAP_3727 ();
 sky130_as_sc_hs__tap_1 TAP_3728 ();
 sky130_as_sc_hs__tap_1 TAP_3729 ();
 sky130_as_sc_hs__tap_1 TAP_3730 ();
 sky130_as_sc_hs__tap_1 TAP_3731 ();
 sky130_as_sc_hs__tap_1 TAP_3732 ();
 sky130_as_sc_hs__tap_1 TAP_3733 ();
 sky130_as_sc_hs__tap_1 TAP_3734 ();
 sky130_as_sc_hs__tap_1 TAP_3735 ();
 sky130_as_sc_hs__tap_1 TAP_3736 ();
 sky130_as_sc_hs__tap_1 TAP_3737 ();
 sky130_as_sc_hs__tap_1 TAP_3738 ();
 sky130_as_sc_hs__tap_1 TAP_3739 ();
 sky130_as_sc_hs__tap_1 TAP_3740 ();
 sky130_as_sc_hs__tap_1 TAP_3741 ();
 sky130_as_sc_hs__tap_1 TAP_3742 ();
 sky130_as_sc_hs__tap_1 TAP_3743 ();
 sky130_as_sc_hs__tap_1 TAP_3744 ();
 sky130_as_sc_hs__tap_1 TAP_3745 ();
 sky130_as_sc_hs__tap_1 TAP_3746 ();
 sky130_as_sc_hs__tap_1 TAP_3747 ();
 sky130_as_sc_hs__tap_1 TAP_3748 ();
 sky130_as_sc_hs__tap_1 TAP_3749 ();
 sky130_as_sc_hs__tap_1 TAP_3750 ();
 sky130_as_sc_hs__tap_1 TAP_3751 ();
 sky130_as_sc_hs__tap_1 TAP_3752 ();
 sky130_as_sc_hs__tap_1 TAP_3753 ();
 sky130_as_sc_hs__tap_1 TAP_3754 ();
 sky130_as_sc_hs__tap_1 TAP_3755 ();
 sky130_as_sc_hs__tap_1 TAP_3756 ();
 sky130_as_sc_hs__tap_1 TAP_3757 ();
 sky130_as_sc_hs__tap_1 TAP_3758 ();
 sky130_as_sc_hs__tap_1 TAP_3759 ();
 sky130_as_sc_hs__tap_1 TAP_3760 ();
 sky130_as_sc_hs__tap_1 TAP_3761 ();
 sky130_as_sc_hs__tap_1 TAP_3762 ();
 sky130_as_sc_hs__tap_1 TAP_3763 ();
 sky130_as_sc_hs__tap_1 TAP_3764 ();
 sky130_as_sc_hs__tap_1 TAP_3765 ();
 sky130_as_sc_hs__tap_1 TAP_3766 ();
 sky130_as_sc_hs__tap_1 TAP_3767 ();
 sky130_as_sc_hs__tap_1 TAP_3768 ();
 sky130_as_sc_hs__tap_1 TAP_3769 ();
 sky130_as_sc_hs__tap_1 TAP_3770 ();
 sky130_as_sc_hs__tap_1 TAP_3771 ();
 sky130_as_sc_hs__tap_1 TAP_3772 ();
 sky130_as_sc_hs__tap_1 TAP_3773 ();
 sky130_as_sc_hs__tap_1 TAP_3774 ();
 sky130_as_sc_hs__tap_1 TAP_3775 ();
 sky130_as_sc_hs__tap_1 TAP_3776 ();
 sky130_as_sc_hs__tap_1 TAP_3777 ();
 sky130_as_sc_hs__tap_1 TAP_3778 ();
 sky130_as_sc_hs__tap_1 TAP_3779 ();
 sky130_as_sc_hs__tap_1 TAP_3780 ();
 sky130_as_sc_hs__tap_1 TAP_3781 ();
 sky130_as_sc_hs__tap_1 TAP_3782 ();
 sky130_as_sc_hs__tap_1 TAP_3783 ();
 sky130_as_sc_hs__tap_1 TAP_3784 ();
 sky130_as_sc_hs__tap_1 TAP_3785 ();
 sky130_as_sc_hs__tap_1 TAP_3786 ();
 sky130_as_sc_hs__tap_1 TAP_3787 ();
 sky130_as_sc_hs__tap_1 TAP_3788 ();
 sky130_as_sc_hs__tap_1 TAP_3789 ();
 sky130_as_sc_hs__tap_1 TAP_3790 ();
 sky130_as_sc_hs__tap_1 TAP_3791 ();
 sky130_as_sc_hs__tap_1 TAP_3792 ();
 sky130_as_sc_hs__tap_1 TAP_3793 ();
 sky130_as_sc_hs__tap_1 TAP_3794 ();
 sky130_as_sc_hs__tap_1 TAP_3795 ();
 sky130_as_sc_hs__tap_1 TAP_3796 ();
 sky130_as_sc_hs__tap_1 TAP_3797 ();
 sky130_as_sc_hs__tap_1 TAP_3798 ();
 sky130_as_sc_hs__tap_1 TAP_3799 ();
 sky130_as_sc_hs__tap_1 TAP_3800 ();
 sky130_as_sc_hs__tap_1 TAP_3801 ();
 sky130_as_sc_hs__tap_1 TAP_3802 ();
 sky130_as_sc_hs__tap_1 TAP_3803 ();
 sky130_as_sc_hs__tap_1 TAP_3804 ();
 sky130_as_sc_hs__tap_1 TAP_3805 ();
 sky130_as_sc_hs__tap_1 TAP_3806 ();
 sky130_as_sc_hs__tap_1 TAP_3807 ();
 sky130_as_sc_hs__tap_1 TAP_3808 ();
 sky130_as_sc_hs__tap_1 TAP_3809 ();
 sky130_as_sc_hs__tap_1 TAP_3810 ();
 sky130_as_sc_hs__tap_1 TAP_3811 ();
 sky130_as_sc_hs__tap_1 TAP_3812 ();
 sky130_as_sc_hs__tap_1 TAP_3813 ();
 sky130_as_sc_hs__tap_1 TAP_3814 ();
 sky130_as_sc_hs__tap_1 TAP_3815 ();
 sky130_as_sc_hs__tap_1 TAP_3816 ();
 sky130_as_sc_hs__tap_1 TAP_3817 ();
 sky130_as_sc_hs__tap_1 TAP_3818 ();
 sky130_as_sc_hs__tap_1 TAP_3819 ();
 sky130_as_sc_hs__tap_1 TAP_3820 ();
 sky130_as_sc_hs__tap_1 TAP_3821 ();
 sky130_as_sc_hs__tap_1 TAP_3822 ();
 sky130_as_sc_hs__tap_1 TAP_3823 ();
 sky130_as_sc_hs__tap_1 TAP_3824 ();
 sky130_as_sc_hs__tap_1 TAP_3825 ();
 sky130_as_sc_hs__tap_1 TAP_3826 ();
 sky130_as_sc_hs__tap_1 TAP_3827 ();
 sky130_as_sc_hs__tap_1 TAP_3828 ();
 sky130_as_sc_hs__tap_1 TAP_3829 ();
 sky130_as_sc_hs__tap_1 TAP_3830 ();
 sky130_as_sc_hs__tap_1 TAP_3831 ();
 sky130_as_sc_hs__tap_1 TAP_3832 ();
 sky130_as_sc_hs__tap_1 TAP_3833 ();
 sky130_as_sc_hs__tap_1 TAP_3834 ();
 sky130_as_sc_hs__tap_1 TAP_3835 ();
 sky130_as_sc_hs__tap_1 TAP_3836 ();
 sky130_as_sc_hs__tap_1 TAP_3837 ();
 sky130_as_sc_hs__tap_1 TAP_3838 ();
 sky130_as_sc_hs__tap_1 TAP_3839 ();
 sky130_as_sc_hs__tap_1 TAP_3840 ();
 sky130_as_sc_hs__tap_1 TAP_3841 ();
 sky130_as_sc_hs__tap_1 TAP_3842 ();
 sky130_as_sc_hs__tap_1 TAP_3843 ();
 sky130_as_sc_hs__tap_1 TAP_3844 ();
 sky130_as_sc_hs__tap_1 TAP_3845 ();
 sky130_as_sc_hs__tap_1 TAP_3846 ();
 sky130_as_sc_hs__tap_1 TAP_3847 ();
 sky130_as_sc_hs__tap_1 TAP_3848 ();
 sky130_as_sc_hs__tap_1 TAP_3849 ();
 sky130_as_sc_hs__tap_1 TAP_3850 ();
 sky130_as_sc_hs__tap_1 TAP_3851 ();
 sky130_as_sc_hs__tap_1 TAP_3852 ();
 sky130_as_sc_hs__tap_1 TAP_3853 ();
 sky130_as_sc_hs__tap_1 TAP_3854 ();
 sky130_as_sc_hs__tap_1 TAP_3855 ();
 sky130_as_sc_hs__tap_1 TAP_3856 ();
 sky130_as_sc_hs__tap_1 TAP_3857 ();
 sky130_as_sc_hs__tap_1 TAP_3858 ();
 sky130_as_sc_hs__tap_1 TAP_3859 ();
 sky130_as_sc_hs__tap_1 TAP_3860 ();
 sky130_as_sc_hs__tap_1 TAP_3861 ();
 sky130_as_sc_hs__tap_1 TAP_3862 ();
 sky130_as_sc_hs__tap_1 TAP_3863 ();
 sky130_as_sc_hs__tap_1 TAP_3864 ();
 sky130_as_sc_hs__tap_1 TAP_3865 ();
 sky130_as_sc_hs__tap_1 TAP_3866 ();
 sky130_as_sc_hs__tap_1 TAP_3867 ();
 sky130_as_sc_hs__tap_1 TAP_3868 ();
 sky130_as_sc_hs__tap_1 TAP_3869 ();
 sky130_as_sc_hs__tap_1 TAP_3870 ();
 sky130_as_sc_hs__tap_1 TAP_3871 ();
 sky130_as_sc_hs__tap_1 TAP_3872 ();
 sky130_as_sc_hs__tap_1 TAP_3873 ();
 sky130_as_sc_hs__tap_1 TAP_3874 ();
 sky130_as_sc_hs__tap_1 TAP_3875 ();
 sky130_as_sc_hs__tap_1 TAP_3876 ();
 sky130_as_sc_hs__tap_1 TAP_3877 ();
 sky130_as_sc_hs__tap_1 TAP_3878 ();
 sky130_as_sc_hs__tap_1 TAP_3879 ();
 sky130_as_sc_hs__tap_1 TAP_3880 ();
 sky130_as_sc_hs__tap_1 TAP_3881 ();
 sky130_as_sc_hs__tap_1 TAP_3882 ();
 sky130_as_sc_hs__tap_1 TAP_3883 ();
 sky130_as_sc_hs__tap_1 TAP_3884 ();
 sky130_as_sc_hs__tap_1 TAP_3885 ();
 sky130_as_sc_hs__tap_1 TAP_3886 ();
 sky130_as_sc_hs__tap_1 TAP_3887 ();
 sky130_as_sc_hs__tap_1 TAP_3888 ();
 sky130_as_sc_hs__tap_1 TAP_3889 ();
 sky130_as_sc_hs__tap_1 TAP_3890 ();
 sky130_as_sc_hs__tap_1 TAP_3891 ();
 sky130_as_sc_hs__tap_1 TAP_3892 ();
 sky130_as_sc_hs__tap_1 TAP_3893 ();
 sky130_as_sc_hs__tap_1 TAP_3894 ();
 sky130_as_sc_hs__tap_1 TAP_3895 ();
 sky130_as_sc_hs__tap_1 TAP_3896 ();
 sky130_as_sc_hs__tap_1 TAP_3897 ();
 sky130_as_sc_hs__tap_1 TAP_3898 ();
 sky130_as_sc_hs__tap_1 TAP_3899 ();
 sky130_as_sc_hs__tap_1 TAP_3900 ();
 sky130_as_sc_hs__tap_1 TAP_3901 ();
 sky130_as_sc_hs__tap_1 TAP_3902 ();
 sky130_as_sc_hs__tap_1 TAP_3903 ();
 sky130_as_sc_hs__tap_1 TAP_3904 ();
 sky130_as_sc_hs__tap_1 TAP_3905 ();
 sky130_as_sc_hs__tap_1 TAP_3906 ();
 sky130_as_sc_hs__tap_1 TAP_3907 ();
 sky130_as_sc_hs__tap_1 TAP_3908 ();
 sky130_as_sc_hs__tap_1 TAP_3909 ();
 sky130_as_sc_hs__tap_1 TAP_3910 ();
 sky130_as_sc_hs__tap_1 TAP_3911 ();
 sky130_as_sc_hs__tap_1 TAP_3912 ();
 sky130_as_sc_hs__tap_1 TAP_3913 ();
 sky130_as_sc_hs__tap_1 TAP_3914 ();
 sky130_as_sc_hs__tap_1 TAP_3915 ();
 sky130_as_sc_hs__tap_1 TAP_3916 ();
 sky130_as_sc_hs__tap_1 TAP_3917 ();
 sky130_as_sc_hs__tap_1 TAP_3918 ();
 sky130_as_sc_hs__tap_1 TAP_3919 ();
 sky130_as_sc_hs__tap_1 TAP_3920 ();
 sky130_as_sc_hs__tap_1 TAP_3921 ();
 sky130_as_sc_hs__tap_1 TAP_3922 ();
 sky130_as_sc_hs__tap_1 TAP_3923 ();
 sky130_as_sc_hs__tap_1 TAP_3924 ();
 sky130_as_sc_hs__tap_1 TAP_3925 ();
 sky130_as_sc_hs__tap_1 TAP_3926 ();
 sky130_as_sc_hs__tap_1 TAP_3927 ();
 sky130_as_sc_hs__tap_1 TAP_3928 ();
 sky130_as_sc_hs__tap_1 TAP_3929 ();
 sky130_as_sc_hs__tap_1 TAP_3930 ();
 sky130_as_sc_hs__tap_1 TAP_3931 ();
 sky130_as_sc_hs__tap_1 TAP_3932 ();
 sky130_as_sc_hs__tap_1 TAP_3933 ();
 sky130_as_sc_hs__tap_1 TAP_3934 ();
 sky130_as_sc_hs__tap_1 TAP_3935 ();
 sky130_as_sc_hs__tap_1 TAP_3936 ();
 sky130_as_sc_hs__tap_1 TAP_3937 ();
 sky130_as_sc_hs__tap_1 TAP_3938 ();
 sky130_as_sc_hs__tap_1 TAP_3939 ();
 sky130_as_sc_hs__tap_1 TAP_3940 ();
 sky130_as_sc_hs__tap_1 TAP_3941 ();
 sky130_as_sc_hs__tap_1 TAP_3942 ();
 sky130_as_sc_hs__tap_1 TAP_3943 ();
 sky130_as_sc_hs__tap_1 TAP_3944 ();
 sky130_as_sc_hs__tap_1 TAP_3945 ();
 sky130_as_sc_hs__tap_1 TAP_3946 ();
 sky130_as_sc_hs__tap_1 TAP_3947 ();
 sky130_as_sc_hs__tap_1 TAP_3948 ();
 sky130_as_sc_hs__tap_1 TAP_3949 ();
 sky130_as_sc_hs__tap_1 TAP_3950 ();
 sky130_as_sc_hs__tap_1 TAP_3951 ();
 sky130_as_sc_hs__tap_1 TAP_3952 ();
 sky130_as_sc_hs__tap_1 TAP_3953 ();
 sky130_as_sc_hs__tap_1 TAP_3954 ();
 sky130_as_sc_hs__tap_1 TAP_3955 ();
 sky130_as_sc_hs__tap_1 TAP_3956 ();
 sky130_as_sc_hs__tap_1 TAP_3957 ();
 sky130_as_sc_hs__tap_1 TAP_3958 ();
 sky130_as_sc_hs__tap_1 TAP_3959 ();
 sky130_as_sc_hs__tap_1 TAP_3960 ();
 sky130_as_sc_hs__tap_1 TAP_3961 ();
 sky130_as_sc_hs__tap_1 TAP_3962 ();
 sky130_as_sc_hs__tap_1 TAP_3963 ();
 sky130_as_sc_hs__tap_1 TAP_3964 ();
 sky130_as_sc_hs__tap_1 TAP_3965 ();
 sky130_as_sc_hs__tap_1 TAP_3966 ();
 sky130_as_sc_hs__tap_1 TAP_3967 ();
 sky130_as_sc_hs__tap_1 TAP_3968 ();
 sky130_as_sc_hs__tap_1 TAP_3969 ();
 sky130_as_sc_hs__tap_1 TAP_3970 ();
 sky130_as_sc_hs__tap_1 TAP_3971 ();
 sky130_as_sc_hs__tap_1 TAP_3972 ();
 sky130_as_sc_hs__tap_1 TAP_3973 ();
 sky130_as_sc_hs__tap_1 TAP_3974 ();
 sky130_as_sc_hs__tap_1 TAP_3975 ();
 sky130_as_sc_hs__tap_1 TAP_3976 ();
 sky130_as_sc_hs__tap_1 TAP_3977 ();
 sky130_as_sc_hs__tap_1 TAP_3978 ();
 sky130_as_sc_hs__tap_1 TAP_3979 ();
 sky130_as_sc_hs__tap_1 TAP_3980 ();
 sky130_as_sc_hs__tap_1 TAP_3981 ();
 sky130_as_sc_hs__tap_1 TAP_3982 ();
 sky130_as_sc_hs__tap_1 TAP_3983 ();
 sky130_as_sc_hs__tap_1 TAP_3984 ();
 sky130_as_sc_hs__tap_1 TAP_3985 ();
 sky130_as_sc_hs__tap_1 TAP_3986 ();
 sky130_as_sc_hs__tap_1 TAP_3987 ();
 sky130_as_sc_hs__tap_1 TAP_3988 ();
 sky130_as_sc_hs__tap_1 TAP_3989 ();
 sky130_as_sc_hs__tap_1 TAP_3990 ();
 sky130_as_sc_hs__tap_1 TAP_3991 ();
 sky130_as_sc_hs__tap_1 TAP_3992 ();
 sky130_as_sc_hs__tap_1 TAP_3993 ();
 sky130_as_sc_hs__tap_1 TAP_3994 ();
 sky130_as_sc_hs__tap_1 TAP_3995 ();
 sky130_as_sc_hs__tap_1 TAP_3996 ();
 sky130_as_sc_hs__tap_1 TAP_3997 ();
 sky130_as_sc_hs__tap_1 TAP_3998 ();
 sky130_as_sc_hs__tap_1 TAP_3999 ();
 sky130_as_sc_hs__tap_1 TAP_4000 ();
 sky130_as_sc_hs__tap_1 TAP_4001 ();
 sky130_as_sc_hs__tap_1 TAP_4002 ();
 sky130_as_sc_hs__tap_1 TAP_4003 ();
 sky130_as_sc_hs__tap_1 TAP_4004 ();
 sky130_as_sc_hs__tap_1 TAP_4005 ();
 sky130_as_sc_hs__tap_1 TAP_4006 ();
 sky130_as_sc_hs__tap_1 TAP_4007 ();
 sky130_as_sc_hs__tap_1 TAP_4008 ();
 sky130_as_sc_hs__tap_1 TAP_4009 ();
 sky130_as_sc_hs__tap_1 TAP_4010 ();
 sky130_as_sc_hs__tap_1 TAP_4011 ();
 sky130_as_sc_hs__tap_1 TAP_4012 ();
 sky130_as_sc_hs__tap_1 TAP_4013 ();
 sky130_as_sc_hs__tap_1 TAP_4014 ();
 sky130_as_sc_hs__tap_1 TAP_4015 ();
 sky130_as_sc_hs__tap_1 TAP_4016 ();
 sky130_as_sc_hs__tap_1 TAP_4017 ();
 sky130_as_sc_hs__tap_1 TAP_4018 ();
 sky130_as_sc_hs__tap_1 TAP_4019 ();
 sky130_as_sc_hs__tap_1 TAP_4020 ();
 sky130_as_sc_hs__tap_1 TAP_4021 ();
 sky130_as_sc_hs__tap_1 TAP_4022 ();
 sky130_as_sc_hs__tap_1 TAP_4023 ();
 sky130_as_sc_hs__tap_1 TAP_4024 ();
 sky130_as_sc_hs__tap_1 TAP_4025 ();
 sky130_as_sc_hs__tap_1 TAP_4026 ();
 sky130_as_sc_hs__tap_1 TAP_4027 ();
 sky130_as_sc_hs__tap_1 TAP_4028 ();
 sky130_as_sc_hs__tap_1 TAP_4029 ();
 sky130_as_sc_hs__tap_1 TAP_4030 ();
 sky130_as_sc_hs__tap_1 TAP_4031 ();
 sky130_as_sc_hs__tap_1 TAP_4032 ();
 sky130_as_sc_hs__tap_1 TAP_4033 ();
 sky130_as_sc_hs__tap_1 TAP_4034 ();
 sky130_as_sc_hs__tap_1 TAP_4035 ();
 sky130_as_sc_hs__tap_1 TAP_4036 ();
 sky130_as_sc_hs__tap_1 TAP_4037 ();
 sky130_as_sc_hs__tap_1 TAP_4038 ();
 sky130_as_sc_hs__tap_1 TAP_4039 ();
 sky130_as_sc_hs__tap_1 TAP_4040 ();
 sky130_as_sc_hs__tap_1 TAP_4041 ();
 sky130_as_sc_hs__tap_1 TAP_4042 ();
 sky130_as_sc_hs__tap_1 TAP_4043 ();
 sky130_as_sc_hs__tap_1 TAP_4044 ();
 sky130_as_sc_hs__tap_1 TAP_4045 ();
 sky130_as_sc_hs__tap_1 TAP_4046 ();
 sky130_as_sc_hs__tap_1 TAP_4047 ();
 sky130_as_sc_hs__tap_1 TAP_4048 ();
 sky130_as_sc_hs__tap_1 TAP_4049 ();
 sky130_as_sc_hs__tap_1 TAP_4050 ();
 sky130_as_sc_hs__tap_1 TAP_4051 ();
 sky130_as_sc_hs__tap_1 TAP_4052 ();
 sky130_as_sc_hs__tap_1 TAP_4053 ();
 sky130_as_sc_hs__tap_1 TAP_4054 ();
 sky130_as_sc_hs__tap_1 TAP_4055 ();
 sky130_as_sc_hs__tap_1 TAP_4056 ();
 sky130_as_sc_hs__tap_1 TAP_4057 ();
 sky130_as_sc_hs__tap_1 TAP_4058 ();
 sky130_as_sc_hs__tap_1 TAP_4059 ();
 sky130_as_sc_hs__tap_1 TAP_4060 ();
 sky130_as_sc_hs__tap_1 TAP_4061 ();
 sky130_as_sc_hs__tap_1 TAP_4062 ();
 sky130_as_sc_hs__tap_1 TAP_4063 ();
 sky130_as_sc_hs__tap_1 TAP_4064 ();
 sky130_as_sc_hs__tap_1 TAP_4065 ();
 sky130_as_sc_hs__tap_1 TAP_4066 ();
 sky130_as_sc_hs__tap_1 TAP_4067 ();
 sky130_as_sc_hs__tap_1 TAP_4068 ();
 sky130_as_sc_hs__tap_1 TAP_4069 ();
 sky130_as_sc_hs__tap_1 TAP_4070 ();
 sky130_as_sc_hs__tap_1 TAP_4071 ();
 sky130_as_sc_hs__tap_1 TAP_4072 ();
 sky130_as_sc_hs__tap_1 TAP_4073 ();
 sky130_as_sc_hs__tap_1 TAP_4074 ();
 sky130_as_sc_hs__tap_1 TAP_4075 ();
 sky130_as_sc_hs__tap_1 TAP_4076 ();
 sky130_as_sc_hs__tap_1 TAP_4077 ();
 sky130_as_sc_hs__tap_1 TAP_4078 ();
 sky130_as_sc_hs__tap_1 TAP_4079 ();
 sky130_as_sc_hs__tap_1 TAP_4080 ();
 sky130_as_sc_hs__tap_1 TAP_4081 ();
 sky130_as_sc_hs__tap_1 TAP_4082 ();
 sky130_as_sc_hs__tap_1 TAP_4083 ();
 sky130_as_sc_hs__tap_1 TAP_4084 ();
 sky130_as_sc_hs__tap_1 TAP_4085 ();
 sky130_as_sc_hs__tap_1 TAP_4086 ();
 sky130_as_sc_hs__tap_1 TAP_4087 ();
 sky130_as_sc_hs__tap_1 TAP_4088 ();
 sky130_as_sc_hs__tap_1 TAP_4089 ();
 sky130_as_sc_hs__tap_1 TAP_4090 ();
 sky130_as_sc_hs__tap_1 TAP_4091 ();
 sky130_as_sc_hs__tap_1 TAP_4092 ();
 sky130_as_sc_hs__tap_1 TAP_4093 ();
 sky130_as_sc_hs__tap_1 TAP_4094 ();
 sky130_as_sc_hs__tap_1 TAP_4095 ();
 sky130_as_sc_hs__tap_1 TAP_4096 ();
 sky130_as_sc_hs__tap_1 TAP_4097 ();
 sky130_as_sc_hs__tap_1 TAP_4098 ();
 sky130_as_sc_hs__tap_1 TAP_4099 ();
 sky130_as_sc_hs__tap_1 TAP_4100 ();
 sky130_as_sc_hs__tap_1 TAP_4101 ();
 sky130_as_sc_hs__tap_1 TAP_4102 ();
 sky130_as_sc_hs__tap_1 TAP_4103 ();
 sky130_as_sc_hs__tap_1 TAP_4104 ();
 sky130_as_sc_hs__tap_1 TAP_4105 ();
 sky130_as_sc_hs__tap_1 TAP_4106 ();
 sky130_as_sc_hs__tap_1 TAP_4107 ();
 sky130_as_sc_hs__tap_1 TAP_4108 ();
 sky130_as_sc_hs__tap_1 TAP_4109 ();
 sky130_as_sc_hs__tap_1 TAP_4110 ();
 sky130_as_sc_hs__tap_1 TAP_4111 ();
 sky130_as_sc_hs__tap_1 TAP_4112 ();
 sky130_as_sc_hs__tap_1 TAP_4113 ();
 sky130_as_sc_hs__tap_1 TAP_4114 ();
 sky130_as_sc_hs__tap_1 TAP_4115 ();
 sky130_as_sc_hs__tap_1 TAP_4116 ();
 sky130_as_sc_hs__tap_1 TAP_4117 ();
 sky130_as_sc_hs__tap_1 TAP_4118 ();
 sky130_as_sc_hs__tap_1 TAP_4119 ();
 sky130_as_sc_hs__tap_1 TAP_4120 ();
 sky130_as_sc_hs__tap_1 TAP_4121 ();
 sky130_as_sc_hs__tap_1 TAP_4122 ();
 sky130_as_sc_hs__tap_1 TAP_4123 ();
 sky130_as_sc_hs__tap_1 TAP_4124 ();
 sky130_as_sc_hs__tap_1 TAP_4125 ();
 sky130_as_sc_hs__tap_1 TAP_4126 ();
 sky130_as_sc_hs__tap_1 TAP_4127 ();
 sky130_as_sc_hs__tap_1 TAP_4128 ();
 sky130_as_sc_hs__tap_1 TAP_4129 ();
 sky130_as_sc_hs__tap_1 TAP_4130 ();
 sky130_as_sc_hs__tap_1 TAP_4131 ();
 sky130_as_sc_hs__tap_1 TAP_4132 ();
 sky130_as_sc_hs__tap_1 TAP_4133 ();
 sky130_as_sc_hs__tap_1 TAP_4134 ();
 sky130_as_sc_hs__tap_1 TAP_4135 ();
 sky130_as_sc_hs__tap_1 TAP_4136 ();
 sky130_as_sc_hs__tap_1 TAP_4137 ();
 sky130_as_sc_hs__tap_1 TAP_4138 ();
 sky130_as_sc_hs__tap_1 TAP_4139 ();
 sky130_as_sc_hs__tap_1 TAP_4140 ();
 sky130_as_sc_hs__tap_1 TAP_4141 ();
 sky130_as_sc_hs__tap_1 TAP_4142 ();
 sky130_as_sc_hs__tap_1 TAP_4143 ();
 sky130_as_sc_hs__tap_1 TAP_4144 ();
 sky130_as_sc_hs__tap_1 TAP_4145 ();
 sky130_as_sc_hs__tap_1 TAP_4146 ();
 sky130_as_sc_hs__tap_1 TAP_4147 ();
 sky130_as_sc_hs__tap_1 TAP_4148 ();
 sky130_as_sc_hs__tap_1 TAP_4149 ();
 sky130_as_sc_hs__tap_1 TAP_4150 ();
 sky130_as_sc_hs__tap_1 TAP_4151 ();
 sky130_as_sc_hs__tap_1 TAP_4152 ();
 sky130_as_sc_hs__tap_1 TAP_4153 ();
 sky130_as_sc_hs__tap_1 TAP_4154 ();
 sky130_as_sc_hs__tap_1 TAP_4155 ();
 sky130_as_sc_hs__tap_1 TAP_4156 ();
 sky130_as_sc_hs__tap_1 TAP_4157 ();
 sky130_as_sc_hs__tap_1 TAP_4158 ();
 sky130_as_sc_hs__tap_1 TAP_4159 ();
 sky130_as_sc_hs__tap_1 TAP_4160 ();
 sky130_as_sc_hs__tap_1 TAP_4161 ();
 sky130_as_sc_hs__tap_1 TAP_4162 ();
 sky130_as_sc_hs__tap_1 TAP_4163 ();
 sky130_as_sc_hs__tap_1 TAP_4164 ();
 sky130_as_sc_hs__tap_1 TAP_4165 ();
 sky130_as_sc_hs__tap_1 TAP_4166 ();
 sky130_as_sc_hs__tap_1 TAP_4167 ();
 sky130_as_sc_hs__tap_1 TAP_4168 ();
 sky130_as_sc_hs__tap_1 TAP_4169 ();
 sky130_as_sc_hs__tap_1 TAP_4170 ();
 sky130_as_sc_hs__tap_1 TAP_4171 ();
 sky130_as_sc_hs__tap_1 TAP_4172 ();
 sky130_as_sc_hs__tap_1 TAP_4173 ();
 sky130_as_sc_hs__tap_1 TAP_4174 ();
 sky130_as_sc_hs__tap_1 TAP_4175 ();
 sky130_as_sc_hs__tap_1 TAP_4176 ();
 sky130_as_sc_hs__tap_1 TAP_4177 ();
 sky130_as_sc_hs__tap_1 TAP_4178 ();
 sky130_as_sc_hs__tap_1 TAP_4179 ();
 sky130_as_sc_hs__tap_1 TAP_4180 ();
 sky130_as_sc_hs__tap_1 TAP_4181 ();
 sky130_as_sc_hs__tap_1 TAP_4182 ();
 sky130_as_sc_hs__tap_1 TAP_4183 ();
 sky130_as_sc_hs__tap_1 TAP_4184 ();
 sky130_as_sc_hs__tap_1 TAP_4185 ();
 sky130_as_sc_hs__tap_1 TAP_4186 ();
 sky130_as_sc_hs__tap_1 TAP_4187 ();
 sky130_as_sc_hs__tap_1 TAP_4188 ();
 sky130_as_sc_hs__tap_1 TAP_4189 ();
 sky130_as_sc_hs__tap_1 TAP_4190 ();
 sky130_as_sc_hs__tap_1 TAP_4191 ();
 sky130_as_sc_hs__tap_1 TAP_4192 ();
 sky130_as_sc_hs__tap_1 TAP_4193 ();
 sky130_as_sc_hs__tap_1 TAP_4194 ();
 sky130_as_sc_hs__tap_1 TAP_4195 ();
 sky130_as_sc_hs__tap_1 TAP_4196 ();
 sky130_as_sc_hs__tap_1 TAP_4197 ();
 sky130_as_sc_hs__tap_1 TAP_4198 ();
 sky130_as_sc_hs__tap_1 TAP_4199 ();
 sky130_as_sc_hs__tap_1 TAP_4200 ();
 sky130_as_sc_hs__tap_1 TAP_4201 ();
 sky130_as_sc_hs__tap_1 TAP_4202 ();
 sky130_as_sc_hs__tap_1 TAP_4203 ();
 sky130_as_sc_hs__tap_1 TAP_4204 ();
 sky130_as_sc_hs__tap_1 TAP_4205 ();
 sky130_as_sc_hs__tap_1 TAP_4206 ();
 sky130_as_sc_hs__tap_1 TAP_4207 ();
 sky130_as_sc_hs__tap_1 TAP_4208 ();
 sky130_as_sc_hs__tap_1 TAP_4209 ();
 sky130_as_sc_hs__tap_1 TAP_4210 ();
 sky130_as_sc_hs__tap_1 TAP_4211 ();
 sky130_as_sc_hs__tap_1 TAP_4212 ();
 sky130_as_sc_hs__tap_1 TAP_4213 ();
 sky130_as_sc_hs__tap_1 TAP_4214 ();
 sky130_as_sc_hs__tap_1 TAP_4215 ();
 sky130_as_sc_hs__tap_1 TAP_4216 ();
 sky130_as_sc_hs__tap_1 TAP_4217 ();
 sky130_as_sc_hs__tap_1 TAP_4218 ();
 sky130_as_sc_hs__tap_1 TAP_4219 ();
 sky130_as_sc_hs__tap_1 TAP_4220 ();
 sky130_as_sc_hs__tap_1 TAP_4221 ();
 sky130_as_sc_hs__tap_1 TAP_4222 ();
 sky130_as_sc_hs__tap_1 TAP_4223 ();
 sky130_as_sc_hs__tap_1 TAP_4224 ();
 sky130_as_sc_hs__tap_1 TAP_4225 ();
 sky130_as_sc_hs__tap_1 TAP_4226 ();
 sky130_as_sc_hs__tap_1 TAP_4227 ();
 sky130_as_sc_hs__tap_1 TAP_4228 ();
 sky130_as_sc_hs__tap_1 TAP_4229 ();
 sky130_as_sc_hs__tap_1 TAP_4230 ();
 sky130_as_sc_hs__tap_1 TAP_4231 ();
 sky130_as_sc_hs__tap_1 TAP_4232 ();
 sky130_as_sc_hs__tap_1 TAP_4233 ();
 sky130_as_sc_hs__tap_1 TAP_4234 ();
 sky130_as_sc_hs__tap_1 TAP_4235 ();
 sky130_as_sc_hs__tap_1 TAP_4236 ();
 sky130_as_sc_hs__tap_1 TAP_4237 ();
 sky130_as_sc_hs__tap_1 TAP_4238 ();
 sky130_as_sc_hs__tap_1 TAP_4239 ();
 sky130_as_sc_hs__tap_1 TAP_424 ();
 sky130_as_sc_hs__tap_1 TAP_4240 ();
 sky130_as_sc_hs__tap_1 TAP_4241 ();
 sky130_as_sc_hs__tap_1 TAP_4242 ();
 sky130_as_sc_hs__tap_1 TAP_4243 ();
 sky130_as_sc_hs__tap_1 TAP_4244 ();
 sky130_as_sc_hs__tap_1 TAP_4245 ();
 sky130_as_sc_hs__tap_1 TAP_4246 ();
 sky130_as_sc_hs__tap_1 TAP_4247 ();
 sky130_as_sc_hs__tap_1 TAP_4248 ();
 sky130_as_sc_hs__tap_1 TAP_4249 ();
 sky130_as_sc_hs__tap_1 TAP_425 ();
 sky130_as_sc_hs__tap_1 TAP_4250 ();
 sky130_as_sc_hs__tap_1 TAP_4251 ();
 sky130_as_sc_hs__tap_1 TAP_4252 ();
 sky130_as_sc_hs__tap_1 TAP_4253 ();
 sky130_as_sc_hs__tap_1 TAP_4254 ();
 sky130_as_sc_hs__tap_1 TAP_4255 ();
 sky130_as_sc_hs__tap_1 TAP_4256 ();
 sky130_as_sc_hs__tap_1 TAP_4257 ();
 sky130_as_sc_hs__tap_1 TAP_4258 ();
 sky130_as_sc_hs__tap_1 TAP_4259 ();
 sky130_as_sc_hs__tap_1 TAP_426 ();
 sky130_as_sc_hs__tap_1 TAP_4260 ();
 sky130_as_sc_hs__tap_1 TAP_4261 ();
 sky130_as_sc_hs__tap_1 TAP_4262 ();
 sky130_as_sc_hs__tap_1 TAP_4263 ();
 sky130_as_sc_hs__tap_1 TAP_4264 ();
 sky130_as_sc_hs__tap_1 TAP_4265 ();
 sky130_as_sc_hs__tap_1 TAP_4266 ();
 sky130_as_sc_hs__tap_1 TAP_4267 ();
 sky130_as_sc_hs__tap_1 TAP_4268 ();
 sky130_as_sc_hs__tap_1 TAP_4269 ();
 sky130_as_sc_hs__tap_1 TAP_427 ();
 sky130_as_sc_hs__tap_1 TAP_4270 ();
 sky130_as_sc_hs__tap_1 TAP_4271 ();
 sky130_as_sc_hs__tap_1 TAP_4272 ();
 sky130_as_sc_hs__tap_1 TAP_4273 ();
 sky130_as_sc_hs__tap_1 TAP_4274 ();
 sky130_as_sc_hs__tap_1 TAP_4275 ();
 sky130_as_sc_hs__tap_1 TAP_4276 ();
 sky130_as_sc_hs__tap_1 TAP_4277 ();
 sky130_as_sc_hs__tap_1 TAP_4278 ();
 sky130_as_sc_hs__tap_1 TAP_4279 ();
 sky130_as_sc_hs__tap_1 TAP_428 ();
 sky130_as_sc_hs__tap_1 TAP_4280 ();
 sky130_as_sc_hs__tap_1 TAP_4281 ();
 sky130_as_sc_hs__tap_1 TAP_4282 ();
 sky130_as_sc_hs__tap_1 TAP_4283 ();
 sky130_as_sc_hs__tap_1 TAP_4284 ();
 sky130_as_sc_hs__tap_1 TAP_4285 ();
 sky130_as_sc_hs__tap_1 TAP_4286 ();
 sky130_as_sc_hs__tap_1 TAP_4287 ();
 sky130_as_sc_hs__tap_1 TAP_4288 ();
 sky130_as_sc_hs__tap_1 TAP_4289 ();
 sky130_as_sc_hs__tap_1 TAP_429 ();
 sky130_as_sc_hs__tap_1 TAP_4290 ();
 sky130_as_sc_hs__tap_1 TAP_4291 ();
 sky130_as_sc_hs__tap_1 TAP_4292 ();
 sky130_as_sc_hs__tap_1 TAP_4293 ();
 sky130_as_sc_hs__tap_1 TAP_4294 ();
 sky130_as_sc_hs__tap_1 TAP_4295 ();
 sky130_as_sc_hs__tap_1 TAP_4296 ();
 sky130_as_sc_hs__tap_1 TAP_4297 ();
 sky130_as_sc_hs__tap_1 TAP_4298 ();
 sky130_as_sc_hs__tap_1 TAP_4299 ();
 sky130_as_sc_hs__tap_1 TAP_430 ();
 sky130_as_sc_hs__tap_1 TAP_4300 ();
 sky130_as_sc_hs__tap_1 TAP_4301 ();
 sky130_as_sc_hs__tap_1 TAP_4302 ();
 sky130_as_sc_hs__tap_1 TAP_4303 ();
 sky130_as_sc_hs__tap_1 TAP_4304 ();
 sky130_as_sc_hs__tap_1 TAP_4305 ();
 sky130_as_sc_hs__tap_1 TAP_4306 ();
 sky130_as_sc_hs__tap_1 TAP_4307 ();
 sky130_as_sc_hs__tap_1 TAP_4308 ();
 sky130_as_sc_hs__tap_1 TAP_4309 ();
 sky130_as_sc_hs__tap_1 TAP_431 ();
 sky130_as_sc_hs__tap_1 TAP_4310 ();
 sky130_as_sc_hs__tap_1 TAP_4311 ();
 sky130_as_sc_hs__tap_1 TAP_4312 ();
 sky130_as_sc_hs__tap_1 TAP_4313 ();
 sky130_as_sc_hs__tap_1 TAP_4314 ();
 sky130_as_sc_hs__tap_1 TAP_4315 ();
 sky130_as_sc_hs__tap_1 TAP_4316 ();
 sky130_as_sc_hs__tap_1 TAP_4317 ();
 sky130_as_sc_hs__tap_1 TAP_4318 ();
 sky130_as_sc_hs__tap_1 TAP_4319 ();
 sky130_as_sc_hs__tap_1 TAP_432 ();
 sky130_as_sc_hs__tap_1 TAP_4320 ();
 sky130_as_sc_hs__tap_1 TAP_4321 ();
 sky130_as_sc_hs__tap_1 TAP_4322 ();
 sky130_as_sc_hs__tap_1 TAP_4323 ();
 sky130_as_sc_hs__tap_1 TAP_4324 ();
 sky130_as_sc_hs__tap_1 TAP_4325 ();
 sky130_as_sc_hs__tap_1 TAP_4326 ();
 sky130_as_sc_hs__tap_1 TAP_4327 ();
 sky130_as_sc_hs__tap_1 TAP_4328 ();
 sky130_as_sc_hs__tap_1 TAP_4329 ();
 sky130_as_sc_hs__tap_1 TAP_433 ();
 sky130_as_sc_hs__tap_1 TAP_4330 ();
 sky130_as_sc_hs__tap_1 TAP_4331 ();
 sky130_as_sc_hs__tap_1 TAP_4332 ();
 sky130_as_sc_hs__tap_1 TAP_4333 ();
 sky130_as_sc_hs__tap_1 TAP_4334 ();
 sky130_as_sc_hs__tap_1 TAP_4335 ();
 sky130_as_sc_hs__tap_1 TAP_4336 ();
 sky130_as_sc_hs__tap_1 TAP_4337 ();
 sky130_as_sc_hs__tap_1 TAP_4338 ();
 sky130_as_sc_hs__tap_1 TAP_4339 ();
 sky130_as_sc_hs__tap_1 TAP_434 ();
 sky130_as_sc_hs__tap_1 TAP_4340 ();
 sky130_as_sc_hs__tap_1 TAP_4341 ();
 sky130_as_sc_hs__tap_1 TAP_4342 ();
 sky130_as_sc_hs__tap_1 TAP_4343 ();
 sky130_as_sc_hs__tap_1 TAP_4344 ();
 sky130_as_sc_hs__tap_1 TAP_4345 ();
 sky130_as_sc_hs__tap_1 TAP_4346 ();
 sky130_as_sc_hs__tap_1 TAP_4347 ();
 sky130_as_sc_hs__tap_1 TAP_4348 ();
 sky130_as_sc_hs__tap_1 TAP_4349 ();
 sky130_as_sc_hs__tap_1 TAP_435 ();
 sky130_as_sc_hs__tap_1 TAP_4350 ();
 sky130_as_sc_hs__tap_1 TAP_4351 ();
 sky130_as_sc_hs__tap_1 TAP_4352 ();
 sky130_as_sc_hs__tap_1 TAP_4353 ();
 sky130_as_sc_hs__tap_1 TAP_4354 ();
 sky130_as_sc_hs__tap_1 TAP_4355 ();
 sky130_as_sc_hs__tap_1 TAP_4356 ();
 sky130_as_sc_hs__tap_1 TAP_4357 ();
 sky130_as_sc_hs__tap_1 TAP_4358 ();
 sky130_as_sc_hs__tap_1 TAP_4359 ();
 sky130_as_sc_hs__tap_1 TAP_436 ();
 sky130_as_sc_hs__tap_1 TAP_4360 ();
 sky130_as_sc_hs__tap_1 TAP_4361 ();
 sky130_as_sc_hs__tap_1 TAP_4362 ();
 sky130_as_sc_hs__tap_1 TAP_4363 ();
 sky130_as_sc_hs__tap_1 TAP_4364 ();
 sky130_as_sc_hs__tap_1 TAP_4365 ();
 sky130_as_sc_hs__tap_1 TAP_4366 ();
 sky130_as_sc_hs__tap_1 TAP_4367 ();
 sky130_as_sc_hs__tap_1 TAP_4368 ();
 sky130_as_sc_hs__tap_1 TAP_4369 ();
 sky130_as_sc_hs__tap_1 TAP_437 ();
 sky130_as_sc_hs__tap_1 TAP_4370 ();
 sky130_as_sc_hs__tap_1 TAP_4371 ();
 sky130_as_sc_hs__tap_1 TAP_4372 ();
 sky130_as_sc_hs__tap_1 TAP_4373 ();
 sky130_as_sc_hs__tap_1 TAP_4374 ();
 sky130_as_sc_hs__tap_1 TAP_4375 ();
 sky130_as_sc_hs__tap_1 TAP_4376 ();
 sky130_as_sc_hs__tap_1 TAP_4377 ();
 sky130_as_sc_hs__tap_1 TAP_4378 ();
 sky130_as_sc_hs__tap_1 TAP_4379 ();
 sky130_as_sc_hs__tap_1 TAP_438 ();
 sky130_as_sc_hs__tap_1 TAP_4380 ();
 sky130_as_sc_hs__tap_1 TAP_4381 ();
 sky130_as_sc_hs__tap_1 TAP_4382 ();
 sky130_as_sc_hs__tap_1 TAP_4383 ();
 sky130_as_sc_hs__tap_1 TAP_4384 ();
 sky130_as_sc_hs__tap_1 TAP_4385 ();
 sky130_as_sc_hs__tap_1 TAP_4386 ();
 sky130_as_sc_hs__tap_1 TAP_4387 ();
 sky130_as_sc_hs__tap_1 TAP_4388 ();
 sky130_as_sc_hs__tap_1 TAP_4389 ();
 sky130_as_sc_hs__tap_1 TAP_439 ();
 sky130_as_sc_hs__tap_1 TAP_4390 ();
 sky130_as_sc_hs__tap_1 TAP_4391 ();
 sky130_as_sc_hs__tap_1 TAP_4392 ();
 sky130_as_sc_hs__tap_1 TAP_4393 ();
 sky130_as_sc_hs__tap_1 TAP_4394 ();
 sky130_as_sc_hs__tap_1 TAP_4395 ();
 sky130_as_sc_hs__tap_1 TAP_4396 ();
 sky130_as_sc_hs__tap_1 TAP_4397 ();
 sky130_as_sc_hs__tap_1 TAP_4398 ();
 sky130_as_sc_hs__tap_1 TAP_4399 ();
 sky130_as_sc_hs__tap_1 TAP_440 ();
 sky130_as_sc_hs__tap_1 TAP_4400 ();
 sky130_as_sc_hs__tap_1 TAP_4401 ();
 sky130_as_sc_hs__tap_1 TAP_4402 ();
 sky130_as_sc_hs__tap_1 TAP_4403 ();
 sky130_as_sc_hs__tap_1 TAP_4404 ();
 sky130_as_sc_hs__tap_1 TAP_4405 ();
 sky130_as_sc_hs__tap_1 TAP_4406 ();
 sky130_as_sc_hs__tap_1 TAP_4407 ();
 sky130_as_sc_hs__tap_1 TAP_4408 ();
 sky130_as_sc_hs__tap_1 TAP_4409 ();
 sky130_as_sc_hs__tap_1 TAP_441 ();
 sky130_as_sc_hs__tap_1 TAP_4410 ();
 sky130_as_sc_hs__tap_1 TAP_4411 ();
 sky130_as_sc_hs__tap_1 TAP_4412 ();
 sky130_as_sc_hs__tap_1 TAP_4413 ();
 sky130_as_sc_hs__tap_1 TAP_4414 ();
 sky130_as_sc_hs__tap_1 TAP_4415 ();
 sky130_as_sc_hs__tap_1 TAP_4416 ();
 sky130_as_sc_hs__tap_1 TAP_4417 ();
 sky130_as_sc_hs__tap_1 TAP_4418 ();
 sky130_as_sc_hs__tap_1 TAP_4419 ();
 sky130_as_sc_hs__tap_1 TAP_442 ();
 sky130_as_sc_hs__tap_1 TAP_4420 ();
 sky130_as_sc_hs__tap_1 TAP_4421 ();
 sky130_as_sc_hs__tap_1 TAP_4422 ();
 sky130_as_sc_hs__tap_1 TAP_4423 ();
 sky130_as_sc_hs__tap_1 TAP_4424 ();
 sky130_as_sc_hs__tap_1 TAP_4425 ();
 sky130_as_sc_hs__tap_1 TAP_4426 ();
 sky130_as_sc_hs__tap_1 TAP_4427 ();
 sky130_as_sc_hs__tap_1 TAP_4428 ();
 sky130_as_sc_hs__tap_1 TAP_4429 ();
 sky130_as_sc_hs__tap_1 TAP_443 ();
 sky130_as_sc_hs__tap_1 TAP_4430 ();
 sky130_as_sc_hs__tap_1 TAP_4431 ();
 sky130_as_sc_hs__tap_1 TAP_4432 ();
 sky130_as_sc_hs__tap_1 TAP_4433 ();
 sky130_as_sc_hs__tap_1 TAP_4434 ();
 sky130_as_sc_hs__tap_1 TAP_4435 ();
 sky130_as_sc_hs__tap_1 TAP_4436 ();
 sky130_as_sc_hs__tap_1 TAP_4437 ();
 sky130_as_sc_hs__tap_1 TAP_4438 ();
 sky130_as_sc_hs__tap_1 TAP_4439 ();
 sky130_as_sc_hs__tap_1 TAP_444 ();
 sky130_as_sc_hs__tap_1 TAP_4440 ();
 sky130_as_sc_hs__tap_1 TAP_4441 ();
 sky130_as_sc_hs__tap_1 TAP_4442 ();
 sky130_as_sc_hs__tap_1 TAP_4443 ();
 sky130_as_sc_hs__tap_1 TAP_4444 ();
 sky130_as_sc_hs__tap_1 TAP_4445 ();
 sky130_as_sc_hs__tap_1 TAP_4446 ();
 sky130_as_sc_hs__tap_1 TAP_4447 ();
 sky130_as_sc_hs__tap_1 TAP_4448 ();
 sky130_as_sc_hs__tap_1 TAP_4449 ();
 sky130_as_sc_hs__tap_1 TAP_445 ();
 sky130_as_sc_hs__tap_1 TAP_4450 ();
 sky130_as_sc_hs__tap_1 TAP_4451 ();
 sky130_as_sc_hs__tap_1 TAP_4452 ();
 sky130_as_sc_hs__tap_1 TAP_4453 ();
 sky130_as_sc_hs__tap_1 TAP_4454 ();
 sky130_as_sc_hs__tap_1 TAP_4455 ();
 sky130_as_sc_hs__tap_1 TAP_4456 ();
 sky130_as_sc_hs__tap_1 TAP_4457 ();
 sky130_as_sc_hs__tap_1 TAP_4458 ();
 sky130_as_sc_hs__tap_1 TAP_4459 ();
 sky130_as_sc_hs__tap_1 TAP_446 ();
 sky130_as_sc_hs__tap_1 TAP_4460 ();
 sky130_as_sc_hs__tap_1 TAP_4461 ();
 sky130_as_sc_hs__tap_1 TAP_4462 ();
 sky130_as_sc_hs__tap_1 TAP_4463 ();
 sky130_as_sc_hs__tap_1 TAP_4464 ();
 sky130_as_sc_hs__tap_1 TAP_4465 ();
 sky130_as_sc_hs__tap_1 TAP_4466 ();
 sky130_as_sc_hs__tap_1 TAP_4467 ();
 sky130_as_sc_hs__tap_1 TAP_4468 ();
 sky130_as_sc_hs__tap_1 TAP_4469 ();
 sky130_as_sc_hs__tap_1 TAP_447 ();
 sky130_as_sc_hs__tap_1 TAP_4470 ();
 sky130_as_sc_hs__tap_1 TAP_4471 ();
 sky130_as_sc_hs__tap_1 TAP_4472 ();
 sky130_as_sc_hs__tap_1 TAP_4473 ();
 sky130_as_sc_hs__tap_1 TAP_4474 ();
 sky130_as_sc_hs__tap_1 TAP_4475 ();
 sky130_as_sc_hs__tap_1 TAP_4476 ();
 sky130_as_sc_hs__tap_1 TAP_4477 ();
 sky130_as_sc_hs__tap_1 TAP_4478 ();
 sky130_as_sc_hs__tap_1 TAP_4479 ();
 sky130_as_sc_hs__tap_1 TAP_448 ();
 sky130_as_sc_hs__tap_1 TAP_4480 ();
 sky130_as_sc_hs__tap_1 TAP_4481 ();
 sky130_as_sc_hs__tap_1 TAP_4482 ();
 sky130_as_sc_hs__tap_1 TAP_4483 ();
 sky130_as_sc_hs__tap_1 TAP_4484 ();
 sky130_as_sc_hs__tap_1 TAP_4485 ();
 sky130_as_sc_hs__tap_1 TAP_4486 ();
 sky130_as_sc_hs__tap_1 TAP_4487 ();
 sky130_as_sc_hs__tap_1 TAP_4488 ();
 sky130_as_sc_hs__tap_1 TAP_4489 ();
 sky130_as_sc_hs__tap_1 TAP_449 ();
 sky130_as_sc_hs__tap_1 TAP_4490 ();
 sky130_as_sc_hs__tap_1 TAP_4491 ();
 sky130_as_sc_hs__tap_1 TAP_4492 ();
 sky130_as_sc_hs__tap_1 TAP_4493 ();
 sky130_as_sc_hs__tap_1 TAP_4494 ();
 sky130_as_sc_hs__tap_1 TAP_4495 ();
 sky130_as_sc_hs__tap_1 TAP_4496 ();
 sky130_as_sc_hs__tap_1 TAP_4497 ();
 sky130_as_sc_hs__tap_1 TAP_4498 ();
 sky130_as_sc_hs__tap_1 TAP_4499 ();
 sky130_as_sc_hs__tap_1 TAP_450 ();
 sky130_as_sc_hs__tap_1 TAP_4500 ();
 sky130_as_sc_hs__tap_1 TAP_4501 ();
 sky130_as_sc_hs__tap_1 TAP_4502 ();
 sky130_as_sc_hs__tap_1 TAP_4503 ();
 sky130_as_sc_hs__tap_1 TAP_4504 ();
 sky130_as_sc_hs__tap_1 TAP_4505 ();
 sky130_as_sc_hs__tap_1 TAP_4506 ();
 sky130_as_sc_hs__tap_1 TAP_4507 ();
 sky130_as_sc_hs__tap_1 TAP_4508 ();
 sky130_as_sc_hs__tap_1 TAP_4509 ();
 sky130_as_sc_hs__tap_1 TAP_451 ();
 sky130_as_sc_hs__tap_1 TAP_4510 ();
 sky130_as_sc_hs__tap_1 TAP_4511 ();
 sky130_as_sc_hs__tap_1 TAP_4512 ();
 sky130_as_sc_hs__tap_1 TAP_4513 ();
 sky130_as_sc_hs__tap_1 TAP_4514 ();
 sky130_as_sc_hs__tap_1 TAP_4515 ();
 sky130_as_sc_hs__tap_1 TAP_4516 ();
 sky130_as_sc_hs__tap_1 TAP_4517 ();
 sky130_as_sc_hs__tap_1 TAP_4518 ();
 sky130_as_sc_hs__tap_1 TAP_4519 ();
 sky130_as_sc_hs__tap_1 TAP_452 ();
 sky130_as_sc_hs__tap_1 TAP_4520 ();
 sky130_as_sc_hs__tap_1 TAP_4521 ();
 sky130_as_sc_hs__tap_1 TAP_4522 ();
 sky130_as_sc_hs__tap_1 TAP_4523 ();
 sky130_as_sc_hs__tap_1 TAP_4524 ();
 sky130_as_sc_hs__tap_1 TAP_4525 ();
 sky130_as_sc_hs__tap_1 TAP_4526 ();
 sky130_as_sc_hs__tap_1 TAP_4527 ();
 sky130_as_sc_hs__tap_1 TAP_4528 ();
 sky130_as_sc_hs__tap_1 TAP_4529 ();
 sky130_as_sc_hs__tap_1 TAP_453 ();
 sky130_as_sc_hs__tap_1 TAP_4530 ();
 sky130_as_sc_hs__tap_1 TAP_4531 ();
 sky130_as_sc_hs__tap_1 TAP_4532 ();
 sky130_as_sc_hs__tap_1 TAP_4533 ();
 sky130_as_sc_hs__tap_1 TAP_4534 ();
 sky130_as_sc_hs__tap_1 TAP_4535 ();
 sky130_as_sc_hs__tap_1 TAP_4536 ();
 sky130_as_sc_hs__tap_1 TAP_4537 ();
 sky130_as_sc_hs__tap_1 TAP_4538 ();
 sky130_as_sc_hs__tap_1 TAP_4539 ();
 sky130_as_sc_hs__tap_1 TAP_454 ();
 sky130_as_sc_hs__tap_1 TAP_4540 ();
 sky130_as_sc_hs__tap_1 TAP_4541 ();
 sky130_as_sc_hs__tap_1 TAP_4542 ();
 sky130_as_sc_hs__tap_1 TAP_4543 ();
 sky130_as_sc_hs__tap_1 TAP_4544 ();
 sky130_as_sc_hs__tap_1 TAP_4545 ();
 sky130_as_sc_hs__tap_1 TAP_4546 ();
 sky130_as_sc_hs__tap_1 TAP_4547 ();
 sky130_as_sc_hs__tap_1 TAP_4548 ();
 sky130_as_sc_hs__tap_1 TAP_4549 ();
 sky130_as_sc_hs__tap_1 TAP_455 ();
 sky130_as_sc_hs__tap_1 TAP_4550 ();
 sky130_as_sc_hs__tap_1 TAP_4551 ();
 sky130_as_sc_hs__tap_1 TAP_4552 ();
 sky130_as_sc_hs__tap_1 TAP_4553 ();
 sky130_as_sc_hs__tap_1 TAP_4554 ();
 sky130_as_sc_hs__tap_1 TAP_4555 ();
 sky130_as_sc_hs__tap_1 TAP_4556 ();
 sky130_as_sc_hs__tap_1 TAP_4557 ();
 sky130_as_sc_hs__tap_1 TAP_4558 ();
 sky130_as_sc_hs__tap_1 TAP_4559 ();
 sky130_as_sc_hs__tap_1 TAP_456 ();
 sky130_as_sc_hs__tap_1 TAP_4560 ();
 sky130_as_sc_hs__tap_1 TAP_4561 ();
 sky130_as_sc_hs__tap_1 TAP_4562 ();
 sky130_as_sc_hs__tap_1 TAP_4563 ();
 sky130_as_sc_hs__tap_1 TAP_4564 ();
 sky130_as_sc_hs__tap_1 TAP_4565 ();
 sky130_as_sc_hs__tap_1 TAP_4566 ();
 sky130_as_sc_hs__tap_1 TAP_4567 ();
 sky130_as_sc_hs__tap_1 TAP_4568 ();
 sky130_as_sc_hs__tap_1 TAP_4569 ();
 sky130_as_sc_hs__tap_1 TAP_457 ();
 sky130_as_sc_hs__tap_1 TAP_4570 ();
 sky130_as_sc_hs__tap_1 TAP_4571 ();
 sky130_as_sc_hs__tap_1 TAP_4572 ();
 sky130_as_sc_hs__tap_1 TAP_4573 ();
 sky130_as_sc_hs__tap_1 TAP_4574 ();
 sky130_as_sc_hs__tap_1 TAP_4575 ();
 sky130_as_sc_hs__tap_1 TAP_4576 ();
 sky130_as_sc_hs__tap_1 TAP_4577 ();
 sky130_as_sc_hs__tap_1 TAP_4578 ();
 sky130_as_sc_hs__tap_1 TAP_4579 ();
 sky130_as_sc_hs__tap_1 TAP_458 ();
 sky130_as_sc_hs__tap_1 TAP_4580 ();
 sky130_as_sc_hs__tap_1 TAP_4581 ();
 sky130_as_sc_hs__tap_1 TAP_4582 ();
 sky130_as_sc_hs__tap_1 TAP_4583 ();
 sky130_as_sc_hs__tap_1 TAP_4584 ();
 sky130_as_sc_hs__tap_1 TAP_4585 ();
 sky130_as_sc_hs__tap_1 TAP_4586 ();
 sky130_as_sc_hs__tap_1 TAP_4587 ();
 sky130_as_sc_hs__tap_1 TAP_4588 ();
 sky130_as_sc_hs__tap_1 TAP_4589 ();
 sky130_as_sc_hs__tap_1 TAP_459 ();
 sky130_as_sc_hs__tap_1 TAP_4590 ();
 sky130_as_sc_hs__tap_1 TAP_4591 ();
 sky130_as_sc_hs__tap_1 TAP_4592 ();
 sky130_as_sc_hs__tap_1 TAP_4593 ();
 sky130_as_sc_hs__tap_1 TAP_4594 ();
 sky130_as_sc_hs__tap_1 TAP_4595 ();
 sky130_as_sc_hs__tap_1 TAP_4596 ();
 sky130_as_sc_hs__tap_1 TAP_4597 ();
 sky130_as_sc_hs__tap_1 TAP_4598 ();
 sky130_as_sc_hs__tap_1 TAP_4599 ();
 sky130_as_sc_hs__tap_1 TAP_460 ();
 sky130_as_sc_hs__tap_1 TAP_4600 ();
 sky130_as_sc_hs__tap_1 TAP_4601 ();
 sky130_as_sc_hs__tap_1 TAP_4602 ();
 sky130_as_sc_hs__tap_1 TAP_4603 ();
 sky130_as_sc_hs__tap_1 TAP_4604 ();
 sky130_as_sc_hs__tap_1 TAP_4605 ();
 sky130_as_sc_hs__tap_1 TAP_4606 ();
 sky130_as_sc_hs__tap_1 TAP_4607 ();
 sky130_as_sc_hs__tap_1 TAP_4608 ();
 sky130_as_sc_hs__tap_1 TAP_4609 ();
 sky130_as_sc_hs__tap_1 TAP_461 ();
 sky130_as_sc_hs__tap_1 TAP_4610 ();
 sky130_as_sc_hs__tap_1 TAP_4611 ();
 sky130_as_sc_hs__tap_1 TAP_4612 ();
 sky130_as_sc_hs__tap_1 TAP_4613 ();
 sky130_as_sc_hs__tap_1 TAP_4614 ();
 sky130_as_sc_hs__tap_1 TAP_4615 ();
 sky130_as_sc_hs__tap_1 TAP_4616 ();
 sky130_as_sc_hs__tap_1 TAP_4617 ();
 sky130_as_sc_hs__tap_1 TAP_4618 ();
 sky130_as_sc_hs__tap_1 TAP_4619 ();
 sky130_as_sc_hs__tap_1 TAP_462 ();
 sky130_as_sc_hs__tap_1 TAP_4620 ();
 sky130_as_sc_hs__tap_1 TAP_4621 ();
 sky130_as_sc_hs__tap_1 TAP_4622 ();
 sky130_as_sc_hs__tap_1 TAP_4623 ();
 sky130_as_sc_hs__tap_1 TAP_4624 ();
 sky130_as_sc_hs__tap_1 TAP_4625 ();
 sky130_as_sc_hs__tap_1 TAP_4626 ();
 sky130_as_sc_hs__tap_1 TAP_4627 ();
 sky130_as_sc_hs__tap_1 TAP_4628 ();
 sky130_as_sc_hs__tap_1 TAP_4629 ();
 sky130_as_sc_hs__tap_1 TAP_463 ();
 sky130_as_sc_hs__tap_1 TAP_4630 ();
 sky130_as_sc_hs__tap_1 TAP_4631 ();
 sky130_as_sc_hs__tap_1 TAP_4632 ();
 sky130_as_sc_hs__tap_1 TAP_4633 ();
 sky130_as_sc_hs__tap_1 TAP_4634 ();
 sky130_as_sc_hs__tap_1 TAP_4635 ();
 sky130_as_sc_hs__tap_1 TAP_4636 ();
 sky130_as_sc_hs__tap_1 TAP_4637 ();
 sky130_as_sc_hs__tap_1 TAP_4638 ();
 sky130_as_sc_hs__tap_1 TAP_4639 ();
 sky130_as_sc_hs__tap_1 TAP_464 ();
 sky130_as_sc_hs__tap_1 TAP_4640 ();
 sky130_as_sc_hs__tap_1 TAP_4641 ();
 sky130_as_sc_hs__tap_1 TAP_4642 ();
 sky130_as_sc_hs__tap_1 TAP_4643 ();
 sky130_as_sc_hs__tap_1 TAP_4644 ();
 sky130_as_sc_hs__tap_1 TAP_4645 ();
 sky130_as_sc_hs__tap_1 TAP_4646 ();
 sky130_as_sc_hs__tap_1 TAP_4647 ();
 sky130_as_sc_hs__tap_1 TAP_4648 ();
 sky130_as_sc_hs__tap_1 TAP_4649 ();
 sky130_as_sc_hs__tap_1 TAP_465 ();
 sky130_as_sc_hs__tap_1 TAP_4650 ();
 sky130_as_sc_hs__tap_1 TAP_4651 ();
 sky130_as_sc_hs__tap_1 TAP_4652 ();
 sky130_as_sc_hs__tap_1 TAP_4653 ();
 sky130_as_sc_hs__tap_1 TAP_4654 ();
 sky130_as_sc_hs__tap_1 TAP_4655 ();
 sky130_as_sc_hs__tap_1 TAP_4656 ();
 sky130_as_sc_hs__tap_1 TAP_4657 ();
 sky130_as_sc_hs__tap_1 TAP_4658 ();
 sky130_as_sc_hs__tap_1 TAP_4659 ();
 sky130_as_sc_hs__tap_1 TAP_466 ();
 sky130_as_sc_hs__tap_1 TAP_4660 ();
 sky130_as_sc_hs__tap_1 TAP_4661 ();
 sky130_as_sc_hs__tap_1 TAP_4662 ();
 sky130_as_sc_hs__tap_1 TAP_4663 ();
 sky130_as_sc_hs__tap_1 TAP_4664 ();
 sky130_as_sc_hs__tap_1 TAP_4665 ();
 sky130_as_sc_hs__tap_1 TAP_4666 ();
 sky130_as_sc_hs__tap_1 TAP_4667 ();
 sky130_as_sc_hs__tap_1 TAP_4668 ();
 sky130_as_sc_hs__tap_1 TAP_4669 ();
 sky130_as_sc_hs__tap_1 TAP_467 ();
 sky130_as_sc_hs__tap_1 TAP_4670 ();
 sky130_as_sc_hs__tap_1 TAP_4671 ();
 sky130_as_sc_hs__tap_1 TAP_4672 ();
 sky130_as_sc_hs__tap_1 TAP_4673 ();
 sky130_as_sc_hs__tap_1 TAP_4674 ();
 sky130_as_sc_hs__tap_1 TAP_4675 ();
 sky130_as_sc_hs__tap_1 TAP_4676 ();
 sky130_as_sc_hs__tap_1 TAP_4677 ();
 sky130_as_sc_hs__tap_1 TAP_4678 ();
 sky130_as_sc_hs__tap_1 TAP_4679 ();
 sky130_as_sc_hs__tap_1 TAP_468 ();
 sky130_as_sc_hs__tap_1 TAP_4680 ();
 sky130_as_sc_hs__tap_1 TAP_4681 ();
 sky130_as_sc_hs__tap_1 TAP_4682 ();
 sky130_as_sc_hs__tap_1 TAP_4683 ();
 sky130_as_sc_hs__tap_1 TAP_4684 ();
 sky130_as_sc_hs__tap_1 TAP_4685 ();
 sky130_as_sc_hs__tap_1 TAP_4686 ();
 sky130_as_sc_hs__tap_1 TAP_4687 ();
 sky130_as_sc_hs__tap_1 TAP_4688 ();
 sky130_as_sc_hs__tap_1 TAP_4689 ();
 sky130_as_sc_hs__tap_1 TAP_469 ();
 sky130_as_sc_hs__tap_1 TAP_4690 ();
 sky130_as_sc_hs__tap_1 TAP_4691 ();
 sky130_as_sc_hs__tap_1 TAP_4692 ();
 sky130_as_sc_hs__tap_1 TAP_4693 ();
 sky130_as_sc_hs__tap_1 TAP_4694 ();
 sky130_as_sc_hs__tap_1 TAP_4695 ();
 sky130_as_sc_hs__tap_1 TAP_4696 ();
 sky130_as_sc_hs__tap_1 TAP_4697 ();
 sky130_as_sc_hs__tap_1 TAP_4698 ();
 sky130_as_sc_hs__tap_1 TAP_4699 ();
 sky130_as_sc_hs__tap_1 TAP_470 ();
 sky130_as_sc_hs__tap_1 TAP_4700 ();
 sky130_as_sc_hs__tap_1 TAP_4701 ();
 sky130_as_sc_hs__tap_1 TAP_4702 ();
 sky130_as_sc_hs__tap_1 TAP_4703 ();
 sky130_as_sc_hs__tap_1 TAP_4704 ();
 sky130_as_sc_hs__tap_1 TAP_4705 ();
 sky130_as_sc_hs__tap_1 TAP_4706 ();
 sky130_as_sc_hs__tap_1 TAP_4707 ();
 sky130_as_sc_hs__tap_1 TAP_4708 ();
 sky130_as_sc_hs__tap_1 TAP_4709 ();
 sky130_as_sc_hs__tap_1 TAP_471 ();
 sky130_as_sc_hs__tap_1 TAP_4710 ();
 sky130_as_sc_hs__tap_1 TAP_4711 ();
 sky130_as_sc_hs__tap_1 TAP_4712 ();
 sky130_as_sc_hs__tap_1 TAP_4713 ();
 sky130_as_sc_hs__tap_1 TAP_4714 ();
 sky130_as_sc_hs__tap_1 TAP_4715 ();
 sky130_as_sc_hs__tap_1 TAP_4716 ();
 sky130_as_sc_hs__tap_1 TAP_4717 ();
 sky130_as_sc_hs__tap_1 TAP_4718 ();
 sky130_as_sc_hs__tap_1 TAP_4719 ();
 sky130_as_sc_hs__tap_1 TAP_472 ();
 sky130_as_sc_hs__tap_1 TAP_4720 ();
 sky130_as_sc_hs__tap_1 TAP_4721 ();
 sky130_as_sc_hs__tap_1 TAP_4722 ();
 sky130_as_sc_hs__tap_1 TAP_4723 ();
 sky130_as_sc_hs__tap_1 TAP_4724 ();
 sky130_as_sc_hs__tap_1 TAP_4725 ();
 sky130_as_sc_hs__tap_1 TAP_4726 ();
 sky130_as_sc_hs__tap_1 TAP_4727 ();
 sky130_as_sc_hs__tap_1 TAP_4728 ();
 sky130_as_sc_hs__tap_1 TAP_4729 ();
 sky130_as_sc_hs__tap_1 TAP_473 ();
 sky130_as_sc_hs__tap_1 TAP_4730 ();
 sky130_as_sc_hs__tap_1 TAP_4731 ();
 sky130_as_sc_hs__tap_1 TAP_4732 ();
 sky130_as_sc_hs__tap_1 TAP_4733 ();
 sky130_as_sc_hs__tap_1 TAP_4734 ();
 sky130_as_sc_hs__tap_1 TAP_4735 ();
 sky130_as_sc_hs__tap_1 TAP_4736 ();
 sky130_as_sc_hs__tap_1 TAP_4737 ();
 sky130_as_sc_hs__tap_1 TAP_4738 ();
 sky130_as_sc_hs__tap_1 TAP_4739 ();
 sky130_as_sc_hs__tap_1 TAP_474 ();
 sky130_as_sc_hs__tap_1 TAP_4740 ();
 sky130_as_sc_hs__tap_1 TAP_4741 ();
 sky130_as_sc_hs__tap_1 TAP_4742 ();
 sky130_as_sc_hs__tap_1 TAP_4743 ();
 sky130_as_sc_hs__tap_1 TAP_4744 ();
 sky130_as_sc_hs__tap_1 TAP_4745 ();
 sky130_as_sc_hs__tap_1 TAP_4746 ();
 sky130_as_sc_hs__tap_1 TAP_4747 ();
 sky130_as_sc_hs__tap_1 TAP_4748 ();
 sky130_as_sc_hs__tap_1 TAP_4749 ();
 sky130_as_sc_hs__tap_1 TAP_475 ();
 sky130_as_sc_hs__tap_1 TAP_4750 ();
 sky130_as_sc_hs__tap_1 TAP_4751 ();
 sky130_as_sc_hs__tap_1 TAP_4752 ();
 sky130_as_sc_hs__tap_1 TAP_4753 ();
 sky130_as_sc_hs__tap_1 TAP_4754 ();
 sky130_as_sc_hs__tap_1 TAP_4755 ();
 sky130_as_sc_hs__tap_1 TAP_4756 ();
 sky130_as_sc_hs__tap_1 TAP_4757 ();
 sky130_as_sc_hs__tap_1 TAP_4758 ();
 sky130_as_sc_hs__tap_1 TAP_4759 ();
 sky130_as_sc_hs__tap_1 TAP_476 ();
 sky130_as_sc_hs__tap_1 TAP_4760 ();
 sky130_as_sc_hs__tap_1 TAP_4761 ();
 sky130_as_sc_hs__tap_1 TAP_4762 ();
 sky130_as_sc_hs__tap_1 TAP_4763 ();
 sky130_as_sc_hs__tap_1 TAP_4764 ();
 sky130_as_sc_hs__tap_1 TAP_4765 ();
 sky130_as_sc_hs__tap_1 TAP_4766 ();
 sky130_as_sc_hs__tap_1 TAP_4767 ();
 sky130_as_sc_hs__tap_1 TAP_4768 ();
 sky130_as_sc_hs__tap_1 TAP_4769 ();
 sky130_as_sc_hs__tap_1 TAP_477 ();
 sky130_as_sc_hs__tap_1 TAP_4770 ();
 sky130_as_sc_hs__tap_1 TAP_4771 ();
 sky130_as_sc_hs__tap_1 TAP_4772 ();
 sky130_as_sc_hs__tap_1 TAP_4773 ();
 sky130_as_sc_hs__tap_1 TAP_4774 ();
 sky130_as_sc_hs__tap_1 TAP_4775 ();
 sky130_as_sc_hs__tap_1 TAP_4776 ();
 sky130_as_sc_hs__tap_1 TAP_4777 ();
 sky130_as_sc_hs__tap_1 TAP_4778 ();
 sky130_as_sc_hs__tap_1 TAP_4779 ();
 sky130_as_sc_hs__tap_1 TAP_478 ();
 sky130_as_sc_hs__tap_1 TAP_4780 ();
 sky130_as_sc_hs__tap_1 TAP_4781 ();
 sky130_as_sc_hs__tap_1 TAP_4782 ();
 sky130_as_sc_hs__tap_1 TAP_4783 ();
 sky130_as_sc_hs__tap_1 TAP_4784 ();
 sky130_as_sc_hs__tap_1 TAP_4785 ();
 sky130_as_sc_hs__tap_1 TAP_4786 ();
 sky130_as_sc_hs__tap_1 TAP_4787 ();
 sky130_as_sc_hs__tap_1 TAP_4788 ();
 sky130_as_sc_hs__tap_1 TAP_4789 ();
 sky130_as_sc_hs__tap_1 TAP_479 ();
 sky130_as_sc_hs__tap_1 TAP_4790 ();
 sky130_as_sc_hs__tap_1 TAP_4791 ();
 sky130_as_sc_hs__tap_1 TAP_4792 ();
 sky130_as_sc_hs__tap_1 TAP_4793 ();
 sky130_as_sc_hs__tap_1 TAP_4794 ();
 sky130_as_sc_hs__tap_1 TAP_4795 ();
 sky130_as_sc_hs__tap_1 TAP_4796 ();
 sky130_as_sc_hs__tap_1 TAP_4797 ();
 sky130_as_sc_hs__tap_1 TAP_4798 ();
 sky130_as_sc_hs__tap_1 TAP_4799 ();
 sky130_as_sc_hs__tap_1 TAP_480 ();
 sky130_as_sc_hs__tap_1 TAP_4800 ();
 sky130_as_sc_hs__tap_1 TAP_4801 ();
 sky130_as_sc_hs__tap_1 TAP_4802 ();
 sky130_as_sc_hs__tap_1 TAP_4803 ();
 sky130_as_sc_hs__tap_1 TAP_4804 ();
 sky130_as_sc_hs__tap_1 TAP_4805 ();
 sky130_as_sc_hs__tap_1 TAP_4806 ();
 sky130_as_sc_hs__tap_1 TAP_4807 ();
 sky130_as_sc_hs__tap_1 TAP_4808 ();
 sky130_as_sc_hs__tap_1 TAP_4809 ();
 sky130_as_sc_hs__tap_1 TAP_481 ();
 sky130_as_sc_hs__tap_1 TAP_4810 ();
 sky130_as_sc_hs__tap_1 TAP_4811 ();
 sky130_as_sc_hs__tap_1 TAP_4812 ();
 sky130_as_sc_hs__tap_1 TAP_4813 ();
 sky130_as_sc_hs__tap_1 TAP_4814 ();
 sky130_as_sc_hs__tap_1 TAP_4815 ();
 sky130_as_sc_hs__tap_1 TAP_4816 ();
 sky130_as_sc_hs__tap_1 TAP_4817 ();
 sky130_as_sc_hs__tap_1 TAP_4818 ();
 sky130_as_sc_hs__tap_1 TAP_4819 ();
 sky130_as_sc_hs__tap_1 TAP_482 ();
 sky130_as_sc_hs__tap_1 TAP_4820 ();
 sky130_as_sc_hs__tap_1 TAP_4821 ();
 sky130_as_sc_hs__tap_1 TAP_4822 ();
 sky130_as_sc_hs__tap_1 TAP_4823 ();
 sky130_as_sc_hs__tap_1 TAP_4824 ();
 sky130_as_sc_hs__tap_1 TAP_4825 ();
 sky130_as_sc_hs__tap_1 TAP_4826 ();
 sky130_as_sc_hs__tap_1 TAP_4827 ();
 sky130_as_sc_hs__tap_1 TAP_4828 ();
 sky130_as_sc_hs__tap_1 TAP_4829 ();
 sky130_as_sc_hs__tap_1 TAP_483 ();
 sky130_as_sc_hs__tap_1 TAP_4830 ();
 sky130_as_sc_hs__tap_1 TAP_4831 ();
 sky130_as_sc_hs__tap_1 TAP_4832 ();
 sky130_as_sc_hs__tap_1 TAP_4833 ();
 sky130_as_sc_hs__tap_1 TAP_4834 ();
 sky130_as_sc_hs__tap_1 TAP_4835 ();
 sky130_as_sc_hs__tap_1 TAP_4836 ();
 sky130_as_sc_hs__tap_1 TAP_4837 ();
 sky130_as_sc_hs__tap_1 TAP_4838 ();
 sky130_as_sc_hs__tap_1 TAP_4839 ();
 sky130_as_sc_hs__tap_1 TAP_484 ();
 sky130_as_sc_hs__tap_1 TAP_4840 ();
 sky130_as_sc_hs__tap_1 TAP_4841 ();
 sky130_as_sc_hs__tap_1 TAP_4842 ();
 sky130_as_sc_hs__tap_1 TAP_4843 ();
 sky130_as_sc_hs__tap_1 TAP_4844 ();
 sky130_as_sc_hs__tap_1 TAP_4845 ();
 sky130_as_sc_hs__tap_1 TAP_4846 ();
 sky130_as_sc_hs__tap_1 TAP_4847 ();
 sky130_as_sc_hs__tap_1 TAP_4848 ();
 sky130_as_sc_hs__tap_1 TAP_4849 ();
 sky130_as_sc_hs__tap_1 TAP_485 ();
 sky130_as_sc_hs__tap_1 TAP_4850 ();
 sky130_as_sc_hs__tap_1 TAP_4851 ();
 sky130_as_sc_hs__tap_1 TAP_4852 ();
 sky130_as_sc_hs__tap_1 TAP_4853 ();
 sky130_as_sc_hs__tap_1 TAP_4854 ();
 sky130_as_sc_hs__tap_1 TAP_4855 ();
 sky130_as_sc_hs__tap_1 TAP_4856 ();
 sky130_as_sc_hs__tap_1 TAP_4857 ();
 sky130_as_sc_hs__tap_1 TAP_4858 ();
 sky130_as_sc_hs__tap_1 TAP_4859 ();
 sky130_as_sc_hs__tap_1 TAP_486 ();
 sky130_as_sc_hs__tap_1 TAP_4860 ();
 sky130_as_sc_hs__tap_1 TAP_4861 ();
 sky130_as_sc_hs__tap_1 TAP_4862 ();
 sky130_as_sc_hs__tap_1 TAP_4863 ();
 sky130_as_sc_hs__tap_1 TAP_4864 ();
 sky130_as_sc_hs__tap_1 TAP_4865 ();
 sky130_as_sc_hs__tap_1 TAP_4866 ();
 sky130_as_sc_hs__tap_1 TAP_4867 ();
 sky130_as_sc_hs__tap_1 TAP_4868 ();
 sky130_as_sc_hs__tap_1 TAP_4869 ();
 sky130_as_sc_hs__tap_1 TAP_487 ();
 sky130_as_sc_hs__tap_1 TAP_4870 ();
 sky130_as_sc_hs__tap_1 TAP_4871 ();
 sky130_as_sc_hs__tap_1 TAP_4872 ();
 sky130_as_sc_hs__tap_1 TAP_4873 ();
 sky130_as_sc_hs__tap_1 TAP_4874 ();
 sky130_as_sc_hs__tap_1 TAP_4875 ();
 sky130_as_sc_hs__tap_1 TAP_4876 ();
 sky130_as_sc_hs__tap_1 TAP_4877 ();
 sky130_as_sc_hs__tap_1 TAP_4878 ();
 sky130_as_sc_hs__tap_1 TAP_4879 ();
 sky130_as_sc_hs__tap_1 TAP_488 ();
 sky130_as_sc_hs__tap_1 TAP_4880 ();
 sky130_as_sc_hs__tap_1 TAP_4881 ();
 sky130_as_sc_hs__tap_1 TAP_4882 ();
 sky130_as_sc_hs__tap_1 TAP_4883 ();
 sky130_as_sc_hs__tap_1 TAP_4884 ();
 sky130_as_sc_hs__tap_1 TAP_4885 ();
 sky130_as_sc_hs__tap_1 TAP_4886 ();
 sky130_as_sc_hs__tap_1 TAP_4887 ();
 sky130_as_sc_hs__tap_1 TAP_4888 ();
 sky130_as_sc_hs__tap_1 TAP_4889 ();
 sky130_as_sc_hs__tap_1 TAP_489 ();
 sky130_as_sc_hs__tap_1 TAP_4890 ();
 sky130_as_sc_hs__tap_1 TAP_4891 ();
 sky130_as_sc_hs__tap_1 TAP_4892 ();
 sky130_as_sc_hs__tap_1 TAP_4893 ();
 sky130_as_sc_hs__tap_1 TAP_4894 ();
 sky130_as_sc_hs__tap_1 TAP_4895 ();
 sky130_as_sc_hs__tap_1 TAP_4896 ();
 sky130_as_sc_hs__tap_1 TAP_4897 ();
 sky130_as_sc_hs__tap_1 TAP_4898 ();
 sky130_as_sc_hs__tap_1 TAP_4899 ();
 sky130_as_sc_hs__tap_1 TAP_490 ();
 sky130_as_sc_hs__tap_1 TAP_4900 ();
 sky130_as_sc_hs__tap_1 TAP_4901 ();
 sky130_as_sc_hs__tap_1 TAP_4902 ();
 sky130_as_sc_hs__tap_1 TAP_4903 ();
 sky130_as_sc_hs__tap_1 TAP_4904 ();
 sky130_as_sc_hs__tap_1 TAP_4905 ();
 sky130_as_sc_hs__tap_1 TAP_4906 ();
 sky130_as_sc_hs__tap_1 TAP_4907 ();
 sky130_as_sc_hs__tap_1 TAP_4908 ();
 sky130_as_sc_hs__tap_1 TAP_4909 ();
 sky130_as_sc_hs__tap_1 TAP_491 ();
 sky130_as_sc_hs__tap_1 TAP_4910 ();
 sky130_as_sc_hs__tap_1 TAP_4911 ();
 sky130_as_sc_hs__tap_1 TAP_4912 ();
 sky130_as_sc_hs__tap_1 TAP_4913 ();
 sky130_as_sc_hs__tap_1 TAP_4914 ();
 sky130_as_sc_hs__tap_1 TAP_4915 ();
 sky130_as_sc_hs__tap_1 TAP_4916 ();
 sky130_as_sc_hs__tap_1 TAP_4917 ();
 sky130_as_sc_hs__tap_1 TAP_4918 ();
 sky130_as_sc_hs__tap_1 TAP_4919 ();
 sky130_as_sc_hs__tap_1 TAP_492 ();
 sky130_as_sc_hs__tap_1 TAP_4920 ();
 sky130_as_sc_hs__tap_1 TAP_4921 ();
 sky130_as_sc_hs__tap_1 TAP_4922 ();
 sky130_as_sc_hs__tap_1 TAP_4923 ();
 sky130_as_sc_hs__tap_1 TAP_4924 ();
 sky130_as_sc_hs__tap_1 TAP_4925 ();
 sky130_as_sc_hs__tap_1 TAP_4926 ();
 sky130_as_sc_hs__tap_1 TAP_4927 ();
 sky130_as_sc_hs__tap_1 TAP_4928 ();
 sky130_as_sc_hs__tap_1 TAP_4929 ();
 sky130_as_sc_hs__tap_1 TAP_493 ();
 sky130_as_sc_hs__tap_1 TAP_4930 ();
 sky130_as_sc_hs__tap_1 TAP_4931 ();
 sky130_as_sc_hs__tap_1 TAP_4932 ();
 sky130_as_sc_hs__tap_1 TAP_4933 ();
 sky130_as_sc_hs__tap_1 TAP_4934 ();
 sky130_as_sc_hs__tap_1 TAP_4935 ();
 sky130_as_sc_hs__tap_1 TAP_4936 ();
 sky130_as_sc_hs__tap_1 TAP_4937 ();
 sky130_as_sc_hs__tap_1 TAP_4938 ();
 sky130_as_sc_hs__tap_1 TAP_4939 ();
 sky130_as_sc_hs__tap_1 TAP_494 ();
 sky130_as_sc_hs__tap_1 TAP_4940 ();
 sky130_as_sc_hs__tap_1 TAP_4941 ();
 sky130_as_sc_hs__tap_1 TAP_4942 ();
 sky130_as_sc_hs__tap_1 TAP_4943 ();
 sky130_as_sc_hs__tap_1 TAP_4944 ();
 sky130_as_sc_hs__tap_1 TAP_4945 ();
 sky130_as_sc_hs__tap_1 TAP_4946 ();
 sky130_as_sc_hs__tap_1 TAP_4947 ();
 sky130_as_sc_hs__tap_1 TAP_4948 ();
 sky130_as_sc_hs__tap_1 TAP_4949 ();
 sky130_as_sc_hs__tap_1 TAP_495 ();
 sky130_as_sc_hs__tap_1 TAP_4950 ();
 sky130_as_sc_hs__tap_1 TAP_4951 ();
 sky130_as_sc_hs__tap_1 TAP_4952 ();
 sky130_as_sc_hs__tap_1 TAP_4953 ();
 sky130_as_sc_hs__tap_1 TAP_4954 ();
 sky130_as_sc_hs__tap_1 TAP_4955 ();
 sky130_as_sc_hs__tap_1 TAP_4956 ();
 sky130_as_sc_hs__tap_1 TAP_4957 ();
 sky130_as_sc_hs__tap_1 TAP_4958 ();
 sky130_as_sc_hs__tap_1 TAP_4959 ();
 sky130_as_sc_hs__tap_1 TAP_496 ();
 sky130_as_sc_hs__tap_1 TAP_4960 ();
 sky130_as_sc_hs__tap_1 TAP_4961 ();
 sky130_as_sc_hs__tap_1 TAP_4962 ();
 sky130_as_sc_hs__tap_1 TAP_4963 ();
 sky130_as_sc_hs__tap_1 TAP_4964 ();
 sky130_as_sc_hs__tap_1 TAP_4965 ();
 sky130_as_sc_hs__tap_1 TAP_4966 ();
 sky130_as_sc_hs__tap_1 TAP_4967 ();
 sky130_as_sc_hs__tap_1 TAP_4968 ();
 sky130_as_sc_hs__tap_1 TAP_4969 ();
 sky130_as_sc_hs__tap_1 TAP_497 ();
 sky130_as_sc_hs__tap_1 TAP_4970 ();
 sky130_as_sc_hs__tap_1 TAP_4971 ();
 sky130_as_sc_hs__tap_1 TAP_4972 ();
 sky130_as_sc_hs__tap_1 TAP_4973 ();
 sky130_as_sc_hs__tap_1 TAP_4974 ();
 sky130_as_sc_hs__tap_1 TAP_4975 ();
 sky130_as_sc_hs__tap_1 TAP_4976 ();
 sky130_as_sc_hs__tap_1 TAP_4977 ();
 sky130_as_sc_hs__tap_1 TAP_4978 ();
 sky130_as_sc_hs__tap_1 TAP_4979 ();
 sky130_as_sc_hs__tap_1 TAP_498 ();
 sky130_as_sc_hs__tap_1 TAP_4980 ();
 sky130_as_sc_hs__tap_1 TAP_4981 ();
 sky130_as_sc_hs__tap_1 TAP_4982 ();
 sky130_as_sc_hs__tap_1 TAP_4983 ();
 sky130_as_sc_hs__tap_1 TAP_4984 ();
 sky130_as_sc_hs__tap_1 TAP_4985 ();
 sky130_as_sc_hs__tap_1 TAP_4986 ();
 sky130_as_sc_hs__tap_1 TAP_4987 ();
 sky130_as_sc_hs__tap_1 TAP_4988 ();
 sky130_as_sc_hs__tap_1 TAP_4989 ();
 sky130_as_sc_hs__tap_1 TAP_499 ();
 sky130_as_sc_hs__tap_1 TAP_4990 ();
 sky130_as_sc_hs__tap_1 TAP_4991 ();
 sky130_as_sc_hs__tap_1 TAP_4992 ();
 sky130_as_sc_hs__tap_1 TAP_4993 ();
 sky130_as_sc_hs__tap_1 TAP_4994 ();
 sky130_as_sc_hs__tap_1 TAP_4995 ();
 sky130_as_sc_hs__tap_1 TAP_4996 ();
 sky130_as_sc_hs__tap_1 TAP_4997 ();
 sky130_as_sc_hs__tap_1 TAP_4998 ();
 sky130_as_sc_hs__tap_1 TAP_4999 ();
 sky130_as_sc_hs__tap_1 TAP_500 ();
 sky130_as_sc_hs__tap_1 TAP_5000 ();
 sky130_as_sc_hs__tap_1 TAP_5001 ();
 sky130_as_sc_hs__tap_1 TAP_5002 ();
 sky130_as_sc_hs__tap_1 TAP_5003 ();
 sky130_as_sc_hs__tap_1 TAP_5004 ();
 sky130_as_sc_hs__tap_1 TAP_5005 ();
 sky130_as_sc_hs__tap_1 TAP_5006 ();
 sky130_as_sc_hs__tap_1 TAP_5007 ();
 sky130_as_sc_hs__tap_1 TAP_5008 ();
 sky130_as_sc_hs__tap_1 TAP_5009 ();
 sky130_as_sc_hs__tap_1 TAP_501 ();
 sky130_as_sc_hs__tap_1 TAP_5010 ();
 sky130_as_sc_hs__tap_1 TAP_5011 ();
 sky130_as_sc_hs__tap_1 TAP_5012 ();
 sky130_as_sc_hs__tap_1 TAP_5013 ();
 sky130_as_sc_hs__tap_1 TAP_5014 ();
 sky130_as_sc_hs__tap_1 TAP_5015 ();
 sky130_as_sc_hs__tap_1 TAP_5016 ();
 sky130_as_sc_hs__tap_1 TAP_5017 ();
 sky130_as_sc_hs__tap_1 TAP_5018 ();
 sky130_as_sc_hs__tap_1 TAP_5019 ();
 sky130_as_sc_hs__tap_1 TAP_502 ();
 sky130_as_sc_hs__tap_1 TAP_5020 ();
 sky130_as_sc_hs__tap_1 TAP_5021 ();
 sky130_as_sc_hs__tap_1 TAP_5022 ();
 sky130_as_sc_hs__tap_1 TAP_5023 ();
 sky130_as_sc_hs__tap_1 TAP_5024 ();
 sky130_as_sc_hs__tap_1 TAP_5025 ();
 sky130_as_sc_hs__tap_1 TAP_5026 ();
 sky130_as_sc_hs__tap_1 TAP_5027 ();
 sky130_as_sc_hs__tap_1 TAP_5028 ();
 sky130_as_sc_hs__tap_1 TAP_5029 ();
 sky130_as_sc_hs__tap_1 TAP_503 ();
 sky130_as_sc_hs__tap_1 TAP_5030 ();
 sky130_as_sc_hs__tap_1 TAP_5031 ();
 sky130_as_sc_hs__tap_1 TAP_5032 ();
 sky130_as_sc_hs__tap_1 TAP_5033 ();
 sky130_as_sc_hs__tap_1 TAP_5034 ();
 sky130_as_sc_hs__tap_1 TAP_5035 ();
 sky130_as_sc_hs__tap_1 TAP_5036 ();
 sky130_as_sc_hs__tap_1 TAP_5037 ();
 sky130_as_sc_hs__tap_1 TAP_5038 ();
 sky130_as_sc_hs__tap_1 TAP_5039 ();
 sky130_as_sc_hs__tap_1 TAP_504 ();
 sky130_as_sc_hs__tap_1 TAP_5040 ();
 sky130_as_sc_hs__tap_1 TAP_5041 ();
 sky130_as_sc_hs__tap_1 TAP_5042 ();
 sky130_as_sc_hs__tap_1 TAP_5043 ();
 sky130_as_sc_hs__tap_1 TAP_5044 ();
 sky130_as_sc_hs__tap_1 TAP_5045 ();
 sky130_as_sc_hs__tap_1 TAP_5046 ();
 sky130_as_sc_hs__tap_1 TAP_5047 ();
 sky130_as_sc_hs__tap_1 TAP_5048 ();
 sky130_as_sc_hs__tap_1 TAP_5049 ();
 sky130_as_sc_hs__tap_1 TAP_505 ();
 sky130_as_sc_hs__tap_1 TAP_5050 ();
 sky130_as_sc_hs__tap_1 TAP_5051 ();
 sky130_as_sc_hs__tap_1 TAP_5052 ();
 sky130_as_sc_hs__tap_1 TAP_5053 ();
 sky130_as_sc_hs__tap_1 TAP_5054 ();
 sky130_as_sc_hs__tap_1 TAP_5055 ();
 sky130_as_sc_hs__tap_1 TAP_5056 ();
 sky130_as_sc_hs__tap_1 TAP_5057 ();
 sky130_as_sc_hs__tap_1 TAP_5058 ();
 sky130_as_sc_hs__tap_1 TAP_5059 ();
 sky130_as_sc_hs__tap_1 TAP_506 ();
 sky130_as_sc_hs__tap_1 TAP_5060 ();
 sky130_as_sc_hs__tap_1 TAP_5061 ();
 sky130_as_sc_hs__tap_1 TAP_5062 ();
 sky130_as_sc_hs__tap_1 TAP_5063 ();
 sky130_as_sc_hs__tap_1 TAP_5064 ();
 sky130_as_sc_hs__tap_1 TAP_5065 ();
 sky130_as_sc_hs__tap_1 TAP_5066 ();
 sky130_as_sc_hs__tap_1 TAP_5067 ();
 sky130_as_sc_hs__tap_1 TAP_5068 ();
 sky130_as_sc_hs__tap_1 TAP_5069 ();
 sky130_as_sc_hs__tap_1 TAP_507 ();
 sky130_as_sc_hs__tap_1 TAP_5070 ();
 sky130_as_sc_hs__tap_1 TAP_5071 ();
 sky130_as_sc_hs__tap_1 TAP_5072 ();
 sky130_as_sc_hs__tap_1 TAP_5073 ();
 sky130_as_sc_hs__tap_1 TAP_5074 ();
 sky130_as_sc_hs__tap_1 TAP_5075 ();
 sky130_as_sc_hs__tap_1 TAP_5076 ();
 sky130_as_sc_hs__tap_1 TAP_5077 ();
 sky130_as_sc_hs__tap_1 TAP_5078 ();
 sky130_as_sc_hs__tap_1 TAP_5079 ();
 sky130_as_sc_hs__tap_1 TAP_508 ();
 sky130_as_sc_hs__tap_1 TAP_5080 ();
 sky130_as_sc_hs__tap_1 TAP_5081 ();
 sky130_as_sc_hs__tap_1 TAP_5082 ();
 sky130_as_sc_hs__tap_1 TAP_5083 ();
 sky130_as_sc_hs__tap_1 TAP_5084 ();
 sky130_as_sc_hs__tap_1 TAP_5085 ();
 sky130_as_sc_hs__tap_1 TAP_5086 ();
 sky130_as_sc_hs__tap_1 TAP_5087 ();
 sky130_as_sc_hs__tap_1 TAP_5088 ();
 sky130_as_sc_hs__tap_1 TAP_5089 ();
 sky130_as_sc_hs__tap_1 TAP_509 ();
 sky130_as_sc_hs__tap_1 TAP_5090 ();
 sky130_as_sc_hs__tap_1 TAP_5091 ();
 sky130_as_sc_hs__tap_1 TAP_5092 ();
 sky130_as_sc_hs__tap_1 TAP_5093 ();
 sky130_as_sc_hs__tap_1 TAP_5094 ();
 sky130_as_sc_hs__tap_1 TAP_5095 ();
 sky130_as_sc_hs__tap_1 TAP_5096 ();
 sky130_as_sc_hs__tap_1 TAP_5097 ();
 sky130_as_sc_hs__tap_1 TAP_5098 ();
 sky130_as_sc_hs__tap_1 TAP_5099 ();
 sky130_as_sc_hs__tap_1 TAP_510 ();
 sky130_as_sc_hs__tap_1 TAP_5100 ();
 sky130_as_sc_hs__tap_1 TAP_5101 ();
 sky130_as_sc_hs__tap_1 TAP_5102 ();
 sky130_as_sc_hs__tap_1 TAP_5103 ();
 sky130_as_sc_hs__tap_1 TAP_5104 ();
 sky130_as_sc_hs__tap_1 TAP_5105 ();
 sky130_as_sc_hs__tap_1 TAP_5106 ();
 sky130_as_sc_hs__tap_1 TAP_5107 ();
 sky130_as_sc_hs__tap_1 TAP_5108 ();
 sky130_as_sc_hs__tap_1 TAP_5109 ();
 sky130_as_sc_hs__tap_1 TAP_511 ();
 sky130_as_sc_hs__tap_1 TAP_5110 ();
 sky130_as_sc_hs__tap_1 TAP_5111 ();
 sky130_as_sc_hs__tap_1 TAP_5112 ();
 sky130_as_sc_hs__tap_1 TAP_5113 ();
 sky130_as_sc_hs__tap_1 TAP_5114 ();
 sky130_as_sc_hs__tap_1 TAP_5115 ();
 sky130_as_sc_hs__tap_1 TAP_5116 ();
 sky130_as_sc_hs__tap_1 TAP_5117 ();
 sky130_as_sc_hs__tap_1 TAP_5118 ();
 sky130_as_sc_hs__tap_1 TAP_5119 ();
 sky130_as_sc_hs__tap_1 TAP_512 ();
 sky130_as_sc_hs__tap_1 TAP_5120 ();
 sky130_as_sc_hs__tap_1 TAP_5121 ();
 sky130_as_sc_hs__tap_1 TAP_5122 ();
 sky130_as_sc_hs__tap_1 TAP_5123 ();
 sky130_as_sc_hs__tap_1 TAP_5124 ();
 sky130_as_sc_hs__tap_1 TAP_5125 ();
 sky130_as_sc_hs__tap_1 TAP_5126 ();
 sky130_as_sc_hs__tap_1 TAP_5127 ();
 sky130_as_sc_hs__tap_1 TAP_5128 ();
 sky130_as_sc_hs__tap_1 TAP_5129 ();
 sky130_as_sc_hs__tap_1 TAP_513 ();
 sky130_as_sc_hs__tap_1 TAP_5130 ();
 sky130_as_sc_hs__tap_1 TAP_5131 ();
 sky130_as_sc_hs__tap_1 TAP_5132 ();
 sky130_as_sc_hs__tap_1 TAP_5133 ();
 sky130_as_sc_hs__tap_1 TAP_5134 ();
 sky130_as_sc_hs__tap_1 TAP_5135 ();
 sky130_as_sc_hs__tap_1 TAP_5136 ();
 sky130_as_sc_hs__tap_1 TAP_5137 ();
 sky130_as_sc_hs__tap_1 TAP_5138 ();
 sky130_as_sc_hs__tap_1 TAP_5139 ();
 sky130_as_sc_hs__tap_1 TAP_514 ();
 sky130_as_sc_hs__tap_1 TAP_5140 ();
 sky130_as_sc_hs__tap_1 TAP_5141 ();
 sky130_as_sc_hs__tap_1 TAP_5142 ();
 sky130_as_sc_hs__tap_1 TAP_5143 ();
 sky130_as_sc_hs__tap_1 TAP_5144 ();
 sky130_as_sc_hs__tap_1 TAP_5145 ();
 sky130_as_sc_hs__tap_1 TAP_5146 ();
 sky130_as_sc_hs__tap_1 TAP_5147 ();
 sky130_as_sc_hs__tap_1 TAP_5148 ();
 sky130_as_sc_hs__tap_1 TAP_5149 ();
 sky130_as_sc_hs__tap_1 TAP_515 ();
 sky130_as_sc_hs__tap_1 TAP_5150 ();
 sky130_as_sc_hs__tap_1 TAP_5151 ();
 sky130_as_sc_hs__tap_1 TAP_5152 ();
 sky130_as_sc_hs__tap_1 TAP_5153 ();
 sky130_as_sc_hs__tap_1 TAP_5154 ();
 sky130_as_sc_hs__tap_1 TAP_5155 ();
 sky130_as_sc_hs__tap_1 TAP_5156 ();
 sky130_as_sc_hs__tap_1 TAP_5157 ();
 sky130_as_sc_hs__tap_1 TAP_5158 ();
 sky130_as_sc_hs__tap_1 TAP_5159 ();
 sky130_as_sc_hs__tap_1 TAP_516 ();
 sky130_as_sc_hs__tap_1 TAP_5160 ();
 sky130_as_sc_hs__tap_1 TAP_5161 ();
 sky130_as_sc_hs__tap_1 TAP_5162 ();
 sky130_as_sc_hs__tap_1 TAP_5163 ();
 sky130_as_sc_hs__tap_1 TAP_5164 ();
 sky130_as_sc_hs__tap_1 TAP_5165 ();
 sky130_as_sc_hs__tap_1 TAP_5166 ();
 sky130_as_sc_hs__tap_1 TAP_5167 ();
 sky130_as_sc_hs__tap_1 TAP_5168 ();
 sky130_as_sc_hs__tap_1 TAP_5169 ();
 sky130_as_sc_hs__tap_1 TAP_517 ();
 sky130_as_sc_hs__tap_1 TAP_5170 ();
 sky130_as_sc_hs__tap_1 TAP_5171 ();
 sky130_as_sc_hs__tap_1 TAP_5172 ();
 sky130_as_sc_hs__tap_1 TAP_5173 ();
 sky130_as_sc_hs__tap_1 TAP_5174 ();
 sky130_as_sc_hs__tap_1 TAP_5175 ();
 sky130_as_sc_hs__tap_1 TAP_5176 ();
 sky130_as_sc_hs__tap_1 TAP_5177 ();
 sky130_as_sc_hs__tap_1 TAP_5178 ();
 sky130_as_sc_hs__tap_1 TAP_5179 ();
 sky130_as_sc_hs__tap_1 TAP_518 ();
 sky130_as_sc_hs__tap_1 TAP_5180 ();
 sky130_as_sc_hs__tap_1 TAP_5181 ();
 sky130_as_sc_hs__tap_1 TAP_5182 ();
 sky130_as_sc_hs__tap_1 TAP_5183 ();
 sky130_as_sc_hs__tap_1 TAP_5184 ();
 sky130_as_sc_hs__tap_1 TAP_5185 ();
 sky130_as_sc_hs__tap_1 TAP_5186 ();
 sky130_as_sc_hs__tap_1 TAP_5187 ();
 sky130_as_sc_hs__tap_1 TAP_5188 ();
 sky130_as_sc_hs__tap_1 TAP_5189 ();
 sky130_as_sc_hs__tap_1 TAP_519 ();
 sky130_as_sc_hs__tap_1 TAP_5190 ();
 sky130_as_sc_hs__tap_1 TAP_5191 ();
 sky130_as_sc_hs__tap_1 TAP_5192 ();
 sky130_as_sc_hs__tap_1 TAP_5193 ();
 sky130_as_sc_hs__tap_1 TAP_5194 ();
 sky130_as_sc_hs__tap_1 TAP_5195 ();
 sky130_as_sc_hs__tap_1 TAP_5196 ();
 sky130_as_sc_hs__tap_1 TAP_5197 ();
 sky130_as_sc_hs__tap_1 TAP_5198 ();
 sky130_as_sc_hs__tap_1 TAP_5199 ();
 sky130_as_sc_hs__tap_1 TAP_520 ();
 sky130_as_sc_hs__tap_1 TAP_5200 ();
 sky130_as_sc_hs__tap_1 TAP_5201 ();
 sky130_as_sc_hs__tap_1 TAP_5202 ();
 sky130_as_sc_hs__tap_1 TAP_5203 ();
 sky130_as_sc_hs__tap_1 TAP_5204 ();
 sky130_as_sc_hs__tap_1 TAP_5205 ();
 sky130_as_sc_hs__tap_1 TAP_5206 ();
 sky130_as_sc_hs__tap_1 TAP_5207 ();
 sky130_as_sc_hs__tap_1 TAP_5208 ();
 sky130_as_sc_hs__tap_1 TAP_5209 ();
 sky130_as_sc_hs__tap_1 TAP_521 ();
 sky130_as_sc_hs__tap_1 TAP_5210 ();
 sky130_as_sc_hs__tap_1 TAP_5211 ();
 sky130_as_sc_hs__tap_1 TAP_5212 ();
 sky130_as_sc_hs__tap_1 TAP_5213 ();
 sky130_as_sc_hs__tap_1 TAP_5214 ();
 sky130_as_sc_hs__tap_1 TAP_5215 ();
 sky130_as_sc_hs__tap_1 TAP_5216 ();
 sky130_as_sc_hs__tap_1 TAP_5217 ();
 sky130_as_sc_hs__tap_1 TAP_5218 ();
 sky130_as_sc_hs__tap_1 TAP_5219 ();
 sky130_as_sc_hs__tap_1 TAP_522 ();
 sky130_as_sc_hs__tap_1 TAP_5220 ();
 sky130_as_sc_hs__tap_1 TAP_5221 ();
 sky130_as_sc_hs__tap_1 TAP_5222 ();
 sky130_as_sc_hs__tap_1 TAP_5223 ();
 sky130_as_sc_hs__tap_1 TAP_5224 ();
 sky130_as_sc_hs__tap_1 TAP_5225 ();
 sky130_as_sc_hs__tap_1 TAP_5226 ();
 sky130_as_sc_hs__tap_1 TAP_5227 ();
 sky130_as_sc_hs__tap_1 TAP_5228 ();
 sky130_as_sc_hs__tap_1 TAP_5229 ();
 sky130_as_sc_hs__tap_1 TAP_523 ();
 sky130_as_sc_hs__tap_1 TAP_5230 ();
 sky130_as_sc_hs__tap_1 TAP_5231 ();
 sky130_as_sc_hs__tap_1 TAP_5232 ();
 sky130_as_sc_hs__tap_1 TAP_5233 ();
 sky130_as_sc_hs__tap_1 TAP_5234 ();
 sky130_as_sc_hs__tap_1 TAP_5235 ();
 sky130_as_sc_hs__tap_1 TAP_5236 ();
 sky130_as_sc_hs__tap_1 TAP_5237 ();
 sky130_as_sc_hs__tap_1 TAP_5238 ();
 sky130_as_sc_hs__tap_1 TAP_524 ();
 sky130_as_sc_hs__tap_1 TAP_525 ();
 sky130_as_sc_hs__tap_1 TAP_526 ();
 sky130_as_sc_hs__tap_1 TAP_527 ();
 sky130_as_sc_hs__tap_1 TAP_528 ();
 sky130_as_sc_hs__tap_1 TAP_529 ();
 sky130_as_sc_hs__tap_1 TAP_530 ();
 sky130_as_sc_hs__tap_1 TAP_531 ();
 sky130_as_sc_hs__tap_1 TAP_532 ();
 sky130_as_sc_hs__tap_1 TAP_533 ();
 sky130_as_sc_hs__tap_1 TAP_534 ();
 sky130_as_sc_hs__tap_1 TAP_535 ();
 sky130_as_sc_hs__tap_1 TAP_536 ();
 sky130_as_sc_hs__tap_1 TAP_537 ();
 sky130_as_sc_hs__tap_1 TAP_538 ();
 sky130_as_sc_hs__tap_1 TAP_539 ();
 sky130_as_sc_hs__tap_1 TAP_540 ();
 sky130_as_sc_hs__tap_1 TAP_541 ();
 sky130_as_sc_hs__tap_1 TAP_542 ();
 sky130_as_sc_hs__tap_1 TAP_543 ();
 sky130_as_sc_hs__tap_1 TAP_544 ();
 sky130_as_sc_hs__tap_1 TAP_545 ();
 sky130_as_sc_hs__tap_1 TAP_546 ();
 sky130_as_sc_hs__tap_1 TAP_547 ();
 sky130_as_sc_hs__tap_1 TAP_548 ();
 sky130_as_sc_hs__tap_1 TAP_549 ();
 sky130_as_sc_hs__tap_1 TAP_550 ();
 sky130_as_sc_hs__tap_1 TAP_551 ();
 sky130_as_sc_hs__tap_1 TAP_552 ();
 sky130_as_sc_hs__tap_1 TAP_553 ();
 sky130_as_sc_hs__tap_1 TAP_554 ();
 sky130_as_sc_hs__tap_1 TAP_555 ();
 sky130_as_sc_hs__tap_1 TAP_556 ();
 sky130_as_sc_hs__tap_1 TAP_557 ();
 sky130_as_sc_hs__tap_1 TAP_558 ();
 sky130_as_sc_hs__tap_1 TAP_559 ();
 sky130_as_sc_hs__tap_1 TAP_560 ();
 sky130_as_sc_hs__tap_1 TAP_561 ();
 sky130_as_sc_hs__tap_1 TAP_562 ();
 sky130_as_sc_hs__tap_1 TAP_563 ();
 sky130_as_sc_hs__tap_1 TAP_564 ();
 sky130_as_sc_hs__tap_1 TAP_565 ();
 sky130_as_sc_hs__tap_1 TAP_566 ();
 sky130_as_sc_hs__tap_1 TAP_567 ();
 sky130_as_sc_hs__tap_1 TAP_568 ();
 sky130_as_sc_hs__tap_1 TAP_569 ();
 sky130_as_sc_hs__tap_1 TAP_570 ();
 sky130_as_sc_hs__tap_1 TAP_571 ();
 sky130_as_sc_hs__tap_1 TAP_572 ();
 sky130_as_sc_hs__tap_1 TAP_573 ();
 sky130_as_sc_hs__tap_1 TAP_574 ();
 sky130_as_sc_hs__tap_1 TAP_575 ();
 sky130_as_sc_hs__tap_1 TAP_576 ();
 sky130_as_sc_hs__tap_1 TAP_577 ();
 sky130_as_sc_hs__tap_1 TAP_578 ();
 sky130_as_sc_hs__tap_1 TAP_579 ();
 sky130_as_sc_hs__tap_1 TAP_580 ();
 sky130_as_sc_hs__tap_1 TAP_581 ();
 sky130_as_sc_hs__tap_1 TAP_582 ();
 sky130_as_sc_hs__tap_1 TAP_583 ();
 sky130_as_sc_hs__tap_1 TAP_584 ();
 sky130_as_sc_hs__tap_1 TAP_585 ();
 sky130_as_sc_hs__tap_1 TAP_586 ();
 sky130_as_sc_hs__tap_1 TAP_587 ();
 sky130_as_sc_hs__tap_1 TAP_588 ();
 sky130_as_sc_hs__tap_1 TAP_589 ();
 sky130_as_sc_hs__tap_1 TAP_590 ();
 sky130_as_sc_hs__tap_1 TAP_591 ();
 sky130_as_sc_hs__tap_1 TAP_592 ();
 sky130_as_sc_hs__tap_1 TAP_593 ();
 sky130_as_sc_hs__tap_1 TAP_594 ();
 sky130_as_sc_hs__tap_1 TAP_595 ();
 sky130_as_sc_hs__tap_1 TAP_596 ();
 sky130_as_sc_hs__tap_1 TAP_597 ();
 sky130_as_sc_hs__tap_1 TAP_598 ();
 sky130_as_sc_hs__tap_1 TAP_599 ();
 sky130_as_sc_hs__tap_1 TAP_600 ();
 sky130_as_sc_hs__tap_1 TAP_601 ();
 sky130_as_sc_hs__tap_1 TAP_602 ();
 sky130_as_sc_hs__tap_1 TAP_603 ();
 sky130_as_sc_hs__tap_1 TAP_604 ();
 sky130_as_sc_hs__tap_1 TAP_605 ();
 sky130_as_sc_hs__tap_1 TAP_606 ();
 sky130_as_sc_hs__tap_1 TAP_607 ();
 sky130_as_sc_hs__tap_1 TAP_608 ();
 sky130_as_sc_hs__tap_1 TAP_609 ();
 sky130_as_sc_hs__tap_1 TAP_610 ();
 sky130_as_sc_hs__tap_1 TAP_611 ();
 sky130_as_sc_hs__tap_1 TAP_612 ();
 sky130_as_sc_hs__tap_1 TAP_613 ();
 sky130_as_sc_hs__tap_1 TAP_614 ();
 sky130_as_sc_hs__tap_1 TAP_615 ();
 sky130_as_sc_hs__tap_1 TAP_616 ();
 sky130_as_sc_hs__tap_1 TAP_617 ();
 sky130_as_sc_hs__tap_1 TAP_618 ();
 sky130_as_sc_hs__tap_1 TAP_619 ();
 sky130_as_sc_hs__tap_1 TAP_620 ();
 sky130_as_sc_hs__tap_1 TAP_621 ();
 sky130_as_sc_hs__tap_1 TAP_622 ();
 sky130_as_sc_hs__tap_1 TAP_623 ();
 sky130_as_sc_hs__tap_1 TAP_624 ();
 sky130_as_sc_hs__tap_1 TAP_625 ();
 sky130_as_sc_hs__tap_1 TAP_626 ();
 sky130_as_sc_hs__tap_1 TAP_627 ();
 sky130_as_sc_hs__tap_1 TAP_628 ();
 sky130_as_sc_hs__tap_1 TAP_629 ();
 sky130_as_sc_hs__tap_1 TAP_630 ();
 sky130_as_sc_hs__tap_1 TAP_631 ();
 sky130_as_sc_hs__tap_1 TAP_632 ();
 sky130_as_sc_hs__tap_1 TAP_633 ();
 sky130_as_sc_hs__tap_1 TAP_634 ();
 sky130_as_sc_hs__tap_1 TAP_635 ();
 sky130_as_sc_hs__tap_1 TAP_636 ();
 sky130_as_sc_hs__tap_1 TAP_637 ();
 sky130_as_sc_hs__tap_1 TAP_638 ();
 sky130_as_sc_hs__tap_1 TAP_639 ();
 sky130_as_sc_hs__tap_1 TAP_640 ();
 sky130_as_sc_hs__tap_1 TAP_641 ();
 sky130_as_sc_hs__tap_1 TAP_642 ();
 sky130_as_sc_hs__tap_1 TAP_643 ();
 sky130_as_sc_hs__tap_1 TAP_644 ();
 sky130_as_sc_hs__tap_1 TAP_645 ();
 sky130_as_sc_hs__tap_1 TAP_646 ();
 sky130_as_sc_hs__tap_1 TAP_647 ();
 sky130_as_sc_hs__tap_1 TAP_648 ();
 sky130_as_sc_hs__tap_1 TAP_649 ();
 sky130_as_sc_hs__tap_1 TAP_650 ();
 sky130_as_sc_hs__tap_1 TAP_651 ();
 sky130_as_sc_hs__tap_1 TAP_652 ();
 sky130_as_sc_hs__tap_1 TAP_653 ();
 sky130_as_sc_hs__tap_1 TAP_654 ();
 sky130_as_sc_hs__tap_1 TAP_655 ();
 sky130_as_sc_hs__tap_1 TAP_656 ();
 sky130_as_sc_hs__tap_1 TAP_657 ();
 sky130_as_sc_hs__tap_1 TAP_658 ();
 sky130_as_sc_hs__tap_1 TAP_659 ();
 sky130_as_sc_hs__tap_1 TAP_660 ();
 sky130_as_sc_hs__tap_1 TAP_661 ();
 sky130_as_sc_hs__tap_1 TAP_662 ();
 sky130_as_sc_hs__tap_1 TAP_663 ();
 sky130_as_sc_hs__tap_1 TAP_664 ();
 sky130_as_sc_hs__tap_1 TAP_665 ();
 sky130_as_sc_hs__tap_1 TAP_666 ();
 sky130_as_sc_hs__tap_1 TAP_667 ();
 sky130_as_sc_hs__tap_1 TAP_668 ();
 sky130_as_sc_hs__tap_1 TAP_669 ();
 sky130_as_sc_hs__tap_1 TAP_670 ();
 sky130_as_sc_hs__tap_1 TAP_671 ();
 sky130_as_sc_hs__tap_1 TAP_672 ();
 sky130_as_sc_hs__tap_1 TAP_673 ();
 sky130_as_sc_hs__tap_1 TAP_674 ();
 sky130_as_sc_hs__tap_1 TAP_675 ();
 sky130_as_sc_hs__tap_1 TAP_676 ();
 sky130_as_sc_hs__tap_1 TAP_677 ();
 sky130_as_sc_hs__tap_1 TAP_678 ();
 sky130_as_sc_hs__tap_1 TAP_679 ();
 sky130_as_sc_hs__tap_1 TAP_680 ();
 sky130_as_sc_hs__tap_1 TAP_681 ();
 sky130_as_sc_hs__tap_1 TAP_682 ();
 sky130_as_sc_hs__tap_1 TAP_683 ();
 sky130_as_sc_hs__tap_1 TAP_684 ();
 sky130_as_sc_hs__tap_1 TAP_685 ();
 sky130_as_sc_hs__tap_1 TAP_686 ();
 sky130_as_sc_hs__tap_1 TAP_687 ();
 sky130_as_sc_hs__tap_1 TAP_688 ();
 sky130_as_sc_hs__tap_1 TAP_689 ();
 sky130_as_sc_hs__tap_1 TAP_690 ();
 sky130_as_sc_hs__tap_1 TAP_691 ();
 sky130_as_sc_hs__tap_1 TAP_692 ();
 sky130_as_sc_hs__tap_1 TAP_693 ();
 sky130_as_sc_hs__tap_1 TAP_694 ();
 sky130_as_sc_hs__tap_1 TAP_695 ();
 sky130_as_sc_hs__tap_1 TAP_696 ();
 sky130_as_sc_hs__tap_1 TAP_697 ();
 sky130_as_sc_hs__tap_1 TAP_698 ();
 sky130_as_sc_hs__tap_1 TAP_699 ();
 sky130_as_sc_hs__tap_1 TAP_700 ();
 sky130_as_sc_hs__tap_1 TAP_701 ();
 sky130_as_sc_hs__tap_1 TAP_702 ();
 sky130_as_sc_hs__tap_1 TAP_703 ();
 sky130_as_sc_hs__tap_1 TAP_704 ();
 sky130_as_sc_hs__tap_1 TAP_705 ();
 sky130_as_sc_hs__tap_1 TAP_706 ();
 sky130_as_sc_hs__tap_1 TAP_707 ();
 sky130_as_sc_hs__tap_1 TAP_708 ();
 sky130_as_sc_hs__tap_1 TAP_709 ();
 sky130_as_sc_hs__tap_1 TAP_710 ();
 sky130_as_sc_hs__tap_1 TAP_711 ();
 sky130_as_sc_hs__tap_1 TAP_712 ();
 sky130_as_sc_hs__tap_1 TAP_713 ();
 sky130_as_sc_hs__tap_1 TAP_714 ();
 sky130_as_sc_hs__tap_1 TAP_715 ();
 sky130_as_sc_hs__tap_1 TAP_716 ();
 sky130_as_sc_hs__tap_1 TAP_717 ();
 sky130_as_sc_hs__tap_1 TAP_718 ();
 sky130_as_sc_hs__tap_1 TAP_719 ();
 sky130_as_sc_hs__tap_1 TAP_720 ();
 sky130_as_sc_hs__tap_1 TAP_721 ();
 sky130_as_sc_hs__tap_1 TAP_722 ();
 sky130_as_sc_hs__tap_1 TAP_723 ();
 sky130_as_sc_hs__tap_1 TAP_724 ();
 sky130_as_sc_hs__tap_1 TAP_725 ();
 sky130_as_sc_hs__tap_1 TAP_726 ();
 sky130_as_sc_hs__tap_1 TAP_727 ();
 sky130_as_sc_hs__tap_1 TAP_728 ();
 sky130_as_sc_hs__tap_1 TAP_729 ();
 sky130_as_sc_hs__tap_1 TAP_730 ();
 sky130_as_sc_hs__tap_1 TAP_731 ();
 sky130_as_sc_hs__tap_1 TAP_732 ();
 sky130_as_sc_hs__tap_1 TAP_733 ();
 sky130_as_sc_hs__tap_1 TAP_734 ();
 sky130_as_sc_hs__tap_1 TAP_735 ();
 sky130_as_sc_hs__tap_1 TAP_736 ();
 sky130_as_sc_hs__tap_1 TAP_737 ();
 sky130_as_sc_hs__tap_1 TAP_738 ();
 sky130_as_sc_hs__tap_1 TAP_739 ();
 sky130_as_sc_hs__tap_1 TAP_740 ();
 sky130_as_sc_hs__tap_1 TAP_741 ();
 sky130_as_sc_hs__tap_1 TAP_742 ();
 sky130_as_sc_hs__tap_1 TAP_743 ();
 sky130_as_sc_hs__tap_1 TAP_744 ();
 sky130_as_sc_hs__tap_1 TAP_745 ();
 sky130_as_sc_hs__tap_1 TAP_746 ();
 sky130_as_sc_hs__tap_1 TAP_747 ();
 sky130_as_sc_hs__tap_1 TAP_748 ();
 sky130_as_sc_hs__tap_1 TAP_749 ();
 sky130_as_sc_hs__tap_1 TAP_750 ();
 sky130_as_sc_hs__tap_1 TAP_751 ();
 sky130_as_sc_hs__tap_1 TAP_752 ();
 sky130_as_sc_hs__tap_1 TAP_753 ();
 sky130_as_sc_hs__tap_1 TAP_754 ();
 sky130_as_sc_hs__tap_1 TAP_755 ();
 sky130_as_sc_hs__tap_1 TAP_756 ();
 sky130_as_sc_hs__tap_1 TAP_757 ();
 sky130_as_sc_hs__tap_1 TAP_758 ();
 sky130_as_sc_hs__tap_1 TAP_759 ();
 sky130_as_sc_hs__tap_1 TAP_760 ();
 sky130_as_sc_hs__tap_1 TAP_761 ();
 sky130_as_sc_hs__tap_1 TAP_762 ();
 sky130_as_sc_hs__tap_1 TAP_763 ();
 sky130_as_sc_hs__tap_1 TAP_764 ();
 sky130_as_sc_hs__tap_1 TAP_765 ();
 sky130_as_sc_hs__tap_1 TAP_766 ();
 sky130_as_sc_hs__tap_1 TAP_767 ();
 sky130_as_sc_hs__tap_1 TAP_768 ();
 sky130_as_sc_hs__tap_1 TAP_769 ();
 sky130_as_sc_hs__tap_1 TAP_770 ();
 sky130_as_sc_hs__tap_1 TAP_771 ();
 sky130_as_sc_hs__tap_1 TAP_772 ();
 sky130_as_sc_hs__tap_1 TAP_773 ();
 sky130_as_sc_hs__tap_1 TAP_774 ();
 sky130_as_sc_hs__tap_1 TAP_775 ();
 sky130_as_sc_hs__tap_1 TAP_776 ();
 sky130_as_sc_hs__tap_1 TAP_777 ();
 sky130_as_sc_hs__tap_1 TAP_778 ();
 sky130_as_sc_hs__tap_1 TAP_779 ();
 sky130_as_sc_hs__tap_1 TAP_780 ();
 sky130_as_sc_hs__tap_1 TAP_781 ();
 sky130_as_sc_hs__tap_1 TAP_782 ();
 sky130_as_sc_hs__tap_1 TAP_783 ();
 sky130_as_sc_hs__tap_1 TAP_784 ();
 sky130_as_sc_hs__tap_1 TAP_785 ();
 sky130_as_sc_hs__tap_1 TAP_786 ();
 sky130_as_sc_hs__tap_1 TAP_787 ();
 sky130_as_sc_hs__tap_1 TAP_788 ();
 sky130_as_sc_hs__tap_1 TAP_789 ();
 sky130_as_sc_hs__tap_1 TAP_790 ();
 sky130_as_sc_hs__tap_1 TAP_791 ();
 sky130_as_sc_hs__tap_1 TAP_792 ();
 sky130_as_sc_hs__tap_1 TAP_793 ();
 sky130_as_sc_hs__tap_1 TAP_794 ();
 sky130_as_sc_hs__tap_1 TAP_795 ();
 sky130_as_sc_hs__tap_1 TAP_796 ();
 sky130_as_sc_hs__tap_1 TAP_797 ();
 sky130_as_sc_hs__tap_1 TAP_798 ();
 sky130_as_sc_hs__tap_1 TAP_799 ();
 sky130_as_sc_hs__tap_1 TAP_800 ();
 sky130_as_sc_hs__tap_1 TAP_801 ();
 sky130_as_sc_hs__tap_1 TAP_802 ();
 sky130_as_sc_hs__tap_1 TAP_803 ();
 sky130_as_sc_hs__tap_1 TAP_804 ();
 sky130_as_sc_hs__tap_1 TAP_805 ();
 sky130_as_sc_hs__tap_1 TAP_806 ();
 sky130_as_sc_hs__tap_1 TAP_807 ();
 sky130_as_sc_hs__tap_1 TAP_808 ();
 sky130_as_sc_hs__tap_1 TAP_809 ();
 sky130_as_sc_hs__tap_1 TAP_810 ();
 sky130_as_sc_hs__tap_1 TAP_811 ();
 sky130_as_sc_hs__tap_1 TAP_812 ();
 sky130_as_sc_hs__tap_1 TAP_813 ();
 sky130_as_sc_hs__tap_1 TAP_814 ();
 sky130_as_sc_hs__tap_1 TAP_815 ();
 sky130_as_sc_hs__tap_1 TAP_816 ();
 sky130_as_sc_hs__tap_1 TAP_817 ();
 sky130_as_sc_hs__tap_1 TAP_818 ();
 sky130_as_sc_hs__tap_1 TAP_819 ();
 sky130_as_sc_hs__tap_1 TAP_820 ();
 sky130_as_sc_hs__tap_1 TAP_821 ();
 sky130_as_sc_hs__tap_1 TAP_822 ();
 sky130_as_sc_hs__tap_1 TAP_823 ();
 sky130_as_sc_hs__tap_1 TAP_824 ();
 sky130_as_sc_hs__tap_1 TAP_825 ();
 sky130_as_sc_hs__tap_1 TAP_826 ();
 sky130_as_sc_hs__tap_1 TAP_827 ();
 sky130_as_sc_hs__tap_1 TAP_828 ();
 sky130_as_sc_hs__tap_1 TAP_829 ();
 sky130_as_sc_hs__tap_1 TAP_830 ();
 sky130_as_sc_hs__tap_1 TAP_831 ();
 sky130_as_sc_hs__tap_1 TAP_832 ();
 sky130_as_sc_hs__tap_1 TAP_833 ();
 sky130_as_sc_hs__tap_1 TAP_834 ();
 sky130_as_sc_hs__tap_1 TAP_835 ();
 sky130_as_sc_hs__tap_1 TAP_836 ();
 sky130_as_sc_hs__tap_1 TAP_837 ();
 sky130_as_sc_hs__tap_1 TAP_838 ();
 sky130_as_sc_hs__tap_1 TAP_839 ();
 sky130_as_sc_hs__tap_1 TAP_840 ();
 sky130_as_sc_hs__tap_1 TAP_841 ();
 sky130_as_sc_hs__tap_1 TAP_842 ();
 sky130_as_sc_hs__tap_1 TAP_843 ();
 sky130_as_sc_hs__tap_1 TAP_844 ();
 sky130_as_sc_hs__tap_1 TAP_845 ();
 sky130_as_sc_hs__tap_1 TAP_846 ();
 sky130_as_sc_hs__tap_1 TAP_847 ();
 sky130_as_sc_hs__tap_1 TAP_848 ();
 sky130_as_sc_hs__tap_1 TAP_849 ();
 sky130_as_sc_hs__tap_1 TAP_850 ();
 sky130_as_sc_hs__tap_1 TAP_851 ();
 sky130_as_sc_hs__tap_1 TAP_852 ();
 sky130_as_sc_hs__tap_1 TAP_853 ();
 sky130_as_sc_hs__tap_1 TAP_854 ();
 sky130_as_sc_hs__tap_1 TAP_855 ();
 sky130_as_sc_hs__tap_1 TAP_856 ();
 sky130_as_sc_hs__tap_1 TAP_857 ();
 sky130_as_sc_hs__tap_1 TAP_858 ();
 sky130_as_sc_hs__tap_1 TAP_859 ();
 sky130_as_sc_hs__tap_1 TAP_860 ();
 sky130_as_sc_hs__tap_1 TAP_861 ();
 sky130_as_sc_hs__tap_1 TAP_862 ();
 sky130_as_sc_hs__tap_1 TAP_863 ();
 sky130_as_sc_hs__tap_1 TAP_864 ();
 sky130_as_sc_hs__tap_1 TAP_865 ();
 sky130_as_sc_hs__tap_1 TAP_866 ();
 sky130_as_sc_hs__tap_1 TAP_867 ();
 sky130_as_sc_hs__tap_1 TAP_868 ();
 sky130_as_sc_hs__tap_1 TAP_869 ();
 sky130_as_sc_hs__tap_1 TAP_870 ();
 sky130_as_sc_hs__tap_1 TAP_871 ();
 sky130_as_sc_hs__tap_1 TAP_872 ();
 sky130_as_sc_hs__tap_1 TAP_873 ();
 sky130_as_sc_hs__tap_1 TAP_874 ();
 sky130_as_sc_hs__tap_1 TAP_875 ();
 sky130_as_sc_hs__tap_1 TAP_876 ();
 sky130_as_sc_hs__tap_1 TAP_877 ();
 sky130_as_sc_hs__tap_1 TAP_878 ();
 sky130_as_sc_hs__tap_1 TAP_879 ();
 sky130_as_sc_hs__tap_1 TAP_880 ();
 sky130_as_sc_hs__tap_1 TAP_881 ();
 sky130_as_sc_hs__tap_1 TAP_882 ();
 sky130_as_sc_hs__tap_1 TAP_883 ();
 sky130_as_sc_hs__tap_1 TAP_884 ();
 sky130_as_sc_hs__tap_1 TAP_885 ();
 sky130_as_sc_hs__tap_1 TAP_886 ();
 sky130_as_sc_hs__tap_1 TAP_887 ();
 sky130_as_sc_hs__tap_1 TAP_888 ();
 sky130_as_sc_hs__tap_1 TAP_889 ();
 sky130_as_sc_hs__tap_1 TAP_890 ();
 sky130_as_sc_hs__tap_1 TAP_891 ();
 sky130_as_sc_hs__tap_1 TAP_892 ();
 sky130_as_sc_hs__tap_1 TAP_893 ();
 sky130_as_sc_hs__tap_1 TAP_894 ();
 sky130_as_sc_hs__tap_1 TAP_895 ();
 sky130_as_sc_hs__tap_1 TAP_896 ();
 sky130_as_sc_hs__tap_1 TAP_897 ();
 sky130_as_sc_hs__tap_1 TAP_898 ();
 sky130_as_sc_hs__tap_1 TAP_899 ();
 sky130_as_sc_hs__tap_1 TAP_900 ();
 sky130_as_sc_hs__tap_1 TAP_901 ();
 sky130_as_sc_hs__tap_1 TAP_902 ();
 sky130_as_sc_hs__tap_1 TAP_903 ();
 sky130_as_sc_hs__tap_1 TAP_904 ();
 sky130_as_sc_hs__tap_1 TAP_905 ();
 sky130_as_sc_hs__tap_1 TAP_906 ();
 sky130_as_sc_hs__tap_1 TAP_907 ();
 sky130_as_sc_hs__tap_1 TAP_908 ();
 sky130_as_sc_hs__tap_1 TAP_909 ();
 sky130_as_sc_hs__tap_1 TAP_910 ();
 sky130_as_sc_hs__tap_1 TAP_911 ();
 sky130_as_sc_hs__tap_1 TAP_912 ();
 sky130_as_sc_hs__tap_1 TAP_913 ();
 sky130_as_sc_hs__tap_1 TAP_914 ();
 sky130_as_sc_hs__tap_1 TAP_915 ();
 sky130_as_sc_hs__tap_1 TAP_916 ();
 sky130_as_sc_hs__tap_1 TAP_917 ();
 sky130_as_sc_hs__tap_1 TAP_918 ();
 sky130_as_sc_hs__tap_1 TAP_919 ();
 sky130_as_sc_hs__tap_1 TAP_920 ();
 sky130_as_sc_hs__tap_1 TAP_921 ();
 sky130_as_sc_hs__tap_1 TAP_922 ();
 sky130_as_sc_hs__tap_1 TAP_923 ();
 sky130_as_sc_hs__tap_1 TAP_924 ();
 sky130_as_sc_hs__tap_1 TAP_925 ();
 sky130_as_sc_hs__tap_1 TAP_926 ();
 sky130_as_sc_hs__tap_1 TAP_927 ();
 sky130_as_sc_hs__tap_1 TAP_928 ();
 sky130_as_sc_hs__tap_1 TAP_929 ();
 sky130_as_sc_hs__tap_1 TAP_930 ();
 sky130_as_sc_hs__tap_1 TAP_931 ();
 sky130_as_sc_hs__tap_1 TAP_932 ();
 sky130_as_sc_hs__tap_1 TAP_933 ();
 sky130_as_sc_hs__tap_1 TAP_934 ();
 sky130_as_sc_hs__tap_1 TAP_935 ();
 sky130_as_sc_hs__tap_1 TAP_936 ();
 sky130_as_sc_hs__tap_1 TAP_937 ();
 sky130_as_sc_hs__tap_1 TAP_938 ();
 sky130_as_sc_hs__tap_1 TAP_939 ();
 sky130_as_sc_hs__tap_1 TAP_940 ();
 sky130_as_sc_hs__tap_1 TAP_941 ();
 sky130_as_sc_hs__tap_1 TAP_942 ();
 sky130_as_sc_hs__tap_1 TAP_943 ();
 sky130_as_sc_hs__tap_1 TAP_944 ();
 sky130_as_sc_hs__tap_1 TAP_945 ();
 sky130_as_sc_hs__tap_1 TAP_946 ();
 sky130_as_sc_hs__tap_1 TAP_947 ();
 sky130_as_sc_hs__tap_1 TAP_948 ();
 sky130_as_sc_hs__tap_1 TAP_949 ();
 sky130_as_sc_hs__tap_1 TAP_950 ();
 sky130_as_sc_hs__tap_1 TAP_951 ();
 sky130_as_sc_hs__tap_1 TAP_952 ();
 sky130_as_sc_hs__tap_1 TAP_953 ();
 sky130_as_sc_hs__tap_1 TAP_954 ();
 sky130_as_sc_hs__tap_1 TAP_955 ();
 sky130_as_sc_hs__tap_1 TAP_956 ();
 sky130_as_sc_hs__tap_1 TAP_957 ();
 sky130_as_sc_hs__tap_1 TAP_958 ();
 sky130_as_sc_hs__tap_1 TAP_959 ();
 sky130_as_sc_hs__tap_1 TAP_960 ();
 sky130_as_sc_hs__tap_1 TAP_961 ();
 sky130_as_sc_hs__tap_1 TAP_962 ();
 sky130_as_sc_hs__tap_1 TAP_963 ();
 sky130_as_sc_hs__tap_1 TAP_964 ();
 sky130_as_sc_hs__tap_1 TAP_965 ();
 sky130_as_sc_hs__tap_1 TAP_966 ();
 sky130_as_sc_hs__tap_1 TAP_967 ();
 sky130_as_sc_hs__tap_1 TAP_968 ();
 sky130_as_sc_hs__tap_1 TAP_969 ();
 sky130_as_sc_hs__tap_1 TAP_970 ();
 sky130_as_sc_hs__tap_1 TAP_971 ();
 sky130_as_sc_hs__tap_1 TAP_972 ();
 sky130_as_sc_hs__tap_1 TAP_973 ();
 sky130_as_sc_hs__tap_1 TAP_974 ();
 sky130_as_sc_hs__tap_1 TAP_975 ();
 sky130_as_sc_hs__tap_1 TAP_976 ();
 sky130_as_sc_hs__tap_1 TAP_977 ();
 sky130_as_sc_hs__tap_1 TAP_978 ();
 sky130_as_sc_hs__tap_1 TAP_979 ();
 sky130_as_sc_hs__tap_1 TAP_980 ();
 sky130_as_sc_hs__tap_1 TAP_981 ();
 sky130_as_sc_hs__tap_1 TAP_982 ();
 sky130_as_sc_hs__tap_1 TAP_983 ();
 sky130_as_sc_hs__tap_1 TAP_984 ();
 sky130_as_sc_hs__tap_1 TAP_985 ();
 sky130_as_sc_hs__tap_1 TAP_986 ();
 sky130_as_sc_hs__tap_1 TAP_987 ();
 sky130_as_sc_hs__tap_1 TAP_988 ();
 sky130_as_sc_hs__tap_1 TAP_989 ();
 sky130_as_sc_hs__tap_1 TAP_990 ();
 sky130_as_sc_hs__tap_1 TAP_991 ();
 sky130_as_sc_hs__tap_1 TAP_992 ();
 sky130_as_sc_hs__tap_1 TAP_993 ();
 sky130_as_sc_hs__tap_1 TAP_994 ();
 sky130_as_sc_hs__tap_1 TAP_995 ();
 sky130_as_sc_hs__tap_1 TAP_996 ();
 sky130_as_sc_hs__tap_1 TAP_997 ();
 sky130_as_sc_hs__tap_1 TAP_998 ();
 sky130_as_sc_hs__tap_1 TAP_999 ();
 sky130_as_sc_hs__inv_2 _25938_ (.Y(_19471_),
    .A(\tholin_riscv.PC[2] ));
 sky130_as_sc_hs__inv_2 _25939_ (.Y(net37),
    .A(\tholin_riscv.PORT_dir[5] ));
 sky130_as_sc_hs__inv_2 _25940_ (.Y(_19472_),
    .A(\tholin_riscv.instr[5] ));
 sky130_as_sc_hs__inv_2 _25941_ (.Y(net36),
    .A(\tholin_riscv.PORT_dir[4] ));
 sky130_as_sc_hs__inv_2 _25942_ (.Y(_19473_),
    .A(\tholin_riscv.instr[4] ));
 sky130_as_sc_hs__inv_2 _25943_ (.Y(net35),
    .A(\tholin_riscv.PORT_dir[3] ));
 sky130_as_sc_hs__inv_2 _25944_ (.Y(_19474_),
    .A(\tholin_riscv.instr[3] ));
 sky130_as_sc_hs__inv_2 _25945_ (.Y(net33),
    .A(\tholin_riscv.PORT_dir[2] ));
 sky130_as_sc_hs__inv_2 _25946_ (.Y(_19475_),
    .A(\tholin_riscv.instr[2] ));
 sky130_as_sc_hs__inv_2 _25947_ (.Y(net32),
    .A(\tholin_riscv.PORT_dir[1] ));
 sky130_as_sc_hs__inv_2 _25948_ (.Y(net31),
    .A(\tholin_riscv.PORT_dir[0] ));
 sky130_as_sc_hs__inv_2 _25949_ (.Y(_19476_),
    .A(\tholin_riscv.Bimm[8] ));
 sky130_as_sc_hs__inv_2 _25950_ (.Y(_19477_),
    .A(\tholin_riscv.Bimm[7] ));
 sky130_as_sc_hs__inv_2 _25951_ (.Y(_19478_),
    .A(\tholin_riscv.Iimm[4] ));
 sky130_as_sc_hs__inv_2 _25952_ (.Y(_19479_),
    .A(\tholin_riscv.Iimm[3] ));
 sky130_as_sc_hs__inv_2 _25953_ (.Y(_19480_),
    .A(\tholin_riscv.Iimm[1] ));
 sky130_as_sc_hs__inv_2 _25954_ (.Y(_19481_),
    .A(\tholin_riscv.Jimm[19] ));
 sky130_as_sc_hs__inv_2 _25955_ (.Y(_19482_),
    .A(net340));
 sky130_as_sc_hs__inv_4 _25956_ (.Y(_19483_),
    .A(net346));
 sky130_as_sc_hs__inv_2 _25957_ (.Y(_19484_),
    .A(net361));
 sky130_as_sc_hs__inv_2 _25958_ (.Y(_19485_),
    .A(net390));
 sky130_as_sc_hs__inv_2 _25959_ (.Y(_19486_),
    .A(net1690));
 sky130_as_sc_hs__inv_2 _25960_ (.Y(_19487_),
    .A(\tholin_riscv.Jimm[12] ));
 sky130_as_sc_hs__inv_2 _25961_ (.Y(_19488_),
    .A(\tholin_riscv.instr[6] ));
 sky130_as_sc_hs__inv_2 _25962_ (.Y(_19489_),
    .A(\tholin_riscv.requested_addr[7] ));
 sky130_as_sc_hs__inv_2 _25963_ (.Y(_19490_),
    .A(\tholin_riscv.requested_addr[5] ));
 sky130_as_sc_hs__inv_2 _25964_ (.Y(_19491_),
    .A(\tholin_riscv.requested_addr[4] ));
 sky130_as_sc_hs__inv_2 _25965_ (.Y(_19492_),
    .A(\tholin_riscv.requested_addr[3] ));
 sky130_as_sc_hs__inv_2 _25966_ (.Y(_19493_),
    .A(\tholin_riscv.requested_addr[2] ));
 sky130_as_sc_hs__inv_2 _25967_ (.Y(_19494_),
    .A(\tholin_riscv.is_write ));
 sky130_as_sc_hs__inv_2 _25968_ (.Y(_19495_),
    .A(\tholin_riscv.ret_cycle[1] ));
 sky130_as_sc_hs__inv_2 _25969_ (.Y(_19496_),
    .A(\tholin_riscv.cycle[3] ));
 sky130_as_sc_hs__inv_2 _25970_ (.Y(_19497_),
    .A(\tholin_riscv.cycle[2] ));
 sky130_as_sc_hs__inv_2 _25971_ (.Y(_19498_),
    .A(\tholin_riscv.cycle[0] ));
 sky130_as_sc_hs__inv_2 _25972_ (.Y(_19499_),
    .A(\tholin_riscv.div_shifter[32] ));
 sky130_as_sc_hs__inv_2 _25973_ (.Y(_19500_),
    .A(\tholin_riscv.div_shifter[31] ));
 sky130_as_sc_hs__inv_2 _25974_ (.Y(_19501_),
    .A(\tholin_riscv.div_counter[0] ));
 sky130_as_sc_hs__inv_2 _25975_ (.Y(_19502_),
    .A(\tholin_riscv.uart.divisor[15] ));
 sky130_as_sc_hs__inv_2 _25976_ (.Y(_19503_),
    .A(\tholin_riscv.uart.divisor[14] ));
 sky130_as_sc_hs__inv_2 _25977_ (.Y(_19504_),
    .A(\tholin_riscv.uart.divisor[13] ));
 sky130_as_sc_hs__inv_2 _25978_ (.Y(_19505_),
    .A(\tholin_riscv.uart.divisor[12] ));
 sky130_as_sc_hs__inv_2 _25979_ (.Y(_19506_),
    .A(\tholin_riscv.uart.divisor[10] ));
 sky130_as_sc_hs__inv_2 _25980_ (.Y(_19507_),
    .A(\tholin_riscv.uart.divisor[9] ));
 sky130_as_sc_hs__inv_2 _25981_ (.Y(_19508_),
    .A(\tholin_riscv.uart.divisor[8] ));
 sky130_as_sc_hs__inv_2 _25982_ (.Y(_19509_),
    .A(\tholin_riscv.uart.divisor[7] ));
 sky130_as_sc_hs__inv_2 _25983_ (.Y(_19510_),
    .A(\tholin_riscv.uart.divisor[6] ));
 sky130_as_sc_hs__inv_2 _25984_ (.Y(_19511_),
    .A(\tholin_riscv.uart.divisor[5] ));
 sky130_as_sc_hs__inv_2 _25985_ (.Y(_19512_),
    .A(\tholin_riscv.uart.divisor[4] ));
 sky130_as_sc_hs__inv_2 _25986_ (.Y(_19513_),
    .A(\tholin_riscv.uart.divisor[3] ));
 sky130_as_sc_hs__inv_2 _25987_ (.Y(_19514_),
    .A(\tholin_riscv.uart.divisor[2] ));
 sky130_as_sc_hs__inv_2 _25988_ (.Y(_19515_),
    .A(\tholin_riscv.uart.divisor[1] ));
 sky130_as_sc_hs__inv_2 _25989_ (.Y(_19516_),
    .A(\tholin_riscv.uart.divisor[0] ));
 sky130_as_sc_hs__inv_2 _25990_ (.Y(_19517_),
    .A(\tholin_riscv.spi.data_in_buff[0] ));
 sky130_as_sc_hs__inv_2 _25991_ (.Y(_19518_),
    .A(\tholin_riscv.spi.div_counter[7] ));
 sky130_as_sc_hs__inv_2 _25992_ (.Y(_19519_),
    .A(\tholin_riscv.spi.div_counter[4] ));
 sky130_as_sc_hs__inv_2 _25993_ (.Y(_19520_),
    .A(\tholin_riscv.spi.div_counter[2] ));
 sky130_as_sc_hs__inv_2 _25994_ (.Y(_19521_),
    .A(\tholin_riscv.spi.div_counter[1] ));
 sky130_as_sc_hs__inv_2 _25995_ (.Y(_19522_),
    .A(\tholin_riscv.spi.div_counter[0] ));
 sky130_as_sc_hs__inv_2 _25996_ (.Y(_19523_),
    .A(\tholin_riscv.uart.receive_div_counter[15] ));
 sky130_as_sc_hs__inv_2 _25997_ (.Y(_19524_),
    .A(\tholin_riscv.uart.receive_div_counter[1] ));
 sky130_as_sc_hs__inv_2 _25998_ (.Y(_19525_),
    .A(net1665));
 sky130_as_sc_hs__inv_2 _25999_ (.Y(_19526_),
    .A(\tholin_riscv.uart.div_counter[1] ));
 sky130_as_sc_hs__inv_2 _26000_ (.Y(_19527_),
    .A(net717));
 sky130_as_sc_hs__inv_4 _26001_ (.Y(_19528_),
    .A(net526));
 sky130_as_sc_hs__inv_2 _26002_ (.Y(_19529_),
    .A(net1721));
 sky130_as_sc_hs__inv_2 _26003_ (.Y(_19530_),
    .A(net1694));
 sky130_as_sc_hs__inv_2 _26004_ (.Y(_19531_),
    .A(\tholin_riscv.uart.receiving ));
 sky130_as_sc_hs__inv_2 _26005_ (.Y(_19532_),
    .A(\tholin_riscv.uart.receive_counter[0] ));
 sky130_as_sc_hs__inv_2 _26006_ (.Y(_19533_),
    .A(\tholin_riscv.uart.receive_counter[3] ));
 sky130_as_sc_hs__inv_4 _26007_ (.Y(_19534_),
    .A(net331));
 sky130_as_sc_hs__inv_4 _26008_ (.Y(_19535_),
    .A(net278));
 sky130_as_sc_hs__inv_2 _26009_ (.Y(_19536_),
    .A(net261));
 sky130_as_sc_hs__inv_2 _26010_ (.Y(_19537_),
    .A(net252));
 sky130_as_sc_hs__inv_4 _26011_ (.Y(_19538_),
    .A(net248));
 sky130_as_sc_hs__inv_2 _26012_ (.Y(_19539_),
    .A(\tholin_riscv.regs[1][23] ));
 sky130_as_sc_hs__inv_2 _26013_ (.Y(_19540_),
    .A(\tholin_riscv.regs[3][23] ));
 sky130_as_sc_hs__inv_2 _26014_ (.Y(_19541_),
    .A(\tholin_riscv.regs[5][23] ));
 sky130_as_sc_hs__inv_2 _26015_ (.Y(_19542_),
    .A(\tholin_riscv.regs[7][23] ));
 sky130_as_sc_hs__inv_2 _26016_ (.Y(_19543_),
    .A(\tholin_riscv.regs[9][23] ));
 sky130_as_sc_hs__inv_2 _26017_ (.Y(_19544_),
    .A(\tholin_riscv.regs[11][23] ));
 sky130_as_sc_hs__inv_2 _26018_ (.Y(_19545_),
    .A(\tholin_riscv.regs[13][23] ));
 sky130_as_sc_hs__inv_2 _26019_ (.Y(_19546_),
    .A(\tholin_riscv.regs[15][23] ));
 sky130_as_sc_hs__inv_2 _26020_ (.Y(_19547_),
    .A(\tholin_riscv.regs[17][23] ));
 sky130_as_sc_hs__inv_2 _26021_ (.Y(_19548_),
    .A(\tholin_riscv.regs[19][23] ));
 sky130_as_sc_hs__inv_2 _26022_ (.Y(_19549_),
    .A(\tholin_riscv.regs[21][23] ));
 sky130_as_sc_hs__inv_2 _26023_ (.Y(_19550_),
    .A(\tholin_riscv.regs[23][23] ));
 sky130_as_sc_hs__inv_2 _26024_ (.Y(_19551_),
    .A(\tholin_riscv.regs[25][23] ));
 sky130_as_sc_hs__inv_2 _26025_ (.Y(_19552_),
    .A(\tholin_riscv.regs[27][23] ));
 sky130_as_sc_hs__inv_2 _26026_ (.Y(_19553_),
    .A(\tholin_riscv.regs[29][23] ));
 sky130_as_sc_hs__inv_2 _26027_ (.Y(_19554_),
    .A(\tholin_riscv.regs[31][23] ));
 sky130_as_sc_hs__inv_2 _26028_ (.Y(_19555_),
    .A(\tholin_riscv.regs[1][22] ));
 sky130_as_sc_hs__inv_2 _26029_ (.Y(_19556_),
    .A(\tholin_riscv.regs[3][22] ));
 sky130_as_sc_hs__inv_2 _26030_ (.Y(_19557_),
    .A(\tholin_riscv.regs[5][22] ));
 sky130_as_sc_hs__inv_2 _26031_ (.Y(_19558_),
    .A(\tholin_riscv.regs[7][22] ));
 sky130_as_sc_hs__inv_2 _26032_ (.Y(_19559_),
    .A(\tholin_riscv.regs[9][22] ));
 sky130_as_sc_hs__inv_2 _26033_ (.Y(_19560_),
    .A(\tholin_riscv.regs[11][22] ));
 sky130_as_sc_hs__inv_2 _26034_ (.Y(_19561_),
    .A(\tholin_riscv.regs[13][22] ));
 sky130_as_sc_hs__inv_2 _26035_ (.Y(_19562_),
    .A(\tholin_riscv.regs[15][22] ));
 sky130_as_sc_hs__inv_2 _26036_ (.Y(_19563_),
    .A(\tholin_riscv.regs[17][22] ));
 sky130_as_sc_hs__inv_2 _26037_ (.Y(_19564_),
    .A(\tholin_riscv.regs[19][22] ));
 sky130_as_sc_hs__inv_2 _26038_ (.Y(_19565_),
    .A(\tholin_riscv.regs[21][22] ));
 sky130_as_sc_hs__inv_2 _26039_ (.Y(_19566_),
    .A(\tholin_riscv.regs[23][22] ));
 sky130_as_sc_hs__inv_2 _26040_ (.Y(_19567_),
    .A(\tholin_riscv.regs[25][22] ));
 sky130_as_sc_hs__inv_2 _26041_ (.Y(_19568_),
    .A(\tholin_riscv.regs[27][22] ));
 sky130_as_sc_hs__inv_2 _26042_ (.Y(_19569_),
    .A(\tholin_riscv.regs[29][22] ));
 sky130_as_sc_hs__inv_2 _26043_ (.Y(_19570_),
    .A(\tholin_riscv.regs[31][22] ));
 sky130_as_sc_hs__inv_2 _26044_ (.Y(_19571_),
    .A(\tholin_riscv.regs[1][21] ));
 sky130_as_sc_hs__inv_2 _26045_ (.Y(_19572_),
    .A(\tholin_riscv.regs[3][21] ));
 sky130_as_sc_hs__inv_2 _26046_ (.Y(_19573_),
    .A(\tholin_riscv.regs[5][21] ));
 sky130_as_sc_hs__inv_2 _26047_ (.Y(_19574_),
    .A(\tholin_riscv.regs[7][21] ));
 sky130_as_sc_hs__inv_2 _26048_ (.Y(_19575_),
    .A(\tholin_riscv.regs[9][21] ));
 sky130_as_sc_hs__inv_2 _26049_ (.Y(_19576_),
    .A(\tholin_riscv.regs[11][21] ));
 sky130_as_sc_hs__inv_2 _26050_ (.Y(_19577_),
    .A(\tholin_riscv.regs[13][21] ));
 sky130_as_sc_hs__inv_2 _26051_ (.Y(_19578_),
    .A(\tholin_riscv.regs[15][21] ));
 sky130_as_sc_hs__inv_2 _26052_ (.Y(_19579_),
    .A(\tholin_riscv.regs[17][21] ));
 sky130_as_sc_hs__inv_2 _26053_ (.Y(_19580_),
    .A(\tholin_riscv.regs[19][21] ));
 sky130_as_sc_hs__inv_2 _26054_ (.Y(_19581_),
    .A(\tholin_riscv.regs[21][21] ));
 sky130_as_sc_hs__inv_2 _26055_ (.Y(_19582_),
    .A(\tholin_riscv.regs[23][21] ));
 sky130_as_sc_hs__inv_2 _26056_ (.Y(_19583_),
    .A(\tholin_riscv.regs[25][21] ));
 sky130_as_sc_hs__inv_2 _26057_ (.Y(_19584_),
    .A(\tholin_riscv.regs[27][21] ));
 sky130_as_sc_hs__inv_2 _26058_ (.Y(_19585_),
    .A(\tholin_riscv.regs[29][21] ));
 sky130_as_sc_hs__inv_2 _26059_ (.Y(_19586_),
    .A(\tholin_riscv.regs[31][21] ));
 sky130_as_sc_hs__inv_2 _26060_ (.Y(_19587_),
    .A(\tholin_riscv.regs[1][20] ));
 sky130_as_sc_hs__inv_2 _26061_ (.Y(_19588_),
    .A(\tholin_riscv.regs[3][20] ));
 sky130_as_sc_hs__inv_2 _26062_ (.Y(_19589_),
    .A(\tholin_riscv.regs[5][20] ));
 sky130_as_sc_hs__inv_2 _26063_ (.Y(_19590_),
    .A(\tholin_riscv.regs[7][20] ));
 sky130_as_sc_hs__inv_2 _26064_ (.Y(_19591_),
    .A(\tholin_riscv.regs[9][20] ));
 sky130_as_sc_hs__inv_2 _26065_ (.Y(_19592_),
    .A(\tholin_riscv.regs[11][20] ));
 sky130_as_sc_hs__inv_2 _26066_ (.Y(_19593_),
    .A(\tholin_riscv.regs[13][20] ));
 sky130_as_sc_hs__inv_2 _26067_ (.Y(_19594_),
    .A(\tholin_riscv.regs[15][20] ));
 sky130_as_sc_hs__inv_2 _26068_ (.Y(_19595_),
    .A(\tholin_riscv.regs[17][20] ));
 sky130_as_sc_hs__inv_2 _26069_ (.Y(_19596_),
    .A(\tholin_riscv.regs[19][20] ));
 sky130_as_sc_hs__inv_2 _26070_ (.Y(_19597_),
    .A(\tholin_riscv.regs[21][20] ));
 sky130_as_sc_hs__inv_2 _26071_ (.Y(_19598_),
    .A(\tholin_riscv.regs[23][20] ));
 sky130_as_sc_hs__inv_2 _26072_ (.Y(_19599_),
    .A(\tholin_riscv.regs[25][20] ));
 sky130_as_sc_hs__inv_2 _26073_ (.Y(_19600_),
    .A(\tholin_riscv.regs[27][20] ));
 sky130_as_sc_hs__inv_2 _26074_ (.Y(_19601_),
    .A(\tholin_riscv.regs[29][20] ));
 sky130_as_sc_hs__inv_2 _26075_ (.Y(_19602_),
    .A(\tholin_riscv.regs[31][20] ));
 sky130_as_sc_hs__inv_2 _26076_ (.Y(_19603_),
    .A(\tholin_riscv.regs[1][19] ));
 sky130_as_sc_hs__inv_2 _26077_ (.Y(_19604_),
    .A(\tholin_riscv.regs[3][19] ));
 sky130_as_sc_hs__inv_2 _26078_ (.Y(_19605_),
    .A(\tholin_riscv.regs[5][19] ));
 sky130_as_sc_hs__inv_2 _26079_ (.Y(_19606_),
    .A(\tholin_riscv.regs[7][19] ));
 sky130_as_sc_hs__inv_2 _26080_ (.Y(_19607_),
    .A(\tholin_riscv.regs[9][19] ));
 sky130_as_sc_hs__inv_2 _26081_ (.Y(_19608_),
    .A(\tholin_riscv.regs[11][19] ));
 sky130_as_sc_hs__inv_2 _26082_ (.Y(_19609_),
    .A(\tholin_riscv.regs[13][19] ));
 sky130_as_sc_hs__inv_2 _26083_ (.Y(_19610_),
    .A(\tholin_riscv.regs[15][19] ));
 sky130_as_sc_hs__inv_2 _26084_ (.Y(_19611_),
    .A(\tholin_riscv.regs[17][19] ));
 sky130_as_sc_hs__inv_2 _26085_ (.Y(_19612_),
    .A(\tholin_riscv.regs[19][19] ));
 sky130_as_sc_hs__inv_2 _26086_ (.Y(_19613_),
    .A(\tholin_riscv.regs[21][19] ));
 sky130_as_sc_hs__inv_2 _26087_ (.Y(_19614_),
    .A(\tholin_riscv.regs[23][19] ));
 sky130_as_sc_hs__inv_2 _26088_ (.Y(_19615_),
    .A(\tholin_riscv.regs[25][19] ));
 sky130_as_sc_hs__inv_2 _26089_ (.Y(_19616_),
    .A(\tholin_riscv.regs[27][19] ));
 sky130_as_sc_hs__inv_2 _26090_ (.Y(_19617_),
    .A(\tholin_riscv.regs[29][19] ));
 sky130_as_sc_hs__inv_2 _26091_ (.Y(_19618_),
    .A(\tholin_riscv.regs[31][19] ));
 sky130_as_sc_hs__inv_2 _26092_ (.Y(_19619_),
    .A(\tholin_riscv.regs[1][18] ));
 sky130_as_sc_hs__inv_2 _26093_ (.Y(_19620_),
    .A(\tholin_riscv.regs[3][18] ));
 sky130_as_sc_hs__inv_2 _26094_ (.Y(_19621_),
    .A(\tholin_riscv.regs[5][18] ));
 sky130_as_sc_hs__inv_2 _26095_ (.Y(_19622_),
    .A(\tholin_riscv.regs[7][18] ));
 sky130_as_sc_hs__inv_2 _26096_ (.Y(_19623_),
    .A(\tholin_riscv.regs[9][18] ));
 sky130_as_sc_hs__inv_2 _26097_ (.Y(_19624_),
    .A(\tholin_riscv.regs[11][18] ));
 sky130_as_sc_hs__inv_2 _26098_ (.Y(_19625_),
    .A(\tholin_riscv.regs[13][18] ));
 sky130_as_sc_hs__inv_2 _26099_ (.Y(_19626_),
    .A(\tholin_riscv.regs[15][18] ));
 sky130_as_sc_hs__inv_2 _26100_ (.Y(_19627_),
    .A(\tholin_riscv.regs[17][18] ));
 sky130_as_sc_hs__inv_2 _26101_ (.Y(_19628_),
    .A(\tholin_riscv.regs[19][18] ));
 sky130_as_sc_hs__inv_2 _26102_ (.Y(_19629_),
    .A(\tholin_riscv.regs[21][18] ));
 sky130_as_sc_hs__inv_2 _26103_ (.Y(_19630_),
    .A(\tholin_riscv.regs[23][18] ));
 sky130_as_sc_hs__inv_2 _26104_ (.Y(_19631_),
    .A(\tholin_riscv.regs[25][18] ));
 sky130_as_sc_hs__inv_2 _26105_ (.Y(_19632_),
    .A(\tholin_riscv.regs[27][18] ));
 sky130_as_sc_hs__inv_2 _26106_ (.Y(_19633_),
    .A(\tholin_riscv.regs[29][18] ));
 sky130_as_sc_hs__inv_2 _26107_ (.Y(_19634_),
    .A(\tholin_riscv.regs[31][18] ));
 sky130_as_sc_hs__inv_2 _26108_ (.Y(_19635_),
    .A(\tholin_riscv.regs[1][17] ));
 sky130_as_sc_hs__inv_2 _26109_ (.Y(_19636_),
    .A(\tholin_riscv.regs[3][17] ));
 sky130_as_sc_hs__inv_2 _26110_ (.Y(_19637_),
    .A(\tholin_riscv.regs[5][17] ));
 sky130_as_sc_hs__inv_2 _26111_ (.Y(_19638_),
    .A(\tholin_riscv.regs[7][17] ));
 sky130_as_sc_hs__inv_2 _26112_ (.Y(_19639_),
    .A(\tholin_riscv.regs[9][17] ));
 sky130_as_sc_hs__inv_2 _26113_ (.Y(_19640_),
    .A(\tholin_riscv.regs[11][17] ));
 sky130_as_sc_hs__inv_2 _26114_ (.Y(_19641_),
    .A(\tholin_riscv.regs[13][17] ));
 sky130_as_sc_hs__inv_2 _26115_ (.Y(_19642_),
    .A(\tholin_riscv.regs[15][17] ));
 sky130_as_sc_hs__inv_2 _26116_ (.Y(_19643_),
    .A(\tholin_riscv.regs[17][17] ));
 sky130_as_sc_hs__inv_2 _26117_ (.Y(_19644_),
    .A(\tholin_riscv.regs[19][17] ));
 sky130_as_sc_hs__inv_2 _26118_ (.Y(_19645_),
    .A(\tholin_riscv.regs[21][17] ));
 sky130_as_sc_hs__inv_2 _26119_ (.Y(_19646_),
    .A(\tholin_riscv.regs[23][17] ));
 sky130_as_sc_hs__inv_2 _26120_ (.Y(_19647_),
    .A(\tholin_riscv.regs[25][17] ));
 sky130_as_sc_hs__inv_2 _26121_ (.Y(_19648_),
    .A(\tholin_riscv.regs[27][17] ));
 sky130_as_sc_hs__inv_2 _26122_ (.Y(_19649_),
    .A(\tholin_riscv.regs[29][17] ));
 sky130_as_sc_hs__inv_2 _26123_ (.Y(_19650_),
    .A(\tholin_riscv.regs[31][17] ));
 sky130_as_sc_hs__inv_2 _26124_ (.Y(_19651_),
    .A(\tholin_riscv.regs[1][16] ));
 sky130_as_sc_hs__inv_2 _26125_ (.Y(_19652_),
    .A(\tholin_riscv.regs[3][16] ));
 sky130_as_sc_hs__inv_2 _26126_ (.Y(_19653_),
    .A(\tholin_riscv.regs[5][16] ));
 sky130_as_sc_hs__inv_2 _26127_ (.Y(_19654_),
    .A(\tholin_riscv.regs[7][16] ));
 sky130_as_sc_hs__inv_2 _26128_ (.Y(_19655_),
    .A(\tholin_riscv.regs[9][16] ));
 sky130_as_sc_hs__inv_2 _26129_ (.Y(_19656_),
    .A(\tholin_riscv.regs[11][16] ));
 sky130_as_sc_hs__inv_2 _26130_ (.Y(_19657_),
    .A(\tholin_riscv.regs[13][16] ));
 sky130_as_sc_hs__inv_2 _26131_ (.Y(_19658_),
    .A(\tholin_riscv.regs[15][16] ));
 sky130_as_sc_hs__inv_2 _26132_ (.Y(_19659_),
    .A(\tholin_riscv.regs[17][16] ));
 sky130_as_sc_hs__inv_2 _26133_ (.Y(_19660_),
    .A(\tholin_riscv.regs[19][16] ));
 sky130_as_sc_hs__inv_2 _26134_ (.Y(_19661_),
    .A(\tholin_riscv.regs[21][16] ));
 sky130_as_sc_hs__inv_2 _26135_ (.Y(_19662_),
    .A(\tholin_riscv.regs[23][16] ));
 sky130_as_sc_hs__inv_2 _26136_ (.Y(_19663_),
    .A(\tholin_riscv.regs[25][16] ));
 sky130_as_sc_hs__inv_2 _26137_ (.Y(_19664_),
    .A(\tholin_riscv.regs[27][16] ));
 sky130_as_sc_hs__inv_2 _26138_ (.Y(_19665_),
    .A(\tholin_riscv.regs[29][16] ));
 sky130_as_sc_hs__inv_2 _26139_ (.Y(_19666_),
    .A(\tholin_riscv.regs[31][16] ));
 sky130_as_sc_hs__inv_2 _26140_ (.Y(_19667_),
    .A(\tholin_riscv.regs[1][4] ));
 sky130_as_sc_hs__inv_2 _26141_ (.Y(_19668_),
    .A(\tholin_riscv.regs[3][4] ));
 sky130_as_sc_hs__inv_2 _26142_ (.Y(_19669_),
    .A(\tholin_riscv.regs[5][4] ));
 sky130_as_sc_hs__inv_2 _26143_ (.Y(_19670_),
    .A(\tholin_riscv.regs[7][4] ));
 sky130_as_sc_hs__inv_2 _26144_ (.Y(_19671_),
    .A(\tholin_riscv.regs[9][4] ));
 sky130_as_sc_hs__inv_2 _26145_ (.Y(_19672_),
    .A(\tholin_riscv.regs[11][4] ));
 sky130_as_sc_hs__inv_2 _26146_ (.Y(_19673_),
    .A(\tholin_riscv.regs[13][4] ));
 sky130_as_sc_hs__inv_2 _26147_ (.Y(_19674_),
    .A(\tholin_riscv.regs[15][4] ));
 sky130_as_sc_hs__inv_2 _26148_ (.Y(_19675_),
    .A(\tholin_riscv.regs[17][4] ));
 sky130_as_sc_hs__inv_2 _26149_ (.Y(_19676_),
    .A(\tholin_riscv.regs[19][4] ));
 sky130_as_sc_hs__inv_2 _26150_ (.Y(_19677_),
    .A(\tholin_riscv.regs[21][4] ));
 sky130_as_sc_hs__inv_2 _26151_ (.Y(_19678_),
    .A(\tholin_riscv.regs[23][4] ));
 sky130_as_sc_hs__inv_2 _26152_ (.Y(_19679_),
    .A(\tholin_riscv.regs[25][4] ));
 sky130_as_sc_hs__inv_2 _26153_ (.Y(_19680_),
    .A(\tholin_riscv.regs[27][4] ));
 sky130_as_sc_hs__inv_2 _26154_ (.Y(_19681_),
    .A(\tholin_riscv.regs[29][4] ));
 sky130_as_sc_hs__inv_2 _26155_ (.Y(_19682_),
    .A(\tholin_riscv.regs[31][4] ));
 sky130_as_sc_hs__inv_2 _26156_ (.Y(_19683_),
    .A(\tholin_riscv.tmr1[20] ));
 sky130_as_sc_hs__inv_2 _26157_ (.Y(_19684_),
    .A(\tholin_riscv.tmr0[20] ));
 sky130_as_sc_hs__inv_2 _26158_ (.Y(_19685_),
    .A(net1257));
 sky130_as_sc_hs__inv_2 _26159_ (.Y(_19686_),
    .A(net1286));
 sky130_as_sc_hs__inv_2 _26160_ (.Y(_19687_),
    .A(net818));
 sky130_as_sc_hs__inv_2 _26161_ (.Y(_19688_),
    .A(net971));
 sky130_as_sc_hs__inv_2 _26162_ (.Y(_19689_),
    .A(\tholin_riscv.tmr1[23] ));
 sky130_as_sc_hs__inv_2 _26163_ (.Y(_19690_),
    .A(\tholin_riscv.tmr0[23] ));
 sky130_as_sc_hs__inv_2 _26164_ (.Y(_19691_),
    .A(net1301));
 sky130_as_sc_hs__inv_2 _26165_ (.Y(_19692_),
    .A(net1323));
 sky130_as_sc_hs__inv_2 _26166_ (.Y(_19693_),
    .A(net11));
 sky130_as_sc_hs__inv_2 _26167_ (.Y(_19694_),
    .A(\tholin_riscv.tmr0[31] ));
 sky130_as_sc_hs__inv_2 _26168_ (.Y(_19695_),
    .A(net1042));
 sky130_as_sc_hs__inv_2 _26169_ (.Y(_19696_),
    .A(\tholin_riscv.tmr0[29] ));
 sky130_as_sc_hs__inv_2 _26170_ (.Y(_19697_),
    .A(net923));
 sky130_as_sc_hs__inv_2 _26171_ (.Y(_19698_),
    .A(net1198));
 sky130_as_sc_hs__inv_2 _26172_ (.Y(_19699_),
    .A(\tholin_riscv.tmr0[26] ));
 sky130_as_sc_hs__inv_2 _26173_ (.Y(_19700_),
    .A(net826));
 sky130_as_sc_hs__inv_2 _26174_ (.Y(_19701_),
    .A(net835));
 sky130_as_sc_hs__inv_2 _26175_ (.Y(_19702_),
    .A(net1326));
 sky130_as_sc_hs__inv_2 _26176_ (.Y(_19703_),
    .A(\tholin_riscv.tmr0[17] ));
 sky130_as_sc_hs__inv_2 _26177_ (.Y(_19704_),
    .A(net875));
 sky130_as_sc_hs__inv_2 _26178_ (.Y(_19705_),
    .A(net1211));
 sky130_as_sc_hs__inv_2 _26179_ (.Y(_19706_),
    .A(\tholin_riscv.tmr0[14] ));
 sky130_as_sc_hs__inv_2 _26180_ (.Y(_19707_),
    .A(net794));
 sky130_as_sc_hs__inv_2 _26181_ (.Y(_19708_),
    .A(net1170));
 sky130_as_sc_hs__inv_2 _26182_ (.Y(_19709_),
    .A(\tholin_riscv.tmr0[11] ));
 sky130_as_sc_hs__inv_2 _26183_ (.Y(_19710_),
    .A(net847));
 sky130_as_sc_hs__inv_2 _26184_ (.Y(_19711_),
    .A(net1100));
 sky130_as_sc_hs__inv_2 _26185_ (.Y(_19712_),
    .A(\tholin_riscv.tmr0[8] ));
 sky130_as_sc_hs__inv_2 _26186_ (.Y(_19713_),
    .A(net790));
 sky130_as_sc_hs__inv_2 _26187_ (.Y(_19714_),
    .A(net1082));
 sky130_as_sc_hs__inv_2 _26188_ (.Y(_19715_),
    .A(\tholin_riscv.tmr0[5] ));
 sky130_as_sc_hs__inv_2 _26189_ (.Y(_19716_),
    .A(net806));
 sky130_as_sc_hs__inv_2 _26190_ (.Y(_19717_),
    .A(net1073));
 sky130_as_sc_hs__inv_2 _26191_ (.Y(_19718_),
    .A(\tholin_riscv.tmr0[2] ));
 sky130_as_sc_hs__inv_2 _26192_ (.Y(_19719_),
    .A(\tholin_riscv.tmr0[1] ));
 sky130_as_sc_hs__inv_2 _26193_ (.Y(_19720_),
    .A(\tholin_riscv.tmr0[0] ));
 sky130_as_sc_hs__inv_2 _26194_ (.Y(_19721_),
    .A(\tholin_riscv.tmr1[31] ));
 sky130_as_sc_hs__inv_2 _26195_ (.Y(_19722_),
    .A(net888));
 sky130_as_sc_hs__inv_2 _26196_ (.Y(_19723_),
    .A(\tholin_riscv.tmr1[29] ));
 sky130_as_sc_hs__inv_2 _26197_ (.Y(_19724_),
    .A(net951));
 sky130_as_sc_hs__inv_2 _26198_ (.Y(_19725_),
    .A(net1162));
 sky130_as_sc_hs__inv_2 _26199_ (.Y(_19726_),
    .A(\tholin_riscv.tmr1[26] ));
 sky130_as_sc_hs__inv_2 _26200_ (.Y(_19727_),
    .A(net871));
 sky130_as_sc_hs__inv_2 _26201_ (.Y(_19728_),
    .A(net839));
 sky130_as_sc_hs__inv_2 _26202_ (.Y(_19729_),
    .A(net1334));
 sky130_as_sc_hs__inv_2 _26203_ (.Y(_19730_),
    .A(\tholin_riscv.tmr1[17] ));
 sky130_as_sc_hs__inv_2 _26204_ (.Y(_19731_),
    .A(net830));
 sky130_as_sc_hs__inv_2 _26205_ (.Y(_19732_),
    .A(net1251));
 sky130_as_sc_hs__inv_2 _26206_ (.Y(_19733_),
    .A(\tholin_riscv.tmr1[14] ));
 sky130_as_sc_hs__inv_2 _26207_ (.Y(_19734_),
    .A(net798));
 sky130_as_sc_hs__inv_2 _26208_ (.Y(_19735_),
    .A(net1310));
 sky130_as_sc_hs__inv_2 _26209_ (.Y(_19736_),
    .A(\tholin_riscv.tmr1[11] ));
 sky130_as_sc_hs__inv_2 _26210_ (.Y(_19737_),
    .A(net814));
 sky130_as_sc_hs__inv_2 _26211_ (.Y(_19738_),
    .A(net1069));
 sky130_as_sc_hs__inv_2 _26212_ (.Y(_19739_),
    .A(\tholin_riscv.tmr1[8] ));
 sky130_as_sc_hs__inv_2 _26213_ (.Y(_19740_),
    .A(net855));
 sky130_as_sc_hs__inv_2 _26214_ (.Y(_19741_),
    .A(net1158));
 sky130_as_sc_hs__inv_2 _26215_ (.Y(_19742_),
    .A(\tholin_riscv.tmr1[5] ));
 sky130_as_sc_hs__inv_2 _26216_ (.Y(_19743_),
    .A(net802));
 sky130_as_sc_hs__inv_2 _26217_ (.Y(_19744_),
    .A(net1127));
 sky130_as_sc_hs__inv_2 _26218_ (.Y(_19745_),
    .A(\tholin_riscv.tmr1[2] ));
 sky130_as_sc_hs__inv_2 _26219_ (.Y(_19746_),
    .A(\tholin_riscv.tmr1[1] ));
 sky130_as_sc_hs__inv_2 _26220_ (.Y(_19747_),
    .A(\tholin_riscv.tmr1[0] ));
 sky130_as_sc_hs__and2_2 _26221_ (.A(_19496_),
    .B(\tholin_riscv.cycle[2] ),
    .Y(_19748_));
 sky130_as_sc_hs__nor2_2 _26222_ (.A(\tholin_riscv.cycle[1] ),
    .B(_19498_),
    .Y(_19749_));
 sky130_as_sc_hs__and2_2 _26223_ (.A(_19748_),
    .B(_19749_),
    .Y(_19750_));
 sky130_as_sc_hs__and2_2 _26225_ (.A(\tholin_riscv.cycle[1] ),
    .B(\tholin_riscv.cycle[0] ),
    .Y(_19752_));
 sky130_as_sc_hs__nor2_2 _26226_ (.A(\tholin_riscv.cycle[3] ),
    .B(\tholin_riscv.cycle[2] ),
    .Y(_19753_));
 sky130_as_sc_hs__and2_2 _26227_ (.A(_19752_),
    .B(_19753_),
    .Y(_19754_));
 sky130_as_sc_hs__and2_2 _26229_ (.A(_19751_),
    .B(_19755_),
    .Y(_19756_));
 sky130_as_sc_hs__or2_2 _26230_ (.A(\tholin_riscv.is_write ),
    .B(_19756_),
    .Y(net55));
 sky130_as_sc_hs__or2_2 _26231_ (.A(_19494_),
    .B(_19756_),
    .Y(_19757_));
 sky130_as_sc_hs__and2_2 _26232_ (.A(_19749_),
    .B(_19753_),
    .Y(_19758_));
 sky130_as_sc_hs__nor2_2 _26234_ (.A(\tholin_riscv.cycle[1] ),
    .B(\tholin_riscv.cycle[0] ),
    .Y(_19760_));
 sky130_as_sc_hs__and2_2 _26237_ (.A(\tholin_riscv.cycle[1] ),
    .B(_19498_),
    .Y(_19763_));
 sky130_as_sc_hs__and2_2 _26238_ (.A(_19753_),
    .B(_19763_),
    .Y(_19764_));
 sky130_as_sc_hs__nor2_2 _26239_ (.A(_19762_),
    .B(_19764_),
    .Y(_19765_));
 sky130_as_sc_hs__and2_2 _26240_ (.A(_19757_),
    .B(_19765_),
    .Y(net29));
 sky130_as_sc_hs__and2_2 _26241_ (.A(clknet_leaf_175_wb_clk_i),
    .B(_19764_),
    .Y(net53));
 sky130_as_sc_hs__and2_2 _26242_ (.A(clknet_leaf_175_wb_clk_i),
    .B(_19762_),
    .Y(net52));
 sky130_as_sc_hs__nor2_2 _26243_ (.A(net371),
    .B(\tholin_riscv.io_size[0] ),
    .Y(_19766_));
 sky130_as_sc_hs__or2_2 _26244_ (.A(net371),
    .B(\tholin_riscv.io_size[0] ),
    .Y(_19767_));
 sky130_as_sc_hs__and2_2 _26245_ (.A(\tholin_riscv.requested_addr[0] ),
    .B(_19766_),
    .Y(_19768_));
 sky130_as_sc_hs__or2_2 _26248_ (.A(net2),
    .B(_19770_),
    .Y(_19771_));
 sky130_as_sc_hs__nor2_2 _26249_ (.A(clknet_4_0__leaf_wb_clk_i),
    .B(net1),
    .Y(_19772_));
 sky130_as_sc_hs__nor2_2 _26252_ (.A(_19757_),
    .B(_19774_),
    .Y(_19775_));
 sky130_as_sc_hs__or2_2 _26254_ (.A(\tholin_riscv.requested_addr[0] ),
    .B(_19767_),
    .Y(_19776_));
 sky130_as_sc_hs__and2_2 _26256_ (.A(_19754_),
    .B(_19769_),
    .Y(_19777_));
 sky130_as_sc_hs__and2_2 _26259_ (.A(_19761_),
    .B(_19779_),
    .Y(_19780_));
 sky130_as_sc_hs__and2_2 _26262_ (.A(_19781_),
    .B(_19782_),
    .Y(_19783_));
 sky130_as_sc_hs__nand3_2 _26263_ (.A(_19778_),
    .B(_19780_),
    .C(_19783_),
    .Y(net45));
 sky130_as_sc_hs__and2_2 _26264_ (.A(\tholin_riscv.requested_addr[2] ),
    .B(_19762_),
    .Y(_19784_));
 sky130_as_sc_hs__nand3_2 _26268_ (.A(_19785_),
    .B(_19786_),
    .C(_19787_),
    .Y(_19788_));
 sky130_as_sc_hs__or2_2 _26269_ (.A(_19784_),
    .B(_19788_),
    .Y(net56));
 sky130_as_sc_hs__and2_2 _26271_ (.A(\tholin_riscv.requested_addr[3] ),
    .B(_19762_),
    .Y(_19790_));
 sky130_as_sc_hs__nand3_2 _26274_ (.A(_19789_),
    .B(_19791_),
    .C(_19792_),
    .Y(_19793_));
 sky130_as_sc_hs__or2_2 _26275_ (.A(_19790_),
    .B(_19793_),
    .Y(net63));
 sky130_as_sc_hs__and2_2 _26277_ (.A(\tholin_riscv.requested_addr[4] ),
    .B(_19762_),
    .Y(_19795_));
 sky130_as_sc_hs__nand3_2 _26280_ (.A(_19794_),
    .B(_19796_),
    .C(_19797_),
    .Y(_19798_));
 sky130_as_sc_hs__or2_2 _26281_ (.A(_19795_),
    .B(_19798_),
    .Y(net67));
 sky130_as_sc_hs__and2_2 _26283_ (.A(\tholin_riscv.requested_addr[5] ),
    .B(_19762_),
    .Y(_19800_));
 sky130_as_sc_hs__nand3_2 _26286_ (.A(_19799_),
    .B(_19801_),
    .C(_19802_),
    .Y(_19803_));
 sky130_as_sc_hs__or2_2 _26287_ (.A(_19800_),
    .B(_19803_),
    .Y(net68));
 sky130_as_sc_hs__and2_2 _26289_ (.A(\tholin_riscv.requested_addr[6] ),
    .B(_19762_),
    .Y(_19805_));
 sky130_as_sc_hs__nand3_2 _26292_ (.A(_19804_),
    .B(_19806_),
    .C(_19807_),
    .Y(_19808_));
 sky130_as_sc_hs__or2_2 _26293_ (.A(_19805_),
    .B(_19808_),
    .Y(net69));
 sky130_as_sc_hs__and2_2 _26295_ (.A(\tholin_riscv.requested_addr[7] ),
    .B(_19762_),
    .Y(_19810_));
 sky130_as_sc_hs__nand3_2 _26298_ (.A(_19809_),
    .B(_19811_),
    .C(_19812_),
    .Y(_19813_));
 sky130_as_sc_hs__or2_2 _26299_ (.A(_19810_),
    .B(_19813_),
    .Y(net70));
 sky130_as_sc_hs__and2_2 _26301_ (.A(\tholin_riscv.requested_addr[8] ),
    .B(_19762_),
    .Y(_19815_));
 sky130_as_sc_hs__nand3_2 _26304_ (.A(_19814_),
    .B(_19816_),
    .C(_19817_),
    .Y(_19818_));
 sky130_as_sc_hs__or2_2 _26305_ (.A(_19815_),
    .B(_19818_),
    .Y(net71));
 sky130_as_sc_hs__and2_2 _26306_ (.A(\tholin_riscv.Bimm[1] ),
    .B(_19767_),
    .Y(_19819_));
 sky130_as_sc_hs__and2_2 _26307_ (.A(\tholin_riscv.instr[0] ),
    .B(_19768_),
    .Y(_19820_));
 sky130_as_sc_hs__or2_2 _26308_ (.A(_19819_),
    .B(_19820_),
    .Y(_19821_));
 sky130_as_sc_hs__and2_2 _26313_ (.A(_19824_),
    .B(_19825_),
    .Y(_19826_));
 sky130_as_sc_hs__nand3_2 _26314_ (.A(_19822_),
    .B(_19823_),
    .C(_19826_),
    .Y(net72));
 sky130_as_sc_hs__and2_2 _26315_ (.A(\tholin_riscv.Bimm[2] ),
    .B(_19767_),
    .Y(_19827_));
 sky130_as_sc_hs__and2_2 _26316_ (.A(\tholin_riscv.instr[1] ),
    .B(_19768_),
    .Y(_19828_));
 sky130_as_sc_hs__or2_2 _26317_ (.A(_19827_),
    .B(_19828_),
    .Y(_19829_));
 sky130_as_sc_hs__and2_2 _26322_ (.A(_19832_),
    .B(_19833_),
    .Y(_19834_));
 sky130_as_sc_hs__nand3_2 _26323_ (.A(_19830_),
    .B(_19831_),
    .C(_19834_),
    .Y(net73));
 sky130_as_sc_hs__and2_2 _26324_ (.A(\tholin_riscv.Bimm[3] ),
    .B(_19767_),
    .Y(_19835_));
 sky130_as_sc_hs__and2_2 _26325_ (.A(\tholin_riscv.instr[2] ),
    .B(_19768_),
    .Y(_19836_));
 sky130_as_sc_hs__or2_2 _26326_ (.A(_19835_),
    .B(_19836_),
    .Y(_19837_));
 sky130_as_sc_hs__and2_2 _26331_ (.A(_19840_),
    .B(_19841_),
    .Y(_19842_));
 sky130_as_sc_hs__nand3_2 _26332_ (.A(_19838_),
    .B(_19839_),
    .C(_19842_),
    .Y(net46));
 sky130_as_sc_hs__and2_2 _26333_ (.A(\tholin_riscv.Bimm[4] ),
    .B(_19767_),
    .Y(_19843_));
 sky130_as_sc_hs__and2_2 _26334_ (.A(\tholin_riscv.instr[3] ),
    .B(_19768_),
    .Y(_19844_));
 sky130_as_sc_hs__or2_2 _26335_ (.A(_19843_),
    .B(_19844_),
    .Y(_19845_));
 sky130_as_sc_hs__and2_2 _26340_ (.A(_19848_),
    .B(_19849_),
    .Y(_19850_));
 sky130_as_sc_hs__nand3_2 _26341_ (.A(_19846_),
    .B(_19847_),
    .C(_19850_),
    .Y(net47));
 sky130_as_sc_hs__and2_2 _26342_ (.A(\tholin_riscv.Jimm[12] ),
    .B(_19767_),
    .Y(_19851_));
 sky130_as_sc_hs__and2_2 _26343_ (.A(\tholin_riscv.instr[4] ),
    .B(_19768_),
    .Y(_19852_));
 sky130_as_sc_hs__or2_2 _26344_ (.A(_19851_),
    .B(_19852_),
    .Y(_19853_));
 sky130_as_sc_hs__and2_2 _26349_ (.A(_19856_),
    .B(_19857_),
    .Y(_19858_));
 sky130_as_sc_hs__nand3_2 _26350_ (.A(_19854_),
    .B(_19855_),
    .C(_19858_),
    .Y(net48));
 sky130_as_sc_hs__and2_2 _26351_ (.A(\tholin_riscv.Jimm[13] ),
    .B(_19767_),
    .Y(_19859_));
 sky130_as_sc_hs__and2_2 _26352_ (.A(\tholin_riscv.instr[5] ),
    .B(_19768_),
    .Y(_19860_));
 sky130_as_sc_hs__or2_2 _26353_ (.A(_19859_),
    .B(_19860_),
    .Y(_19861_));
 sky130_as_sc_hs__and2_2 _26358_ (.A(_19864_),
    .B(_19865_),
    .Y(_19866_));
 sky130_as_sc_hs__nand3_2 _26359_ (.A(_19862_),
    .B(_19863_),
    .C(_19866_),
    .Y(net49));
 sky130_as_sc_hs__and2_2 _26360_ (.A(net411),
    .B(_19767_),
    .Y(_19867_));
 sky130_as_sc_hs__and2_2 _26361_ (.A(\tholin_riscv.instr[6] ),
    .B(_19768_),
    .Y(_19868_));
 sky130_as_sc_hs__or2_2 _26362_ (.A(_19867_),
    .B(_19868_),
    .Y(_19869_));
 sky130_as_sc_hs__and2_2 _26367_ (.A(_19872_),
    .B(_19873_),
    .Y(_19874_));
 sky130_as_sc_hs__nand3_2 _26368_ (.A(_19870_),
    .B(_19871_),
    .C(_19874_),
    .Y(net50));
 sky130_as_sc_hs__and2_2 _26369_ (.A(net382),
    .B(_19767_),
    .Y(_19875_));
 sky130_as_sc_hs__and2_2 _26370_ (.A(\tholin_riscv.Bimm[11] ),
    .B(_19766_),
    .Y(_19876_));
 sky130_as_sc_hs__and2_2 _26371_ (.A(\tholin_riscv.requested_addr[0] ),
    .B(_19876_),
    .Y(_19877_));
 sky130_as_sc_hs__or2_2 _26372_ (.A(_19875_),
    .B(_19877_),
    .Y(_19878_));
 sky130_as_sc_hs__nand3_2 _26376_ (.A(_19879_),
    .B(_19880_),
    .C(_19881_),
    .Y(net51));
 sky130_as_sc_hs__and2_2 _26378_ (.A(\tholin_riscv.requested_addr[11] ),
    .B(\tholin_riscv.requested_addr[10] ),
    .Y(_19883_));
 sky130_as_sc_hs__nand3_2 _26379_ (.A(\tholin_riscv.requested_addr[9] ),
    .B(\tholin_riscv.requested_addr[8] ),
    .C(_19883_),
    .Y(_19884_));
 sky130_as_sc_hs__and2_2 _26380_ (.A(\tholin_riscv.requested_addr[15] ),
    .B(\tholin_riscv.requested_addr[14] ),
    .Y(_19885_));
 sky130_as_sc_hs__nand3_2 _26381_ (.A(\tholin_riscv.requested_addr[13] ),
    .B(\tholin_riscv.requested_addr[12] ),
    .C(_19885_),
    .Y(_19886_));
 sky130_as_sc_hs__nor2_2 _26382_ (.A(_19884_),
    .B(_19886_),
    .Y(_19887_));
 sky130_as_sc_hs__and2_2 _26383_ (.A(\tholin_riscv.requested_addr[27] ),
    .B(\tholin_riscv.requested_addr[26] ),
    .Y(_19888_));
 sky130_as_sc_hs__nand3_2 _26384_ (.A(\tholin_riscv.requested_addr[25] ),
    .B(\tholin_riscv.requested_addr[24] ),
    .C(_19888_),
    .Y(_19889_));
 sky130_as_sc_hs__and2_2 _26385_ (.A(\tholin_riscv.requested_addr[31] ),
    .B(\tholin_riscv.requested_addr[30] ),
    .Y(_19890_));
 sky130_as_sc_hs__nand3_2 _26386_ (.A(\tholin_riscv.requested_addr[29] ),
    .B(\tholin_riscv.requested_addr[28] ),
    .C(_19890_),
    .Y(_19891_));
 sky130_as_sc_hs__nor2_2 _26387_ (.A(_19889_),
    .B(_19891_),
    .Y(_19892_));
 sky130_as_sc_hs__and2_2 _26388_ (.A(\tholin_riscv.requested_addr[19] ),
    .B(\tholin_riscv.requested_addr[18] ),
    .Y(_19893_));
 sky130_as_sc_hs__nand3_2 _26389_ (.A(\tholin_riscv.requested_addr[17] ),
    .B(\tholin_riscv.requested_addr[16] ),
    .C(_19893_),
    .Y(_19894_));
 sky130_as_sc_hs__and2_2 _26390_ (.A(\tholin_riscv.requested_addr[23] ),
    .B(\tholin_riscv.requested_addr[22] ),
    .Y(_19895_));
 sky130_as_sc_hs__nand3_2 _26391_ (.A(\tholin_riscv.requested_addr[21] ),
    .B(\tholin_riscv.requested_addr[20] ),
    .C(_19895_),
    .Y(_19896_));
 sky130_as_sc_hs__nor2_2 _26392_ (.A(_19894_),
    .B(_19896_),
    .Y(_19897_));
 sky130_as_sc_hs__and2_2 _26393_ (.A(_19892_),
    .B(_19897_),
    .Y(_19898_));
 sky130_as_sc_hs__nand3_2 _26394_ (.A(_19758_),
    .B(_19887_),
    .C(_19898_),
    .Y(_19899_));
 sky130_as_sc_hs__inv_2 _26395_ (.Y(_19900_),
    .A(_19899_));
 sky130_as_sc_hs__nor2_2 _26396_ (.A(_19494_),
    .B(_19899_),
    .Y(_19901_));
 sky130_as_sc_hs__nor2_2 _26397_ (.A(\tholin_riscv.requested_addr[7] ),
    .B(\tholin_riscv.requested_addr[6] ),
    .Y(_19902_));
 sky130_as_sc_hs__nor2_2 _26398_ (.A(\tholin_riscv.requested_addr[5] ),
    .B(\tholin_riscv.requested_addr[4] ),
    .Y(_19903_));
 sky130_as_sc_hs__and2_2 _26399_ (.A(_19902_),
    .B(_19903_),
    .Y(_19904_));
 sky130_as_sc_hs__and2_2 _26401_ (.A(\tholin_riscv.requested_addr[5] ),
    .B(_19902_),
    .Y(_19906_));
 sky130_as_sc_hs__and2_2 _26402_ (.A(_19491_),
    .B(_19906_),
    .Y(_19907_));
 sky130_as_sc_hs__and2_2 _26403_ (.A(_19492_),
    .B(\tholin_riscv.requested_addr[2] ),
    .Y(_19908_));
 sky130_as_sc_hs__and2_2 _26404_ (.A(_19907_),
    .B(_19908_),
    .Y(_19909_));
 sky130_as_sc_hs__and2_2 _26405_ (.A(_19490_),
    .B(\tholin_riscv.requested_addr[4] ),
    .Y(_19910_));
 sky130_as_sc_hs__and2_2 _26406_ (.A(_19902_),
    .B(_19910_),
    .Y(_19911_));
 sky130_as_sc_hs__and2_2 _26407_ (.A(\tholin_riscv.requested_addr[3] ),
    .B(_19493_),
    .Y(_19912_));
 sky130_as_sc_hs__and2_2 _26408_ (.A(_19907_),
    .B(_19912_),
    .Y(_19913_));
 sky130_as_sc_hs__or2_2 _26409_ (.A(_19909_),
    .B(_19913_),
    .Y(_19914_));
 sky130_as_sc_hs__or2_2 _26410_ (.A(_19911_),
    .B(_19914_),
    .Y(_19915_));
 sky130_as_sc_hs__and2_2 _26411_ (.A(\tholin_riscv.requested_addr[3] ),
    .B(\tholin_riscv.requested_addr[2] ),
    .Y(_19916_));
 sky130_as_sc_hs__and2_2 _26413_ (.A(_19489_),
    .B(\tholin_riscv.requested_addr[6] ),
    .Y(_19918_));
 sky130_as_sc_hs__nor2_2 _26414_ (.A(\tholin_riscv.requested_addr[3] ),
    .B(\tholin_riscv.requested_addr[2] ),
    .Y(_19919_));
 sky130_as_sc_hs__nand3_2 _26415_ (.A(_19910_),
    .B(_19918_),
    .C(_19919_),
    .Y(_19920_));
 sky130_as_sc_hs__and2_2 _26416_ (.A(_19903_),
    .B(_19918_),
    .Y(_19921_));
 sky130_as_sc_hs__nand3_2 _26418_ (.A(_19917_),
    .B(_19920_),
    .C(_19922_),
    .Y(_19923_));
 sky130_as_sc_hs__or2_2 _26419_ (.A(_19915_),
    .B(_19923_),
    .Y(_19924_));
 sky130_as_sc_hs__or2_2 _26420_ (.A(_19904_),
    .B(_19924_),
    .Y(_19925_));
 sky130_as_sc_hs__and2_2 _26422_ (.A(_19882_),
    .B(_19926_),
    .Y(_19927_));
 sky130_as_sc_hs__and2_2 _26423_ (.A(_19907_),
    .B(_19919_),
    .Y(_19928_));
 sky130_as_sc_hs__inv_2 _26424_ (.Y(_19929_),
    .A(_19928_));
 sky130_as_sc_hs__and2_2 _26425_ (.A(_19901_),
    .B(_19928_),
    .Y(_19930_));
 sky130_as_sc_hs__and2_2 _26427_ (.A(\tholin_riscv.cycle[2] ),
    .B(\tholin_riscv.cycle[1] ),
    .Y(_19932_));
 sky130_as_sc_hs__nor2_2 _26428_ (.A(\tholin_riscv.cycle[3] ),
    .B(\tholin_riscv.cycle[0] ),
    .Y(_19933_));
 sky130_as_sc_hs__and2_2 _26429_ (.A(_19932_),
    .B(_19933_),
    .Y(_19934_));
 sky130_as_sc_hs__and2_2 _26431_ (.A(_19753_),
    .B(_19760_),
    .Y(_19936_));
 sky130_as_sc_hs__or2_2 _26433_ (.A(\tholin_riscv.irqs[1] ),
    .B(\tholin_riscv.irqs[2] ),
    .Y(_19938_));
 sky130_as_sc_hs__or2_2 _26434_ (.A(\tholin_riscv.irqs[0] ),
    .B(_19938_),
    .Y(_19939_));
 sky130_as_sc_hs__and2_2 _26435_ (.A(\tholin_riscv.int_enabled ),
    .B(_19939_),
    .Y(_19940_));
 sky130_as_sc_hs__and2_2 _26436_ (.A(_19936_),
    .B(_19940_),
    .Y(_19941_));
 sky130_as_sc_hs__and2_2 _26438_ (.A(_19935_),
    .B(_19942_),
    .Y(_19943_));
 sky130_as_sc_hs__and2_2 _26440_ (.A(\tholin_riscv.instr[5] ),
    .B(\tholin_riscv.instr[6] ),
    .Y(_19945_));
 sky130_as_sc_hs__and2_2 _26441_ (.A(\tholin_riscv.instr[1] ),
    .B(\tholin_riscv.instr[0] ),
    .Y(_19946_));
 sky130_as_sc_hs__and2_2 _26442_ (.A(_19473_),
    .B(\tholin_riscv.instr[2] ),
    .Y(_19947_));
 sky130_as_sc_hs__nand3_2 _26443_ (.A(_19945_),
    .B(_19946_),
    .C(_19947_),
    .Y(_19948_));
 sky130_as_sc_hs__nand3_2 _26446_ (.A(_19751_),
    .B(_19931_),
    .C(_19950_),
    .Y(_19951_));
 sky130_as_sc_hs__and2_2 _26447_ (.A(\tholin_riscv.requested_addr[4] ),
    .B(_19906_),
    .Y(_19952_));
 sky130_as_sc_hs__inv_2 _26448_ (.Y(_19953_),
    .A(_19952_));
 sky130_as_sc_hs__and2_2 _26449_ (.A(_19912_),
    .B(_19952_),
    .Y(_19954_));
 sky130_as_sc_hs__and2_2 _26450_ (.A(_19901_),
    .B(_19954_),
    .Y(_19955_));
 sky130_as_sc_hs__and2_2 _26452_ (.A(_19908_),
    .B(_19952_),
    .Y(_19957_));
 sky130_as_sc_hs__and2_2 _26453_ (.A(_19901_),
    .B(_19957_),
    .Y(_19958_));
 sky130_as_sc_hs__and2_2 _26455_ (.A(_19919_),
    .B(_19952_),
    .Y(_19960_));
 sky130_as_sc_hs__and2_2 _26456_ (.A(_19901_),
    .B(_19960_),
    .Y(_19961_));
 sky130_as_sc_hs__nand3_2 _26458_ (.A(_19956_),
    .B(_19959_),
    .C(_19962_),
    .Y(_19963_));
 sky130_as_sc_hs__or2_2 _26459_ (.A(_19951_),
    .B(_19963_),
    .Y(_19964_));
 sky130_as_sc_hs__nor2_2 _26461_ (.A(\tholin_riscv.instr[2] ),
    .B(_19965_),
    .Y(_19966_));
 sky130_as_sc_hs__and2_2 _26462_ (.A(_19945_),
    .B(_19966_),
    .Y(_19967_));
 sky130_as_sc_hs__inv_2 _26464_ (.Y(_19969_),
    .A(_19968_));
 sky130_as_sc_hs__nor2_2 _26465_ (.A(\tholin_riscv.instr[4] ),
    .B(\tholin_riscv.instr[6] ),
    .Y(_19970_));
 sky130_as_sc_hs__and2_2 _26466_ (.A(_19966_),
    .B(_19970_),
    .Y(_19971_));
 sky130_as_sc_hs__and2_2 _26468_ (.A(_19968_),
    .B(_19972_),
    .Y(_19973_));
 sky130_as_sc_hs__or2_2 _26472_ (.A(_19965_),
    .B(_19976_),
    .Y(_19977_));
 sky130_as_sc_hs__nor2_2 _26473_ (.A(\tholin_riscv.instr[2] ),
    .B(_19977_),
    .Y(_19978_));
 sky130_as_sc_hs__and2_2 _26474_ (.A(\tholin_riscv.instr[5] ),
    .B(_19978_),
    .Y(_19979_));
 sky130_as_sc_hs__nor2_2 _26476_ (.A(net334),
    .B(\tholin_riscv.Bimm[10] ),
    .Y(_19981_));
 sky130_as_sc_hs__nor2_2 _26477_ (.A(\tholin_riscv.Bimm[9] ),
    .B(\tholin_riscv.Bimm[8] ),
    .Y(_19982_));
 sky130_as_sc_hs__and2_2 _26478_ (.A(_19981_),
    .B(_19982_),
    .Y(_19983_));
 sky130_as_sc_hs__nor2_2 _26479_ (.A(\tholin_riscv.Bimm[7] ),
    .B(\tholin_riscv.Bimm[6] ),
    .Y(_19984_));
 sky130_as_sc_hs__and2_2 _26480_ (.A(\tholin_riscv.Bimm[5] ),
    .B(_19984_),
    .Y(_19985_));
 sky130_as_sc_hs__and2_2 _26481_ (.A(_19983_),
    .B(_19985_),
    .Y(_19986_));
 sky130_as_sc_hs__and2_2 _26482_ (.A(_19979_),
    .B(_19986_),
    .Y(_19987_));
 sky130_as_sc_hs__and2_2 _26484_ (.A(\tholin_riscv.instr[4] ),
    .B(_19967_),
    .Y(_19989_));
 sky130_as_sc_hs__nand3_2 _26489_ (.A(_19901_),
    .B(_19916_),
    .C(_19921_),
    .Y(_19994_));
 sky130_as_sc_hs__or2_2 _26490_ (.A(_19758_),
    .B(_19764_),
    .Y(_19995_));
 sky130_as_sc_hs__or2_2 _26492_ (.A(_19937_),
    .B(_19940_),
    .Y(_19997_));
 sky130_as_sc_hs__and2_2 _26493_ (.A(_19920_),
    .B(_19993_),
    .Y(_19998_));
 sky130_as_sc_hs__nand3_2 _26494_ (.A(_19922_),
    .B(_19953_),
    .C(_19998_),
    .Y(_19999_));
 sky130_as_sc_hs__and2_2 _26495_ (.A(_19907_),
    .B(_19916_),
    .Y(_20000_));
 sky130_as_sc_hs__nor2_2 _26496_ (.A(_19905_),
    .B(_19912_),
    .Y(_20001_));
 sky130_as_sc_hs__or2_2 _26497_ (.A(_20000_),
    .B(_20001_),
    .Y(_20002_));
 sky130_as_sc_hs__or2_2 _26498_ (.A(_19999_),
    .B(_20002_),
    .Y(_20003_));
 sky130_as_sc_hs__nor2_2 _26499_ (.A(_19915_),
    .B(_20003_),
    .Y(_20004_));
 sky130_as_sc_hs__inv_2 _26501_ (.Y(_20006_),
    .A(_20005_));
 sky130_as_sc_hs__nand3_2 _26502_ (.A(_19900_),
    .B(_19929_),
    .C(_19993_),
    .Y(_20007_));
 sky130_as_sc_hs__nor2_2 _26503_ (.A(_20005_),
    .B(_20007_),
    .Y(_20008_));
 sky130_as_sc_hs__nor2_2 _26504_ (.A(_19971_),
    .B(_19987_),
    .Y(_20009_));
 sky130_as_sc_hs__and2_2 _26505_ (.A(net145),
    .B(_19990_),
    .Y(_20010_));
 sky130_as_sc_hs__and2_2 _26506_ (.A(_19948_),
    .B(_20010_),
    .Y(_20011_));
 sky130_as_sc_hs__and2_2 _26507_ (.A(_20009_),
    .B(_20011_),
    .Y(_20012_));
 sky130_as_sc_hs__nand3_2 _26509_ (.A(_19761_),
    .B(_19992_),
    .C(_19997_),
    .Y(_20014_));
 sky130_as_sc_hs__nor2_2 _26510_ (.A(_20008_),
    .B(_20014_),
    .Y(_20015_));
 sky130_as_sc_hs__nand3_2 _26511_ (.A(_19496_),
    .B(_19975_),
    .C(_19996_),
    .Y(_20016_));
 sky130_as_sc_hs__nor2_2 _26512_ (.A(_19964_),
    .B(_20016_),
    .Y(_20017_));
 sky130_as_sc_hs__and2_2 _26513_ (.A(_20015_),
    .B(_20017_),
    .Y(_20018_));
 sky130_as_sc_hs__and2_2 _26514_ (.A(_19994_),
    .B(_20013_),
    .Y(_20019_));
 sky130_as_sc_hs__and2_2 _26515_ (.A(_19927_),
    .B(_20019_),
    .Y(_20020_));
 sky130_as_sc_hs__and2_2 _26516_ (.A(_20018_),
    .B(_20020_),
    .Y(_20021_));
 sky130_as_sc_hs__and2_2 _26521_ (.A(_20024_),
    .B(_20025_),
    .Y(_20026_));
 sky130_as_sc_hs__nand3_2 _26522_ (.A(_20022_),
    .B(_20023_),
    .C(_20026_),
    .Y(_20027_));
 sky130_as_sc_hs__and2_2 _26523_ (.A(_19916_),
    .B(_19952_),
    .Y(_20028_));
 sky130_as_sc_hs__and2_2 _26527_ (.A(_19919_),
    .B(_19921_),
    .Y(_20032_));
 sky130_as_sc_hs__and2_2 _26529_ (.A(_19912_),
    .B(_19921_),
    .Y(_20034_));
 sky130_as_sc_hs__nand3_2 _26531_ (.A(_19920_),
    .B(_20033_),
    .C(_20035_),
    .Y(_20036_));
 sky130_as_sc_hs__or2_2 _26532_ (.A(_20031_),
    .B(_20036_),
    .Y(_20037_));
 sky130_as_sc_hs__or2_2 _26533_ (.A(_20027_),
    .B(_20037_),
    .Y(_20038_));
 sky130_as_sc_hs__nor2_2 _26535_ (.A(_19508_),
    .B(_20039_),
    .Y(_20040_));
 sky130_as_sc_hs__or2_2 _26536_ (.A(_20038_),
    .B(_20040_),
    .Y(_20041_));
 sky130_as_sc_hs__or2_2 _26538_ (.A(_19534_),
    .B(\tholin_riscv.regs[25][8] ),
    .Y(_20043_));
 sky130_as_sc_hs__or2_2 _26539_ (.A(net325),
    .B(\tholin_riscv.regs[24][8] ),
    .Y(_20044_));
 sky130_as_sc_hs__nand3_2 _26540_ (.A(net180),
    .B(_20043_),
    .C(_20044_),
    .Y(_20045_));
 sky130_as_sc_hs__or2_2 _26541_ (.A(net196),
    .B(\tholin_riscv.regs[27][8] ),
    .Y(_20046_));
 sky130_as_sc_hs__or2_2 _26542_ (.A(net325),
    .B(\tholin_riscv.regs[26][8] ),
    .Y(_20047_));
 sky130_as_sc_hs__nand3_2 _26543_ (.A(net276),
    .B(_20046_),
    .C(_20047_),
    .Y(_20048_));
 sky130_as_sc_hs__nand3_2 _26544_ (.A(net164),
    .B(_20045_),
    .C(_20048_),
    .Y(_20049_));
 sky130_as_sc_hs__or2_2 _26545_ (.A(net196),
    .B(\tholin_riscv.regs[29][8] ),
    .Y(_20050_));
 sky130_as_sc_hs__or2_2 _26546_ (.A(net326),
    .B(\tholin_riscv.regs[28][8] ),
    .Y(_20051_));
 sky130_as_sc_hs__nand3_2 _26547_ (.A(net181),
    .B(_20050_),
    .C(_20051_),
    .Y(_20052_));
 sky130_as_sc_hs__or2_2 _26548_ (.A(_19534_),
    .B(\tholin_riscv.regs[31][8] ),
    .Y(_20053_));
 sky130_as_sc_hs__or2_2 _26549_ (.A(net325),
    .B(\tholin_riscv.regs[30][8] ),
    .Y(_20054_));
 sky130_as_sc_hs__nand3_2 _26550_ (.A(net281),
    .B(_20053_),
    .C(_20054_),
    .Y(_20055_));
 sky130_as_sc_hs__nand3_2 _26551_ (.A(net260),
    .B(_20052_),
    .C(_20055_),
    .Y(_20056_));
 sky130_as_sc_hs__or2_2 _26552_ (.A(net196),
    .B(\tholin_riscv.regs[17][8] ),
    .Y(_20057_));
 sky130_as_sc_hs__or2_2 _26553_ (.A(net325),
    .B(\tholin_riscv.regs[16][8] ),
    .Y(_20058_));
 sky130_as_sc_hs__nand3_2 _26554_ (.A(net181),
    .B(_20057_),
    .C(_20058_),
    .Y(_20059_));
 sky130_as_sc_hs__or2_2 _26555_ (.A(net200),
    .B(\tholin_riscv.regs[19][8] ),
    .Y(_20060_));
 sky130_as_sc_hs__or2_2 _26556_ (.A(net330),
    .B(\tholin_riscv.regs[18][8] ),
    .Y(_20061_));
 sky130_as_sc_hs__nand3_2 _26557_ (.A(net280),
    .B(_20060_),
    .C(_20061_),
    .Y(_20062_));
 sky130_as_sc_hs__nand3_2 _26558_ (.A(net164),
    .B(_20059_),
    .C(_20062_),
    .Y(_20063_));
 sky130_as_sc_hs__or2_2 _26559_ (.A(net200),
    .B(\tholin_riscv.regs[23][8] ),
    .Y(_20064_));
 sky130_as_sc_hs__or2_2 _26560_ (.A(net330),
    .B(\tholin_riscv.regs[22][8] ),
    .Y(_20065_));
 sky130_as_sc_hs__nand3_2 _26561_ (.A(net280),
    .B(_20064_),
    .C(_20065_),
    .Y(_20066_));
 sky130_as_sc_hs__or2_2 _26562_ (.A(net200),
    .B(\tholin_riscv.regs[21][8] ),
    .Y(_20067_));
 sky130_as_sc_hs__or2_2 _26563_ (.A(net325),
    .B(\tholin_riscv.regs[20][8] ),
    .Y(_20068_));
 sky130_as_sc_hs__nand3_2 _26564_ (.A(net180),
    .B(_20067_),
    .C(_20068_),
    .Y(_20069_));
 sky130_as_sc_hs__nand3_2 _26565_ (.A(net262),
    .B(_20066_),
    .C(_20069_),
    .Y(_20070_));
 sky130_as_sc_hs__nand3_2 _26566_ (.A(net155),
    .B(_20063_),
    .C(_20070_),
    .Y(_20071_));
 sky130_as_sc_hs__nand3_2 _26567_ (.A(net252),
    .B(_20049_),
    .C(_20056_),
    .Y(_20072_));
 sky130_as_sc_hs__nand3_2 _26568_ (.A(net247),
    .B(_20071_),
    .C(_20072_),
    .Y(_20073_));
 sky130_as_sc_hs__or2_2 _26569_ (.A(net196),
    .B(\tholin_riscv.regs[9][8] ),
    .Y(_20074_));
 sky130_as_sc_hs__or2_2 _26570_ (.A(net323),
    .B(\tholin_riscv.regs[8][8] ),
    .Y(_20075_));
 sky130_as_sc_hs__nand3_2 _26571_ (.A(net182),
    .B(_20074_),
    .C(_20075_),
    .Y(_20076_));
 sky130_as_sc_hs__or2_2 _26572_ (.A(net196),
    .B(\tholin_riscv.regs[11][8] ),
    .Y(_20077_));
 sky130_as_sc_hs__or2_2 _26573_ (.A(net323),
    .B(\tholin_riscv.regs[10][8] ),
    .Y(_20078_));
 sky130_as_sc_hs__nand3_2 _26574_ (.A(net277),
    .B(_20077_),
    .C(_20078_),
    .Y(_20079_));
 sky130_as_sc_hs__nand3_2 _26575_ (.A(net163),
    .B(_20076_),
    .C(_20079_),
    .Y(_20080_));
 sky130_as_sc_hs__or2_2 _26576_ (.A(net196),
    .B(\tholin_riscv.regs[13][8] ),
    .Y(_20081_));
 sky130_as_sc_hs__or2_2 _26577_ (.A(net325),
    .B(\tholin_riscv.regs[12][8] ),
    .Y(_20082_));
 sky130_as_sc_hs__nand3_2 _26578_ (.A(net180),
    .B(_20081_),
    .C(_20082_),
    .Y(_20083_));
 sky130_as_sc_hs__or2_2 _26579_ (.A(net196),
    .B(\tholin_riscv.regs[15][8] ),
    .Y(_20084_));
 sky130_as_sc_hs__or2_2 _26580_ (.A(net325),
    .B(\tholin_riscv.regs[14][8] ),
    .Y(_20085_));
 sky130_as_sc_hs__nand3_2 _26581_ (.A(net281),
    .B(_20084_),
    .C(_20085_),
    .Y(_20086_));
 sky130_as_sc_hs__nand3_2 _26582_ (.A(net260),
    .B(_20083_),
    .C(_20086_),
    .Y(_20087_));
 sky130_as_sc_hs__or2_2 _26583_ (.A(net198),
    .B(\tholin_riscv.regs[1][8] ),
    .Y(_20088_));
 sky130_as_sc_hs__or2_2 _26584_ (.A(net323),
    .B(\tholin_riscv.regs[0][8] ),
    .Y(_20089_));
 sky130_as_sc_hs__nand3_2 _26585_ (.A(net182),
    .B(_20088_),
    .C(_20089_),
    .Y(_20090_));
 sky130_as_sc_hs__or2_2 _26586_ (.A(net196),
    .B(\tholin_riscv.regs[3][8] ),
    .Y(_20091_));
 sky130_as_sc_hs__or2_2 _26587_ (.A(net323),
    .B(\tholin_riscv.regs[2][8] ),
    .Y(_20092_));
 sky130_as_sc_hs__nand3_2 _26588_ (.A(net277),
    .B(_20091_),
    .C(_20092_),
    .Y(_20093_));
 sky130_as_sc_hs__nand3_2 _26589_ (.A(net163),
    .B(_20090_),
    .C(_20093_),
    .Y(_20094_));
 sky130_as_sc_hs__or2_2 _26590_ (.A(net198),
    .B(\tholin_riscv.regs[7][8] ),
    .Y(_20095_));
 sky130_as_sc_hs__or2_2 _26591_ (.A(net327),
    .B(\tholin_riscv.regs[6][8] ),
    .Y(_20096_));
 sky130_as_sc_hs__nand3_2 _26592_ (.A(net278),
    .B(_20095_),
    .C(_20096_),
    .Y(_20097_));
 sky130_as_sc_hs__or2_2 _26593_ (.A(net200),
    .B(\tholin_riscv.regs[5][8] ),
    .Y(_20098_));
 sky130_as_sc_hs__or2_2 _26594_ (.A(net330),
    .B(\tholin_riscv.regs[4][8] ),
    .Y(_20099_));
 sky130_as_sc_hs__nand3_2 _26595_ (.A(net185),
    .B(_20098_),
    .C(_20099_),
    .Y(_20100_));
 sky130_as_sc_hs__nand3_2 _26596_ (.A(net262),
    .B(_20097_),
    .C(_20100_),
    .Y(_20101_));
 sky130_as_sc_hs__nand3_2 _26597_ (.A(net155),
    .B(_20094_),
    .C(_20101_),
    .Y(_20102_));
 sky130_as_sc_hs__nand3_2 _26598_ (.A(net253),
    .B(_20080_),
    .C(_20087_),
    .Y(_20103_));
 sky130_as_sc_hs__nand3_2 _26599_ (.A(net150),
    .B(_20102_),
    .C(_20103_),
    .Y(_20104_));
 sky130_as_sc_hs__inv_2 _26601_ (.Y(_20106_),
    .A(_20105_));
 sky130_as_sc_hs__or2_2 _26603_ (.A(net20),
    .B(_19755_),
    .Y(_20108_));
 sky130_as_sc_hs__nand3_2 _26604_ (.A(_19759_),
    .B(_20107_),
    .C(_20108_),
    .Y(_20109_));
 sky130_as_sc_hs__or2_2 _26605_ (.A(net1710),
    .B(_20021_),
    .Y(_20110_));
 sky130_as_sc_hs__nand3_2 _26606_ (.A(_20021_),
    .B(_20042_),
    .C(_20109_),
    .Y(_20111_));
 sky130_as_sc_hs__and2_2 _26607_ (.A(net497),
    .B(_20111_),
    .Y(_20112_));
 sky130_as_sc_hs__and2_2 _26608_ (.A(_20110_),
    .B(_20112_),
    .Y(_00005_));
 sky130_as_sc_hs__nand3_2 _26618_ (.A(_20114_),
    .B(_20116_),
    .C(_20119_),
    .Y(_20122_));
 sky130_as_sc_hs__nand3_2 _26619_ (.A(_20117_),
    .B(_20118_),
    .C(_20120_),
    .Y(_20123_));
 sky130_as_sc_hs__or2_2 _26620_ (.A(_20121_),
    .B(_20123_),
    .Y(_20124_));
 sky130_as_sc_hs__nor2_2 _26621_ (.A(_20122_),
    .B(_20124_),
    .Y(_20125_));
 sky130_as_sc_hs__or2_2 _26622_ (.A(_19507_),
    .B(_20039_),
    .Y(_20126_));
 sky130_as_sc_hs__or2_2 _26625_ (.A(net193),
    .B(\tholin_riscv.regs[25][9] ),
    .Y(_20129_));
 sky130_as_sc_hs__or2_2 _26626_ (.A(net318),
    .B(\tholin_riscv.regs[24][9] ),
    .Y(_20130_));
 sky130_as_sc_hs__nand3_2 _26627_ (.A(net178),
    .B(_20129_),
    .C(_20130_),
    .Y(_20131_));
 sky130_as_sc_hs__or2_2 _26628_ (.A(net193),
    .B(\tholin_riscv.regs[27][9] ),
    .Y(_20132_));
 sky130_as_sc_hs__or2_2 _26629_ (.A(net333),
    .B(\tholin_riscv.regs[26][9] ),
    .Y(_20133_));
 sky130_as_sc_hs__nand3_2 _26630_ (.A(net271),
    .B(_20132_),
    .C(_20133_),
    .Y(_20134_));
 sky130_as_sc_hs__nand3_2 _26631_ (.A(net159),
    .B(_20131_),
    .C(_20134_),
    .Y(_20135_));
 sky130_as_sc_hs__or2_2 _26632_ (.A(net198),
    .B(\tholin_riscv.regs[29][9] ),
    .Y(_20136_));
 sky130_as_sc_hs__or2_2 _26633_ (.A(net327),
    .B(\tholin_riscv.regs[28][9] ),
    .Y(_20137_));
 sky130_as_sc_hs__nand3_2 _26634_ (.A(net183),
    .B(_20136_),
    .C(_20137_),
    .Y(_20138_));
 sky130_as_sc_hs__or2_2 _26635_ (.A(net198),
    .B(\tholin_riscv.regs[31][9] ),
    .Y(_20139_));
 sky130_as_sc_hs__or2_2 _26636_ (.A(net327),
    .B(\tholin_riscv.regs[30][9] ),
    .Y(_20140_));
 sky130_as_sc_hs__nand3_2 _26637_ (.A(net278),
    .B(_20139_),
    .C(_20140_),
    .Y(_20141_));
 sky130_as_sc_hs__nand3_2 _26638_ (.A(net261),
    .B(_20138_),
    .C(_20141_),
    .Y(_20142_));
 sky130_as_sc_hs__or2_2 _26639_ (.A(net193),
    .B(\tholin_riscv.regs[17][9] ),
    .Y(_20143_));
 sky130_as_sc_hs__or2_2 _26640_ (.A(net318),
    .B(\tholin_riscv.regs[16][9] ),
    .Y(_20144_));
 sky130_as_sc_hs__nand3_2 _26641_ (.A(net178),
    .B(_20143_),
    .C(_20144_),
    .Y(_20145_));
 sky130_as_sc_hs__or2_2 _26642_ (.A(net193),
    .B(\tholin_riscv.regs[19][9] ),
    .Y(_20146_));
 sky130_as_sc_hs__or2_2 _26643_ (.A(net320),
    .B(\tholin_riscv.regs[18][9] ),
    .Y(_20147_));
 sky130_as_sc_hs__nand3_2 _26644_ (.A(net273),
    .B(_20146_),
    .C(_20147_),
    .Y(_20148_));
 sky130_as_sc_hs__nand3_2 _26645_ (.A(net160),
    .B(_20145_),
    .C(_20148_),
    .Y(_20149_));
 sky130_as_sc_hs__or2_2 _26646_ (.A(net193),
    .B(\tholin_riscv.regs[23][9] ),
    .Y(_20150_));
 sky130_as_sc_hs__or2_2 _26647_ (.A(net319),
    .B(\tholin_riscv.regs[22][9] ),
    .Y(_20151_));
 sky130_as_sc_hs__nand3_2 _26648_ (.A(net274),
    .B(_20150_),
    .C(_20151_),
    .Y(_20152_));
 sky130_as_sc_hs__or2_2 _26649_ (.A(net198),
    .B(\tholin_riscv.regs[21][9] ),
    .Y(_20153_));
 sky130_as_sc_hs__or2_2 _26650_ (.A(net327),
    .B(\tholin_riscv.regs[20][9] ),
    .Y(_20154_));
 sky130_as_sc_hs__nand3_2 _26651_ (.A(net183),
    .B(_20153_),
    .C(_20154_),
    .Y(_20155_));
 sky130_as_sc_hs__nand3_2 _26652_ (.A(net259),
    .B(_20152_),
    .C(_20155_),
    .Y(_20156_));
 sky130_as_sc_hs__nand3_2 _26653_ (.A(net153),
    .B(_20149_),
    .C(_20156_),
    .Y(_20157_));
 sky130_as_sc_hs__nand3_2 _26654_ (.A(net250),
    .B(_20135_),
    .C(_20142_),
    .Y(_20158_));
 sky130_as_sc_hs__nand3_2 _26655_ (.A(net248),
    .B(_20157_),
    .C(_20158_),
    .Y(_20159_));
 sky130_as_sc_hs__or2_2 _26656_ (.A(net198),
    .B(\tholin_riscv.regs[9][9] ),
    .Y(_20160_));
 sky130_as_sc_hs__or2_2 _26657_ (.A(net333),
    .B(\tholin_riscv.regs[8][9] ),
    .Y(_20161_));
 sky130_as_sc_hs__nand3_2 _26658_ (.A(net182),
    .B(_20160_),
    .C(_20161_),
    .Y(_20162_));
 sky130_as_sc_hs__or2_2 _26659_ (.A(net198),
    .B(\tholin_riscv.regs[11][9] ),
    .Y(_20163_));
 sky130_as_sc_hs__or2_2 _26660_ (.A(net327),
    .B(\tholin_riscv.regs[10][9] ),
    .Y(_20164_));
 sky130_as_sc_hs__nand3_2 _26661_ (.A(net278),
    .B(_20163_),
    .C(_20164_),
    .Y(_20165_));
 sky130_as_sc_hs__nand3_2 _26662_ (.A(net163),
    .B(_20162_),
    .C(_20165_),
    .Y(_20166_));
 sky130_as_sc_hs__or2_2 _26663_ (.A(net196),
    .B(\tholin_riscv.regs[13][9] ),
    .Y(_20167_));
 sky130_as_sc_hs__or2_2 _26664_ (.A(net323),
    .B(\tholin_riscv.regs[12][9] ),
    .Y(_20168_));
 sky130_as_sc_hs__nand3_2 _26665_ (.A(net182),
    .B(_20167_),
    .C(_20168_),
    .Y(_20169_));
 sky130_as_sc_hs__or2_2 _26666_ (.A(net198),
    .B(\tholin_riscv.regs[15][9] ),
    .Y(_20170_));
 sky130_as_sc_hs__or2_2 _26667_ (.A(net323),
    .B(\tholin_riscv.regs[14][9] ),
    .Y(_20171_));
 sky130_as_sc_hs__nand3_2 _26668_ (.A(net277),
    .B(_20170_),
    .C(_20171_),
    .Y(_20172_));
 sky130_as_sc_hs__nand3_2 _26669_ (.A(net260),
    .B(_20169_),
    .C(_20172_),
    .Y(_20173_));
 sky130_as_sc_hs__or2_2 _26670_ (.A(net196),
    .B(\tholin_riscv.regs[1][9] ),
    .Y(_20174_));
 sky130_as_sc_hs__or2_2 _26671_ (.A(net323),
    .B(\tholin_riscv.regs[0][9] ),
    .Y(_20175_));
 sky130_as_sc_hs__nand3_2 _26672_ (.A(net182),
    .B(_20174_),
    .C(_20175_),
    .Y(_20176_));
 sky130_as_sc_hs__or2_2 _26673_ (.A(net196),
    .B(\tholin_riscv.regs[3][9] ),
    .Y(_20177_));
 sky130_as_sc_hs__or2_2 _26674_ (.A(net323),
    .B(\tholin_riscv.regs[2][9] ),
    .Y(_20178_));
 sky130_as_sc_hs__nand3_2 _26675_ (.A(net277),
    .B(_20177_),
    .C(_20178_),
    .Y(_20179_));
 sky130_as_sc_hs__nand3_2 _26676_ (.A(net163),
    .B(_20176_),
    .C(_20179_),
    .Y(_20180_));
 sky130_as_sc_hs__or2_2 _26677_ (.A(net196),
    .B(\tholin_riscv.regs[7][9] ),
    .Y(_20181_));
 sky130_as_sc_hs__or2_2 _26678_ (.A(net323),
    .B(\tholin_riscv.regs[6][9] ),
    .Y(_20182_));
 sky130_as_sc_hs__nand3_2 _26679_ (.A(net277),
    .B(_20181_),
    .C(_20182_),
    .Y(_20183_));
 sky130_as_sc_hs__or2_2 _26680_ (.A(net196),
    .B(\tholin_riscv.regs[5][9] ),
    .Y(_20184_));
 sky130_as_sc_hs__or2_2 _26681_ (.A(net323),
    .B(\tholin_riscv.regs[4][9] ),
    .Y(_20185_));
 sky130_as_sc_hs__nand3_2 _26682_ (.A(net182),
    .B(_20184_),
    .C(_20185_),
    .Y(_20186_));
 sky130_as_sc_hs__nand3_2 _26683_ (.A(net260),
    .B(_20183_),
    .C(_20186_),
    .Y(_20187_));
 sky130_as_sc_hs__nand3_2 _26684_ (.A(net155),
    .B(_20180_),
    .C(_20187_),
    .Y(_20188_));
 sky130_as_sc_hs__nand3_2 _26685_ (.A(net252),
    .B(_20166_),
    .C(_20173_),
    .Y(_20189_));
 sky130_as_sc_hs__nand3_2 _26686_ (.A(_19538_),
    .B(_20188_),
    .C(_20189_),
    .Y(_20190_));
 sky130_as_sc_hs__inv_2 _26688_ (.Y(_20192_),
    .A(_20191_));
 sky130_as_sc_hs__or2_2 _26690_ (.A(net21),
    .B(_19755_),
    .Y(_20194_));
 sky130_as_sc_hs__nand3_2 _26691_ (.A(_19759_),
    .B(_20193_),
    .C(_20194_),
    .Y(_20195_));
 sky130_as_sc_hs__or2_2 _26692_ (.A(net1780),
    .B(_20021_),
    .Y(_20196_));
 sky130_as_sc_hs__nand3_2 _26693_ (.A(_20021_),
    .B(_20128_),
    .C(_20195_),
    .Y(_20197_));
 sky130_as_sc_hs__and2_2 _26694_ (.A(net497),
    .B(_20197_),
    .Y(_20198_));
 sky130_as_sc_hs__and2_2 _26695_ (.A(_20196_),
    .B(_20198_),
    .Y(_00006_));
 sky130_as_sc_hs__nand3_2 _26705_ (.A(_20200_),
    .B(_20202_),
    .C(_20205_),
    .Y(_20208_));
 sky130_as_sc_hs__nand3_2 _26706_ (.A(_20203_),
    .B(_20204_),
    .C(_20206_),
    .Y(_20209_));
 sky130_as_sc_hs__or2_2 _26707_ (.A(_20207_),
    .B(_20209_),
    .Y(_20210_));
 sky130_as_sc_hs__nor2_2 _26708_ (.A(_20208_),
    .B(_20210_),
    .Y(_20211_));
 sky130_as_sc_hs__or2_2 _26709_ (.A(_19506_),
    .B(_20039_),
    .Y(_20212_));
 sky130_as_sc_hs__or2_2 _26712_ (.A(net193),
    .B(\tholin_riscv.regs[25][10] ),
    .Y(_20215_));
 sky130_as_sc_hs__or2_2 _26713_ (.A(net318),
    .B(\tholin_riscv.regs[24][10] ),
    .Y(_20216_));
 sky130_as_sc_hs__nand3_2 _26714_ (.A(net178),
    .B(_20215_),
    .C(_20216_),
    .Y(_20217_));
 sky130_as_sc_hs__or2_2 _26715_ (.A(net193),
    .B(\tholin_riscv.regs[27][10] ),
    .Y(_20218_));
 sky130_as_sc_hs__or2_2 _26716_ (.A(net319),
    .B(\tholin_riscv.regs[26][10] ),
    .Y(_20219_));
 sky130_as_sc_hs__nand3_2 _26717_ (.A(net274),
    .B(_20218_),
    .C(_20219_),
    .Y(_20220_));
 sky130_as_sc_hs__nand3_2 _26718_ (.A(net159),
    .B(_20217_),
    .C(_20220_),
    .Y(_20221_));
 sky130_as_sc_hs__or2_2 _26719_ (.A(net193),
    .B(\tholin_riscv.regs[29][10] ),
    .Y(_20222_));
 sky130_as_sc_hs__or2_2 _26720_ (.A(net318),
    .B(\tholin_riscv.regs[28][10] ),
    .Y(_20223_));
 sky130_as_sc_hs__nand3_2 _26721_ (.A(net178),
    .B(_20222_),
    .C(_20223_),
    .Y(_20224_));
 sky130_as_sc_hs__or2_2 _26722_ (.A(net193),
    .B(\tholin_riscv.regs[31][10] ),
    .Y(_20225_));
 sky130_as_sc_hs__or2_2 _26723_ (.A(net319),
    .B(\tholin_riscv.regs[30][10] ),
    .Y(_20226_));
 sky130_as_sc_hs__nand3_2 _26724_ (.A(net274),
    .B(_20225_),
    .C(_20226_),
    .Y(_20227_));
 sky130_as_sc_hs__nand3_2 _26725_ (.A(net259),
    .B(_20224_),
    .C(_20227_),
    .Y(_20228_));
 sky130_as_sc_hs__or2_2 _26726_ (.A(net193),
    .B(\tholin_riscv.regs[17][10] ),
    .Y(_20229_));
 sky130_as_sc_hs__or2_2 _26727_ (.A(net318),
    .B(\tholin_riscv.regs[16][10] ),
    .Y(_20230_));
 sky130_as_sc_hs__nand3_2 _26728_ (.A(net178),
    .B(_20229_),
    .C(_20230_),
    .Y(_20231_));
 sky130_as_sc_hs__or2_2 _26729_ (.A(net193),
    .B(\tholin_riscv.regs[19][10] ),
    .Y(_20232_));
 sky130_as_sc_hs__or2_2 _26730_ (.A(net318),
    .B(\tholin_riscv.regs[18][10] ),
    .Y(_20233_));
 sky130_as_sc_hs__nand3_2 _26731_ (.A(net274),
    .B(_20232_),
    .C(_20233_),
    .Y(_20234_));
 sky130_as_sc_hs__nand3_2 _26732_ (.A(net159),
    .B(_20231_),
    .C(_20234_),
    .Y(_20235_));
 sky130_as_sc_hs__or2_2 _26733_ (.A(net188),
    .B(\tholin_riscv.regs[23][10] ),
    .Y(_20236_));
 sky130_as_sc_hs__or2_2 _26734_ (.A(net313),
    .B(\tholin_riscv.regs[22][10] ),
    .Y(_20237_));
 sky130_as_sc_hs__nand3_2 _26735_ (.A(net271),
    .B(_20236_),
    .C(_20237_),
    .Y(_20238_));
 sky130_as_sc_hs__or2_2 _26736_ (.A(net188),
    .B(\tholin_riscv.regs[21][10] ),
    .Y(_20239_));
 sky130_as_sc_hs__or2_2 _26737_ (.A(net333),
    .B(\tholin_riscv.regs[20][10] ),
    .Y(_20240_));
 sky130_as_sc_hs__nand3_2 _26738_ (.A(net175),
    .B(_20239_),
    .C(_20240_),
    .Y(_20241_));
 sky130_as_sc_hs__nand3_2 _26739_ (.A(net259),
    .B(_20238_),
    .C(_20241_),
    .Y(_20242_));
 sky130_as_sc_hs__nand3_2 _26740_ (.A(net152),
    .B(_20235_),
    .C(_20242_),
    .Y(_20243_));
 sky130_as_sc_hs__nand3_2 _26741_ (.A(net249),
    .B(_20221_),
    .C(_20228_),
    .Y(_20244_));
 sky130_as_sc_hs__nand3_2 _26742_ (.A(net248),
    .B(_20243_),
    .C(_20244_),
    .Y(_20245_));
 sky130_as_sc_hs__or2_2 _26743_ (.A(net189),
    .B(\tholin_riscv.regs[9][10] ),
    .Y(_20246_));
 sky130_as_sc_hs__or2_2 _26744_ (.A(net313),
    .B(\tholin_riscv.regs[8][10] ),
    .Y(_20247_));
 sky130_as_sc_hs__nand3_2 _26745_ (.A(net175),
    .B(_20246_),
    .C(_20247_),
    .Y(_20248_));
 sky130_as_sc_hs__or2_2 _26746_ (.A(net189),
    .B(\tholin_riscv.regs[11][10] ),
    .Y(_20249_));
 sky130_as_sc_hs__or2_2 _26747_ (.A(net313),
    .B(\tholin_riscv.regs[10][10] ),
    .Y(_20250_));
 sky130_as_sc_hs__nand3_2 _26748_ (.A(net271),
    .B(_20249_),
    .C(_20250_),
    .Y(_20251_));
 sky130_as_sc_hs__nand3_2 _26749_ (.A(net159),
    .B(_20248_),
    .C(_20251_),
    .Y(_20252_));
 sky130_as_sc_hs__or2_2 _26750_ (.A(net189),
    .B(\tholin_riscv.regs[13][10] ),
    .Y(_20253_));
 sky130_as_sc_hs__or2_2 _26751_ (.A(net313),
    .B(\tholin_riscv.regs[12][10] ),
    .Y(_20254_));
 sky130_as_sc_hs__nand3_2 _26752_ (.A(net175),
    .B(_20253_),
    .C(_20254_),
    .Y(_20255_));
 sky130_as_sc_hs__or2_2 _26753_ (.A(net188),
    .B(\tholin_riscv.regs[15][10] ),
    .Y(_20256_));
 sky130_as_sc_hs__or2_2 _26754_ (.A(net313),
    .B(\tholin_riscv.regs[14][10] ),
    .Y(_20257_));
 sky130_as_sc_hs__nand3_2 _26755_ (.A(net271),
    .B(_20256_),
    .C(_20257_),
    .Y(_20258_));
 sky130_as_sc_hs__nand3_2 _26756_ (.A(net257),
    .B(_20255_),
    .C(_20258_),
    .Y(_20259_));
 sky130_as_sc_hs__or2_2 _26757_ (.A(net188),
    .B(\tholin_riscv.regs[1][10] ),
    .Y(_20260_));
 sky130_as_sc_hs__or2_2 _26758_ (.A(net312),
    .B(\tholin_riscv.regs[0][10] ),
    .Y(_20261_));
 sky130_as_sc_hs__nand3_2 _26759_ (.A(net175),
    .B(_20260_),
    .C(_20261_),
    .Y(_20262_));
 sky130_as_sc_hs__or2_2 _26760_ (.A(net188),
    .B(\tholin_riscv.regs[3][10] ),
    .Y(_20263_));
 sky130_as_sc_hs__or2_2 _26761_ (.A(net313),
    .B(\tholin_riscv.regs[2][10] ),
    .Y(_20264_));
 sky130_as_sc_hs__nand3_2 _26762_ (.A(net271),
    .B(_20263_),
    .C(_20264_),
    .Y(_20265_));
 sky130_as_sc_hs__nand3_2 _26763_ (.A(net159),
    .B(_20262_),
    .C(_20265_),
    .Y(_20266_));
 sky130_as_sc_hs__or2_2 _26764_ (.A(net189),
    .B(\tholin_riscv.regs[7][10] ),
    .Y(_20267_));
 sky130_as_sc_hs__or2_2 _26765_ (.A(net313),
    .B(\tholin_riscv.regs[6][10] ),
    .Y(_20268_));
 sky130_as_sc_hs__nand3_2 _26766_ (.A(net271),
    .B(_20267_),
    .C(_20268_),
    .Y(_20269_));
 sky130_as_sc_hs__or2_2 _26767_ (.A(net196),
    .B(\tholin_riscv.regs[5][10] ),
    .Y(_20270_));
 sky130_as_sc_hs__or2_2 _26768_ (.A(net313),
    .B(\tholin_riscv.regs[4][10] ),
    .Y(_20271_));
 sky130_as_sc_hs__nand3_2 _26769_ (.A(net175),
    .B(_20270_),
    .C(_20271_),
    .Y(_20272_));
 sky130_as_sc_hs__nand3_2 _26770_ (.A(net257),
    .B(_20269_),
    .C(_20272_),
    .Y(_20273_));
 sky130_as_sc_hs__nand3_2 _26771_ (.A(net152),
    .B(_20266_),
    .C(_20273_),
    .Y(_20274_));
 sky130_as_sc_hs__nand3_2 _26772_ (.A(net249),
    .B(_20252_),
    .C(_20259_),
    .Y(_20275_));
 sky130_as_sc_hs__nand3_2 _26773_ (.A(net150),
    .B(_20274_),
    .C(_20275_),
    .Y(_20276_));
 sky130_as_sc_hs__or2_2 _26776_ (.A(net4),
    .B(_19755_),
    .Y(_20279_));
 sky130_as_sc_hs__nand3_2 _26777_ (.A(_19759_),
    .B(_20278_),
    .C(_20279_),
    .Y(_20280_));
 sky130_as_sc_hs__or2_2 _26778_ (.A(net1791),
    .B(_20021_),
    .Y(_20281_));
 sky130_as_sc_hs__nand3_2 _26779_ (.A(_20021_),
    .B(_20214_),
    .C(_20280_),
    .Y(_20282_));
 sky130_as_sc_hs__and2_2 _26780_ (.A(net497),
    .B(_20282_),
    .Y(_20283_));
 sky130_as_sc_hs__and2_2 _26781_ (.A(_20281_),
    .B(_20283_),
    .Y(_00007_));
 sky130_as_sc_hs__and2_2 _26786_ (.A(_20286_),
    .B(_20287_),
    .Y(_20288_));
 sky130_as_sc_hs__nand3_2 _26787_ (.A(_20284_),
    .B(_20285_),
    .C(_20288_),
    .Y(_20289_));
 sky130_as_sc_hs__nand3_2 _26793_ (.A(_19993_),
    .B(_20293_),
    .C(_20294_),
    .Y(_20295_));
 sky130_as_sc_hs__or2_2 _26794_ (.A(_20292_),
    .B(_20295_),
    .Y(_20296_));
 sky130_as_sc_hs__nor2_2 _26795_ (.A(_20289_),
    .B(_20296_),
    .Y(_20297_));
 sky130_as_sc_hs__or2_2 _26796_ (.A(\tholin_riscv.uart.divisor[11] ),
    .B(_20039_),
    .Y(_20298_));
 sky130_as_sc_hs__nand3_2 _26798_ (.A(net137),
    .B(_20298_),
    .C(_20299_),
    .Y(_20300_));
 sky130_as_sc_hs__or2_2 _26799_ (.A(net190),
    .B(\tholin_riscv.regs[25][11] ),
    .Y(_20301_));
 sky130_as_sc_hs__or2_2 _26800_ (.A(net310),
    .B(\tholin_riscv.regs[24][11] ),
    .Y(_20302_));
 sky130_as_sc_hs__nand3_2 _26801_ (.A(net174),
    .B(_20301_),
    .C(_20302_),
    .Y(_20303_));
 sky130_as_sc_hs__or2_2 _26802_ (.A(net190),
    .B(\tholin_riscv.regs[27][11] ),
    .Y(_20304_));
 sky130_as_sc_hs__or2_2 _26803_ (.A(net309),
    .B(\tholin_riscv.regs[26][11] ),
    .Y(_20305_));
 sky130_as_sc_hs__nand3_2 _26804_ (.A(net270),
    .B(_20304_),
    .C(_20305_),
    .Y(_20306_));
 sky130_as_sc_hs__nand3_2 _26805_ (.A(net158),
    .B(_20303_),
    .C(_20306_),
    .Y(_20307_));
 sky130_as_sc_hs__or2_2 _26806_ (.A(net187),
    .B(\tholin_riscv.regs[29][11] ),
    .Y(_20308_));
 sky130_as_sc_hs__or2_2 _26807_ (.A(net310),
    .B(\tholin_riscv.regs[28][11] ),
    .Y(_20309_));
 sky130_as_sc_hs__nand3_2 _26808_ (.A(net174),
    .B(_20308_),
    .C(_20309_),
    .Y(_20310_));
 sky130_as_sc_hs__or2_2 _26809_ (.A(net195),
    .B(\tholin_riscv.regs[31][11] ),
    .Y(_20311_));
 sky130_as_sc_hs__or2_2 _26810_ (.A(net310),
    .B(\tholin_riscv.regs[30][11] ),
    .Y(_20312_));
 sky130_as_sc_hs__nand3_2 _26811_ (.A(net270),
    .B(_20311_),
    .C(_20312_),
    .Y(_20313_));
 sky130_as_sc_hs__nand3_2 _26812_ (.A(net257),
    .B(_20310_),
    .C(_20313_),
    .Y(_20314_));
 sky130_as_sc_hs__or2_2 _26813_ (.A(net187),
    .B(\tholin_riscv.regs[17][11] ),
    .Y(_20315_));
 sky130_as_sc_hs__or2_2 _26814_ (.A(net308),
    .B(\tholin_riscv.regs[16][11] ),
    .Y(_20316_));
 sky130_as_sc_hs__nand3_2 _26815_ (.A(net174),
    .B(_20315_),
    .C(_20316_),
    .Y(_20317_));
 sky130_as_sc_hs__or2_2 _26816_ (.A(net190),
    .B(\tholin_riscv.regs[19][11] ),
    .Y(_20318_));
 sky130_as_sc_hs__or2_2 _26817_ (.A(net310),
    .B(\tholin_riscv.regs[18][11] ),
    .Y(_20319_));
 sky130_as_sc_hs__nand3_2 _26818_ (.A(net270),
    .B(_20318_),
    .C(_20319_),
    .Y(_20320_));
 sky130_as_sc_hs__nand3_2 _26819_ (.A(net158),
    .B(_20317_),
    .C(_20320_),
    .Y(_20321_));
 sky130_as_sc_hs__or2_2 _26820_ (.A(net187),
    .B(\tholin_riscv.regs[23][11] ),
    .Y(_20322_));
 sky130_as_sc_hs__or2_2 _26821_ (.A(net308),
    .B(\tholin_riscv.regs[22][11] ),
    .Y(_20323_));
 sky130_as_sc_hs__nand3_2 _26822_ (.A(net270),
    .B(_20322_),
    .C(_20323_),
    .Y(_20324_));
 sky130_as_sc_hs__or2_2 _26823_ (.A(net187),
    .B(\tholin_riscv.regs[21][11] ),
    .Y(_20325_));
 sky130_as_sc_hs__or2_2 _26824_ (.A(net310),
    .B(\tholin_riscv.regs[20][11] ),
    .Y(_20326_));
 sky130_as_sc_hs__nand3_2 _26825_ (.A(net174),
    .B(_20325_),
    .C(_20326_),
    .Y(_20327_));
 sky130_as_sc_hs__nand3_2 _26826_ (.A(net257),
    .B(_20324_),
    .C(_20327_),
    .Y(_20328_));
 sky130_as_sc_hs__nand3_2 _26827_ (.A(net152),
    .B(_20321_),
    .C(_20328_),
    .Y(_20329_));
 sky130_as_sc_hs__nand3_2 _26828_ (.A(net249),
    .B(_20307_),
    .C(_20314_),
    .Y(_20330_));
 sky130_as_sc_hs__nand3_2 _26829_ (.A(net248),
    .B(_20329_),
    .C(_20330_),
    .Y(_20331_));
 sky130_as_sc_hs__or2_2 _26830_ (.A(net189),
    .B(\tholin_riscv.regs[9][11] ),
    .Y(_20332_));
 sky130_as_sc_hs__or2_2 _26831_ (.A(net313),
    .B(\tholin_riscv.regs[8][11] ),
    .Y(_20333_));
 sky130_as_sc_hs__nand3_2 _26832_ (.A(net175),
    .B(_20332_),
    .C(_20333_),
    .Y(_20334_));
 sky130_as_sc_hs__or2_2 _26833_ (.A(net193),
    .B(\tholin_riscv.regs[11][11] ),
    .Y(_20335_));
 sky130_as_sc_hs__or2_2 _26834_ (.A(net313),
    .B(\tholin_riscv.regs[10][11] ),
    .Y(_20336_));
 sky130_as_sc_hs__nand3_2 _26835_ (.A(net271),
    .B(_20335_),
    .C(_20336_),
    .Y(_20337_));
 sky130_as_sc_hs__nand3_2 _26836_ (.A(net159),
    .B(_20334_),
    .C(_20337_),
    .Y(_20338_));
 sky130_as_sc_hs__or2_2 _26837_ (.A(net188),
    .B(\tholin_riscv.regs[13][11] ),
    .Y(_20339_));
 sky130_as_sc_hs__or2_2 _26838_ (.A(net313),
    .B(\tholin_riscv.regs[12][11] ),
    .Y(_20340_));
 sky130_as_sc_hs__nand3_2 _26839_ (.A(net175),
    .B(_20339_),
    .C(_20340_),
    .Y(_20341_));
 sky130_as_sc_hs__or2_2 _26840_ (.A(net189),
    .B(\tholin_riscv.regs[15][11] ),
    .Y(_20342_));
 sky130_as_sc_hs__or2_2 _26841_ (.A(net313),
    .B(\tholin_riscv.regs[14][11] ),
    .Y(_20343_));
 sky130_as_sc_hs__nand3_2 _26842_ (.A(net271),
    .B(_20342_),
    .C(_20343_),
    .Y(_20344_));
 sky130_as_sc_hs__nand3_2 _26843_ (.A(net257),
    .B(_20341_),
    .C(_20344_),
    .Y(_20345_));
 sky130_as_sc_hs__or2_2 _26844_ (.A(net189),
    .B(\tholin_riscv.regs[1][11] ),
    .Y(_20346_));
 sky130_as_sc_hs__or2_2 _26845_ (.A(net310),
    .B(\tholin_riscv.regs[0][11] ),
    .Y(_20347_));
 sky130_as_sc_hs__nand3_2 _26846_ (.A(net174),
    .B(_20346_),
    .C(_20347_),
    .Y(_20348_));
 sky130_as_sc_hs__or2_2 _26847_ (.A(net190),
    .B(\tholin_riscv.regs[3][11] ),
    .Y(_20349_));
 sky130_as_sc_hs__or2_2 _26848_ (.A(net310),
    .B(\tholin_riscv.regs[2][11] ),
    .Y(_20350_));
 sky130_as_sc_hs__nand3_2 _26849_ (.A(net270),
    .B(_20349_),
    .C(_20350_),
    .Y(_20351_));
 sky130_as_sc_hs__nand3_2 _26850_ (.A(net158),
    .B(_20348_),
    .C(_20351_),
    .Y(_20352_));
 sky130_as_sc_hs__or2_2 _26851_ (.A(net190),
    .B(\tholin_riscv.regs[7][11] ),
    .Y(_20353_));
 sky130_as_sc_hs__or2_2 _26852_ (.A(net310),
    .B(\tholin_riscv.regs[6][11] ),
    .Y(_20354_));
 sky130_as_sc_hs__nand3_2 _26853_ (.A(net270),
    .B(_20353_),
    .C(_20354_),
    .Y(_20355_));
 sky130_as_sc_hs__or2_2 _26854_ (.A(net187),
    .B(\tholin_riscv.regs[5][11] ),
    .Y(_20356_));
 sky130_as_sc_hs__or2_2 _26855_ (.A(net310),
    .B(\tholin_riscv.regs[4][11] ),
    .Y(_20357_));
 sky130_as_sc_hs__nand3_2 _26856_ (.A(net174),
    .B(_20356_),
    .C(_20357_),
    .Y(_20358_));
 sky130_as_sc_hs__nand3_2 _26857_ (.A(net257),
    .B(_20355_),
    .C(_20358_),
    .Y(_20359_));
 sky130_as_sc_hs__nand3_2 _26858_ (.A(net152),
    .B(_20352_),
    .C(_20359_),
    .Y(_20360_));
 sky130_as_sc_hs__nand3_2 _26859_ (.A(net249),
    .B(_20338_),
    .C(_20345_),
    .Y(_20361_));
 sky130_as_sc_hs__nand3_2 _26860_ (.A(net150),
    .B(_20360_),
    .C(_20361_),
    .Y(_20362_));
 sky130_as_sc_hs__inv_2 _26862_ (.Y(_20364_),
    .A(_20363_));
 sky130_as_sc_hs__or2_2 _26864_ (.A(net5),
    .B(_19755_),
    .Y(_20366_));
 sky130_as_sc_hs__nand3_2 _26865_ (.A(_19759_),
    .B(_20365_),
    .C(_20366_),
    .Y(_20367_));
 sky130_as_sc_hs__or2_2 _26866_ (.A(net1792),
    .B(_20021_),
    .Y(_20368_));
 sky130_as_sc_hs__nand3_2 _26867_ (.A(_20021_),
    .B(_20300_),
    .C(_20367_),
    .Y(_20369_));
 sky130_as_sc_hs__and2_2 _26868_ (.A(net502),
    .B(_20369_),
    .Y(_20370_));
 sky130_as_sc_hs__and2_2 _26869_ (.A(_20368_),
    .B(_20370_),
    .Y(_00008_));
 sky130_as_sc_hs__nand3_2 _26879_ (.A(_20372_),
    .B(_20374_),
    .C(_20377_),
    .Y(_20380_));
 sky130_as_sc_hs__nand3_2 _26880_ (.A(_20375_),
    .B(_20376_),
    .C(_20378_),
    .Y(_20381_));
 sky130_as_sc_hs__or2_2 _26881_ (.A(_20379_),
    .B(_20381_),
    .Y(_20382_));
 sky130_as_sc_hs__nor2_2 _26882_ (.A(_20380_),
    .B(_20382_),
    .Y(_20383_));
 sky130_as_sc_hs__or2_2 _26883_ (.A(_19505_),
    .B(_20039_),
    .Y(_20384_));
 sky130_as_sc_hs__nand2b_2 _26886_ (.B(net314),
    .Y(_20387_),
    .A(\tholin_riscv.regs[25][12] ));
 sky130_as_sc_hs__or2_2 _26887_ (.A(net314),
    .B(\tholin_riscv.regs[24][12] ),
    .Y(_20388_));
 sky130_as_sc_hs__nand3_2 _26888_ (.A(net176),
    .B(_20387_),
    .C(_20388_),
    .Y(_20389_));
 sky130_as_sc_hs__nand2b_2 _26889_ (.B(net314),
    .Y(_20390_),
    .A(\tholin_riscv.regs[27][12] ));
 sky130_as_sc_hs__or2_2 _26890_ (.A(net314),
    .B(\tholin_riscv.regs[26][12] ),
    .Y(_20391_));
 sky130_as_sc_hs__nand3_2 _26891_ (.A(net272),
    .B(_20390_),
    .C(_20391_),
    .Y(_20392_));
 sky130_as_sc_hs__nand3_2 _26892_ (.A(net160),
    .B(_20389_),
    .C(_20392_),
    .Y(_20393_));
 sky130_as_sc_hs__nand2b_2 _26893_ (.B(net314),
    .Y(_20394_),
    .A(\tholin_riscv.regs[29][12] ));
 sky130_as_sc_hs__or2_2 _26894_ (.A(net314),
    .B(\tholin_riscv.regs[28][12] ),
    .Y(_20395_));
 sky130_as_sc_hs__nand3_2 _26895_ (.A(net176),
    .B(_20394_),
    .C(_20395_),
    .Y(_20396_));
 sky130_as_sc_hs__nand2b_2 _26896_ (.B(net314),
    .Y(_20397_),
    .A(\tholin_riscv.regs[31][12] ));
 sky130_as_sc_hs__or2_2 _26897_ (.A(net314),
    .B(\tholin_riscv.regs[30][12] ),
    .Y(_20398_));
 sky130_as_sc_hs__nand3_2 _26898_ (.A(net272),
    .B(_20397_),
    .C(_20398_),
    .Y(_20399_));
 sky130_as_sc_hs__nand3_2 _26899_ (.A(net258),
    .B(_20396_),
    .C(_20399_),
    .Y(_20400_));
 sky130_as_sc_hs__nand2b_2 _26900_ (.B(net309),
    .Y(_20401_),
    .A(\tholin_riscv.regs[17][12] ));
 sky130_as_sc_hs__or2_2 _26901_ (.A(net310),
    .B(\tholin_riscv.regs[16][12] ),
    .Y(_20402_));
 sky130_as_sc_hs__nand3_2 _26902_ (.A(net174),
    .B(_20401_),
    .C(_20402_),
    .Y(_20403_));
 sky130_as_sc_hs__nand2b_2 _26903_ (.B(net309),
    .Y(_20404_),
    .A(\tholin_riscv.regs[19][12] ));
 sky130_as_sc_hs__or2_2 _26904_ (.A(net309),
    .B(\tholin_riscv.regs[18][12] ),
    .Y(_20405_));
 sky130_as_sc_hs__nand3_2 _26905_ (.A(net270),
    .B(_20404_),
    .C(_20405_),
    .Y(_20406_));
 sky130_as_sc_hs__nand3_2 _26906_ (.A(net158),
    .B(_20403_),
    .C(_20406_),
    .Y(_20407_));
 sky130_as_sc_hs__nand2b_2 _26907_ (.B(net309),
    .Y(_20408_),
    .A(\tholin_riscv.regs[23][12] ));
 sky130_as_sc_hs__or2_2 _26908_ (.A(net309),
    .B(\tholin_riscv.regs[22][12] ),
    .Y(_20409_));
 sky130_as_sc_hs__nand3_2 _26909_ (.A(net270),
    .B(_20408_),
    .C(_20409_),
    .Y(_20410_));
 sky130_as_sc_hs__nand2b_2 _26910_ (.B(net309),
    .Y(_20411_),
    .A(\tholin_riscv.regs[21][12] ));
 sky130_as_sc_hs__or2_2 _26911_ (.A(net309),
    .B(\tholin_riscv.regs[20][12] ),
    .Y(_20412_));
 sky130_as_sc_hs__nand3_2 _26912_ (.A(net174),
    .B(_20411_),
    .C(_20412_),
    .Y(_20413_));
 sky130_as_sc_hs__nand3_2 _26913_ (.A(net257),
    .B(_20410_),
    .C(_20413_),
    .Y(_20414_));
 sky130_as_sc_hs__nand3_2 _26914_ (.A(net152),
    .B(_20407_),
    .C(_20414_),
    .Y(_20415_));
 sky130_as_sc_hs__nand3_2 _26915_ (.A(net249),
    .B(_20393_),
    .C(_20400_),
    .Y(_20416_));
 sky130_as_sc_hs__nand3_2 _26916_ (.A(net248),
    .B(_20415_),
    .C(_20416_),
    .Y(_20417_));
 sky130_as_sc_hs__nand2b_2 _26917_ (.B(net318),
    .Y(_20418_),
    .A(\tholin_riscv.regs[9][12] ));
 sky130_as_sc_hs__or2_2 _26918_ (.A(net318),
    .B(\tholin_riscv.regs[8][12] ),
    .Y(_20419_));
 sky130_as_sc_hs__nand3_2 _26919_ (.A(net178),
    .B(_20418_),
    .C(_20419_),
    .Y(_20420_));
 sky130_as_sc_hs__nand2b_2 _26920_ (.B(net318),
    .Y(_20421_),
    .A(\tholin_riscv.regs[11][12] ));
 sky130_as_sc_hs__or2_2 _26921_ (.A(net318),
    .B(\tholin_riscv.regs[10][12] ),
    .Y(_20422_));
 sky130_as_sc_hs__nand3_2 _26922_ (.A(net274),
    .B(_20421_),
    .C(_20422_),
    .Y(_20423_));
 sky130_as_sc_hs__nand3_2 _26923_ (.A(net160),
    .B(_20420_),
    .C(_20423_),
    .Y(_20424_));
 sky130_as_sc_hs__nand2b_2 _26924_ (.B(net318),
    .Y(_20425_),
    .A(\tholin_riscv.regs[13][12] ));
 sky130_as_sc_hs__or2_2 _26925_ (.A(net315),
    .B(\tholin_riscv.regs[12][12] ),
    .Y(_20426_));
 sky130_as_sc_hs__nand3_2 _26926_ (.A(net176),
    .B(_20425_),
    .C(_20426_),
    .Y(_20427_));
 sky130_as_sc_hs__nand2b_2 _26927_ (.B(net315),
    .Y(_20428_),
    .A(\tholin_riscv.regs[15][12] ));
 sky130_as_sc_hs__or2_2 _26928_ (.A(net315),
    .B(\tholin_riscv.regs[14][12] ),
    .Y(_20429_));
 sky130_as_sc_hs__nand3_2 _26929_ (.A(net272),
    .B(_20428_),
    .C(_20429_),
    .Y(_20430_));
 sky130_as_sc_hs__nand3_2 _26930_ (.A(net258),
    .B(_20427_),
    .C(_20430_),
    .Y(_20431_));
 sky130_as_sc_hs__nand2b_2 _26931_ (.B(net319),
    .Y(_20432_),
    .A(\tholin_riscv.regs[1][12] ));
 sky130_as_sc_hs__or2_2 _26932_ (.A(net319),
    .B(\tholin_riscv.regs[0][12] ),
    .Y(_20433_));
 sky130_as_sc_hs__nand3_2 _26933_ (.A(net177),
    .B(_20432_),
    .C(_20433_),
    .Y(_20434_));
 sky130_as_sc_hs__nand2b_2 _26934_ (.B(net320),
    .Y(_20435_),
    .A(\tholin_riscv.regs[3][12] ));
 sky130_as_sc_hs__or2_2 _26935_ (.A(net318),
    .B(\tholin_riscv.regs[2][12] ),
    .Y(_20436_));
 sky130_as_sc_hs__nand3_2 _26936_ (.A(net273),
    .B(_20435_),
    .C(_20436_),
    .Y(_20437_));
 sky130_as_sc_hs__nand3_2 _26937_ (.A(net159),
    .B(_20434_),
    .C(_20437_),
    .Y(_20438_));
 sky130_as_sc_hs__nand2b_2 _26938_ (.B(net318),
    .Y(_20439_),
    .A(\tholin_riscv.regs[7][12] ));
 sky130_as_sc_hs__or2_2 _26939_ (.A(net318),
    .B(\tholin_riscv.regs[6][12] ),
    .Y(_20440_));
 sky130_as_sc_hs__nand3_2 _26940_ (.A(net274),
    .B(_20439_),
    .C(_20440_),
    .Y(_20441_));
 sky130_as_sc_hs__nand2b_2 _26941_ (.B(net318),
    .Y(_20442_),
    .A(\tholin_riscv.regs[5][12] ));
 sky130_as_sc_hs__or2_2 _26942_ (.A(net318),
    .B(\tholin_riscv.regs[4][12] ),
    .Y(_20443_));
 sky130_as_sc_hs__nand3_2 _26943_ (.A(net177),
    .B(_20442_),
    .C(_20443_),
    .Y(_20444_));
 sky130_as_sc_hs__nand3_2 _26944_ (.A(net258),
    .B(_20441_),
    .C(_20444_),
    .Y(_20445_));
 sky130_as_sc_hs__nand3_2 _26945_ (.A(net152),
    .B(_20438_),
    .C(_20445_),
    .Y(_20446_));
 sky130_as_sc_hs__nand3_2 _26946_ (.A(net250),
    .B(_20424_),
    .C(_20431_),
    .Y(_20447_));
 sky130_as_sc_hs__nand3_2 _26947_ (.A(net150),
    .B(_20446_),
    .C(_20447_),
    .Y(_20448_));
 sky130_as_sc_hs__or2_2 _26950_ (.A(net6),
    .B(_19755_),
    .Y(_20451_));
 sky130_as_sc_hs__nand3_2 _26951_ (.A(_19759_),
    .B(_20450_),
    .C(_20451_),
    .Y(_20452_));
 sky130_as_sc_hs__or2_2 _26952_ (.A(net1678),
    .B(_20021_),
    .Y(_20453_));
 sky130_as_sc_hs__nand3_2 _26953_ (.A(_20021_),
    .B(_20386_),
    .C(_20452_),
    .Y(_20454_));
 sky130_as_sc_hs__and2_2 _26954_ (.A(net497),
    .B(_20454_),
    .Y(_20455_));
 sky130_as_sc_hs__and2_2 _26955_ (.A(_20453_),
    .B(_20455_),
    .Y(_00009_));
 sky130_as_sc_hs__and2_2 _26960_ (.A(_20458_),
    .B(_20459_),
    .Y(_20460_));
 sky130_as_sc_hs__nand3_2 _26961_ (.A(_20456_),
    .B(_20457_),
    .C(_20460_),
    .Y(_20461_));
 sky130_as_sc_hs__nand3_2 _26967_ (.A(_19920_),
    .B(_20465_),
    .C(_20466_),
    .Y(_20467_));
 sky130_as_sc_hs__or2_2 _26968_ (.A(_20464_),
    .B(_20467_),
    .Y(_20468_));
 sky130_as_sc_hs__or2_2 _26969_ (.A(_20461_),
    .B(_20468_),
    .Y(_20469_));
 sky130_as_sc_hs__nor2_2 _26970_ (.A(_19504_),
    .B(_20039_),
    .Y(_20470_));
 sky130_as_sc_hs__or2_2 _26971_ (.A(_20469_),
    .B(_20470_),
    .Y(_20471_));
 sky130_as_sc_hs__nand2b_2 _26973_ (.B(net309),
    .Y(_20473_),
    .A(\tholin_riscv.regs[25][13] ));
 sky130_as_sc_hs__or2_2 _26974_ (.A(net309),
    .B(\tholin_riscv.regs[24][13] ),
    .Y(_20474_));
 sky130_as_sc_hs__nand3_2 _26975_ (.A(net174),
    .B(_20473_),
    .C(_20474_),
    .Y(_20475_));
 sky130_as_sc_hs__nand2b_2 _26976_ (.B(net309),
    .Y(_20476_),
    .A(\tholin_riscv.regs[27][13] ));
 sky130_as_sc_hs__or2_2 _26977_ (.A(net309),
    .B(\tholin_riscv.regs[26][13] ),
    .Y(_20477_));
 sky130_as_sc_hs__nand3_2 _26978_ (.A(net270),
    .B(_20476_),
    .C(_20477_),
    .Y(_20478_));
 sky130_as_sc_hs__nand3_2 _26979_ (.A(net158),
    .B(_20475_),
    .C(_20478_),
    .Y(_20479_));
 sky130_as_sc_hs__nand2b_2 _26980_ (.B(net309),
    .Y(_20480_),
    .A(\tholin_riscv.regs[29][13] ));
 sky130_as_sc_hs__or2_2 _26981_ (.A(net309),
    .B(\tholin_riscv.regs[28][13] ),
    .Y(_20481_));
 sky130_as_sc_hs__nand3_2 _26982_ (.A(net174),
    .B(_20480_),
    .C(_20481_),
    .Y(_20482_));
 sky130_as_sc_hs__nand2b_2 _26983_ (.B(net309),
    .Y(_20483_),
    .A(\tholin_riscv.regs[31][13] ));
 sky130_as_sc_hs__or2_2 _26984_ (.A(net309),
    .B(\tholin_riscv.regs[30][13] ),
    .Y(_20484_));
 sky130_as_sc_hs__nand3_2 _26985_ (.A(net270),
    .B(_20483_),
    .C(_20484_),
    .Y(_20485_));
 sky130_as_sc_hs__nand3_2 _26986_ (.A(net257),
    .B(_20482_),
    .C(_20485_),
    .Y(_20486_));
 sky130_as_sc_hs__nand2b_2 _26987_ (.B(net308),
    .Y(_20487_),
    .A(\tholin_riscv.regs[17][13] ));
 sky130_as_sc_hs__or2_2 _26988_ (.A(net308),
    .B(\tholin_riscv.regs[16][13] ),
    .Y(_20488_));
 sky130_as_sc_hs__nand3_2 _26989_ (.A(net174),
    .B(_20487_),
    .C(_20488_),
    .Y(_20489_));
 sky130_as_sc_hs__nand2b_2 _26990_ (.B(net308),
    .Y(_20490_),
    .A(\tholin_riscv.regs[19][13] ));
 sky130_as_sc_hs__or2_2 _26991_ (.A(net308),
    .B(\tholin_riscv.regs[18][13] ),
    .Y(_20491_));
 sky130_as_sc_hs__nand3_2 _26992_ (.A(net270),
    .B(_20490_),
    .C(_20491_),
    .Y(_20492_));
 sky130_as_sc_hs__nand3_2 _26993_ (.A(net158),
    .B(_20489_),
    .C(_20492_),
    .Y(_20493_));
 sky130_as_sc_hs__nand2b_2 _26994_ (.B(net308),
    .Y(_20494_),
    .A(\tholin_riscv.regs[23][13] ));
 sky130_as_sc_hs__or2_2 _26995_ (.A(net308),
    .B(\tholin_riscv.regs[22][13] ),
    .Y(_20495_));
 sky130_as_sc_hs__nand3_2 _26996_ (.A(net270),
    .B(_20494_),
    .C(_20495_),
    .Y(_20496_));
 sky130_as_sc_hs__nand2b_2 _26997_ (.B(net308),
    .Y(_20497_),
    .A(\tholin_riscv.regs[21][13] ));
 sky130_as_sc_hs__or2_2 _26998_ (.A(net308),
    .B(\tholin_riscv.regs[20][13] ),
    .Y(_20498_));
 sky130_as_sc_hs__nand3_2 _26999_ (.A(net174),
    .B(_20497_),
    .C(_20498_),
    .Y(_20499_));
 sky130_as_sc_hs__nand3_2 _27000_ (.A(net257),
    .B(_20496_),
    .C(_20499_),
    .Y(_20500_));
 sky130_as_sc_hs__nand3_2 _27001_ (.A(net152),
    .B(_20493_),
    .C(_20500_),
    .Y(_20501_));
 sky130_as_sc_hs__nand3_2 _27002_ (.A(net249),
    .B(_20479_),
    .C(_20486_),
    .Y(_20502_));
 sky130_as_sc_hs__nand3_2 _27003_ (.A(net248),
    .B(_20501_),
    .C(_20502_),
    .Y(_20503_));
 sky130_as_sc_hs__nand2b_2 _27004_ (.B(net314),
    .Y(_20504_),
    .A(\tholin_riscv.regs[9][13] ));
 sky130_as_sc_hs__or2_2 _27005_ (.A(net314),
    .B(\tholin_riscv.regs[8][13] ),
    .Y(_20505_));
 sky130_as_sc_hs__nand3_2 _27006_ (.A(net176),
    .B(_20504_),
    .C(_20505_),
    .Y(_20506_));
 sky130_as_sc_hs__nand2b_2 _27007_ (.B(net314),
    .Y(_20507_),
    .A(\tholin_riscv.regs[11][13] ));
 sky130_as_sc_hs__or2_2 _27008_ (.A(net314),
    .B(\tholin_riscv.regs[10][13] ),
    .Y(_20508_));
 sky130_as_sc_hs__nand3_2 _27009_ (.A(net272),
    .B(_20507_),
    .C(_20508_),
    .Y(_20509_));
 sky130_as_sc_hs__nand3_2 _27010_ (.A(net158),
    .B(_20506_),
    .C(_20509_),
    .Y(_20510_));
 sky130_as_sc_hs__nand2b_2 _27011_ (.B(net315),
    .Y(_20511_),
    .A(\tholin_riscv.regs[13][13] ));
 sky130_as_sc_hs__or2_2 _27012_ (.A(net315),
    .B(\tholin_riscv.regs[12][13] ),
    .Y(_20512_));
 sky130_as_sc_hs__nand3_2 _27013_ (.A(net176),
    .B(_20511_),
    .C(_20512_),
    .Y(_20513_));
 sky130_as_sc_hs__nand2b_2 _27014_ (.B(net315),
    .Y(_20514_),
    .A(\tholin_riscv.regs[15][13] ));
 sky130_as_sc_hs__or2_2 _27015_ (.A(net315),
    .B(\tholin_riscv.regs[14][13] ),
    .Y(_20515_));
 sky130_as_sc_hs__nand3_2 _27016_ (.A(net272),
    .B(_20514_),
    .C(_20515_),
    .Y(_20516_));
 sky130_as_sc_hs__nand3_2 _27017_ (.A(net258),
    .B(_20513_),
    .C(_20516_),
    .Y(_20517_));
 sky130_as_sc_hs__nand2b_2 _27018_ (.B(net315),
    .Y(_20518_),
    .A(\tholin_riscv.regs[1][13] ));
 sky130_as_sc_hs__or2_2 _27019_ (.A(net315),
    .B(\tholin_riscv.regs[0][13] ),
    .Y(_20519_));
 sky130_as_sc_hs__nand3_2 _27020_ (.A(net176),
    .B(_20518_),
    .C(_20519_),
    .Y(_20520_));
 sky130_as_sc_hs__nand2b_2 _27021_ (.B(net315),
    .Y(_20521_),
    .A(\tholin_riscv.regs[3][13] ));
 sky130_as_sc_hs__or2_2 _27022_ (.A(net315),
    .B(\tholin_riscv.regs[2][13] ),
    .Y(_20522_));
 sky130_as_sc_hs__nand3_2 _27023_ (.A(net272),
    .B(_20521_),
    .C(_20522_),
    .Y(_20523_));
 sky130_as_sc_hs__nand3_2 _27024_ (.A(net158),
    .B(_20520_),
    .C(_20523_),
    .Y(_20524_));
 sky130_as_sc_hs__nand2b_2 _27025_ (.B(net315),
    .Y(_20525_),
    .A(\tholin_riscv.regs[7][13] ));
 sky130_as_sc_hs__or2_2 _27026_ (.A(net315),
    .B(\tholin_riscv.regs[6][13] ),
    .Y(_20526_));
 sky130_as_sc_hs__nand3_2 _27027_ (.A(net272),
    .B(_20525_),
    .C(_20526_),
    .Y(_20527_));
 sky130_as_sc_hs__nand2b_2 _27028_ (.B(net315),
    .Y(_20528_),
    .A(\tholin_riscv.regs[5][13] ));
 sky130_as_sc_hs__or2_2 _27029_ (.A(net315),
    .B(\tholin_riscv.regs[4][13] ),
    .Y(_20529_));
 sky130_as_sc_hs__nand3_2 _27030_ (.A(net176),
    .B(_20528_),
    .C(_20529_),
    .Y(_20530_));
 sky130_as_sc_hs__nand3_2 _27031_ (.A(net258),
    .B(_20527_),
    .C(_20530_),
    .Y(_20531_));
 sky130_as_sc_hs__nand3_2 _27032_ (.A(net152),
    .B(_20524_),
    .C(_20531_),
    .Y(_20532_));
 sky130_as_sc_hs__nand3_2 _27033_ (.A(net249),
    .B(_20510_),
    .C(_20517_),
    .Y(_20533_));
 sky130_as_sc_hs__nand3_2 _27034_ (.A(net150),
    .B(_20532_),
    .C(_20533_),
    .Y(_20534_));
 sky130_as_sc_hs__inv_2 _27036_ (.Y(_20536_),
    .A(_20535_));
 sky130_as_sc_hs__or2_2 _27038_ (.A(net7),
    .B(_19755_),
    .Y(_20538_));
 sky130_as_sc_hs__nand3_2 _27039_ (.A(_19759_),
    .B(_20537_),
    .C(_20538_),
    .Y(_20539_));
 sky130_as_sc_hs__or2_2 _27040_ (.A(net1690),
    .B(_20021_),
    .Y(_20540_));
 sky130_as_sc_hs__nand3_2 _27041_ (.A(_20021_),
    .B(_20472_),
    .C(_20539_),
    .Y(_20541_));
 sky130_as_sc_hs__and2_2 _27042_ (.A(net497),
    .B(_20541_),
    .Y(_20542_));
 sky130_as_sc_hs__and2_2 _27043_ (.A(_20540_),
    .B(_20542_),
    .Y(_00010_));
 sky130_as_sc_hs__and2_2 _27048_ (.A(_20545_),
    .B(_20546_),
    .Y(_20547_));
 sky130_as_sc_hs__nand3_2 _27049_ (.A(_20543_),
    .B(_20544_),
    .C(_20547_),
    .Y(_20548_));
 sky130_as_sc_hs__nand3_2 _27055_ (.A(_19993_),
    .B(_20552_),
    .C(_20553_),
    .Y(_20554_));
 sky130_as_sc_hs__or2_2 _27056_ (.A(_20551_),
    .B(_20554_),
    .Y(_20555_));
 sky130_as_sc_hs__or2_2 _27057_ (.A(_20548_),
    .B(_20555_),
    .Y(_20556_));
 sky130_as_sc_hs__nor2_2 _27058_ (.A(_19503_),
    .B(_20039_),
    .Y(_20557_));
 sky130_as_sc_hs__or2_2 _27059_ (.A(_20556_),
    .B(_20557_),
    .Y(_20558_));
 sky130_as_sc_hs__nand2b_2 _27061_ (.B(net283),
    .Y(_20560_),
    .A(\tholin_riscv.regs[25][14] ));
 sky130_as_sc_hs__or2_2 _27062_ (.A(net284),
    .B(\tholin_riscv.regs[24][14] ),
    .Y(_20561_));
 sky130_as_sc_hs__nand3_2 _27063_ (.A(net166),
    .B(_20560_),
    .C(_20561_),
    .Y(_20562_));
 sky130_as_sc_hs__nand2b_2 _27064_ (.B(net283),
    .Y(_20563_),
    .A(\tholin_riscv.regs[27][14] ));
 sky130_as_sc_hs__or2_2 _27065_ (.A(net283),
    .B(\tholin_riscv.regs[26][14] ),
    .Y(_20564_));
 sky130_as_sc_hs__nand3_2 _27066_ (.A(net263),
    .B(_20563_),
    .C(_20564_),
    .Y(_20565_));
 sky130_as_sc_hs__nand3_2 _27067_ (.A(net157),
    .B(_20562_),
    .C(_20565_),
    .Y(_20566_));
 sky130_as_sc_hs__nand2b_2 _27068_ (.B(net283),
    .Y(_20567_),
    .A(\tholin_riscv.regs[29][14] ));
 sky130_as_sc_hs__or2_2 _27069_ (.A(net283),
    .B(\tholin_riscv.regs[28][14] ),
    .Y(_20568_));
 sky130_as_sc_hs__nand3_2 _27070_ (.A(net166),
    .B(_20567_),
    .C(_20568_),
    .Y(_20569_));
 sky130_as_sc_hs__nand2b_2 _27071_ (.B(net283),
    .Y(_20570_),
    .A(\tholin_riscv.regs[31][14] ));
 sky130_as_sc_hs__or2_2 _27072_ (.A(net283),
    .B(\tholin_riscv.regs[30][14] ),
    .Y(_20571_));
 sky130_as_sc_hs__nand3_2 _27073_ (.A(net263),
    .B(_20570_),
    .C(_20571_),
    .Y(_20572_));
 sky130_as_sc_hs__nand3_2 _27074_ (.A(net256),
    .B(_20569_),
    .C(_20572_),
    .Y(_20573_));
 sky130_as_sc_hs__nand2b_2 _27075_ (.B(net283),
    .Y(_20574_),
    .A(\tholin_riscv.regs[17][14] ));
 sky130_as_sc_hs__or2_2 _27076_ (.A(net283),
    .B(\tholin_riscv.regs[16][14] ),
    .Y(_20575_));
 sky130_as_sc_hs__nand3_2 _27077_ (.A(net166),
    .B(_20574_),
    .C(_20575_),
    .Y(_20576_));
 sky130_as_sc_hs__nand2b_2 _27078_ (.B(net283),
    .Y(_20577_),
    .A(\tholin_riscv.regs[19][14] ));
 sky130_as_sc_hs__or2_2 _27079_ (.A(net283),
    .B(\tholin_riscv.regs[18][14] ),
    .Y(_20578_));
 sky130_as_sc_hs__nand3_2 _27080_ (.A(net263),
    .B(_20577_),
    .C(_20578_),
    .Y(_20579_));
 sky130_as_sc_hs__nand3_2 _27081_ (.A(net157),
    .B(_20576_),
    .C(_20579_),
    .Y(_20580_));
 sky130_as_sc_hs__nand2b_2 _27082_ (.B(net283),
    .Y(_20581_),
    .A(\tholin_riscv.regs[23][14] ));
 sky130_as_sc_hs__or2_2 _27083_ (.A(net283),
    .B(\tholin_riscv.regs[22][14] ),
    .Y(_20582_));
 sky130_as_sc_hs__nand3_2 _27084_ (.A(net263),
    .B(_20581_),
    .C(_20582_),
    .Y(_20583_));
 sky130_as_sc_hs__nand2b_2 _27085_ (.B(net283),
    .Y(_20584_),
    .A(\tholin_riscv.regs[21][14] ));
 sky130_as_sc_hs__or2_2 _27086_ (.A(net283),
    .B(\tholin_riscv.regs[20][14] ),
    .Y(_20585_));
 sky130_as_sc_hs__nand3_2 _27087_ (.A(net166),
    .B(_20584_),
    .C(_20585_),
    .Y(_20586_));
 sky130_as_sc_hs__nand3_2 _27088_ (.A(net256),
    .B(_20583_),
    .C(_20586_),
    .Y(_20587_));
 sky130_as_sc_hs__nand3_2 _27089_ (.A(net153),
    .B(_20580_),
    .C(_20587_),
    .Y(_20588_));
 sky130_as_sc_hs__nand3_2 _27090_ (.A(net250),
    .B(_20566_),
    .C(_20573_),
    .Y(_20589_));
 sky130_as_sc_hs__nand3_2 _27091_ (.A(net248),
    .B(_20588_),
    .C(_20589_),
    .Y(_20590_));
 sky130_as_sc_hs__nand2b_2 _27092_ (.B(net284),
    .Y(_20591_),
    .A(\tholin_riscv.regs[9][14] ));
 sky130_as_sc_hs__or2_2 _27093_ (.A(net284),
    .B(\tholin_riscv.regs[8][14] ),
    .Y(_20592_));
 sky130_as_sc_hs__nand3_2 _27094_ (.A(net166),
    .B(_20591_),
    .C(_20592_),
    .Y(_20593_));
 sky130_as_sc_hs__nand2b_2 _27095_ (.B(net284),
    .Y(_20594_),
    .A(\tholin_riscv.regs[11][14] ));
 sky130_as_sc_hs__or2_2 _27096_ (.A(net284),
    .B(\tholin_riscv.regs[10][14] ),
    .Y(_20595_));
 sky130_as_sc_hs__nand3_2 _27097_ (.A(net263),
    .B(_20594_),
    .C(_20595_),
    .Y(_20596_));
 sky130_as_sc_hs__nand3_2 _27098_ (.A(net157),
    .B(_20593_),
    .C(_20596_),
    .Y(_20597_));
 sky130_as_sc_hs__nand2b_2 _27099_ (.B(net284),
    .Y(_20598_),
    .A(\tholin_riscv.regs[13][14] ));
 sky130_as_sc_hs__or2_2 _27100_ (.A(net284),
    .B(\tholin_riscv.regs[12][14] ),
    .Y(_20599_));
 sky130_as_sc_hs__nand3_2 _27101_ (.A(net166),
    .B(_20598_),
    .C(_20599_),
    .Y(_20600_));
 sky130_as_sc_hs__nand2b_2 _27102_ (.B(net287),
    .Y(_20601_),
    .A(\tholin_riscv.regs[15][14] ));
 sky130_as_sc_hs__or2_2 _27103_ (.A(net284),
    .B(\tholin_riscv.regs[14][14] ),
    .Y(_20602_));
 sky130_as_sc_hs__nand3_2 _27104_ (.A(net263),
    .B(_20601_),
    .C(_20602_),
    .Y(_20603_));
 sky130_as_sc_hs__nand3_2 _27105_ (.A(net256),
    .B(_20600_),
    .C(_20603_),
    .Y(_20604_));
 sky130_as_sc_hs__nand2b_2 _27106_ (.B(net284),
    .Y(_20605_),
    .A(\tholin_riscv.regs[1][14] ));
 sky130_as_sc_hs__or2_2 _27107_ (.A(net284),
    .B(\tholin_riscv.regs[0][14] ),
    .Y(_20606_));
 sky130_as_sc_hs__nand3_2 _27108_ (.A(net166),
    .B(_20605_),
    .C(_20606_),
    .Y(_20607_));
 sky130_as_sc_hs__nand2b_2 _27109_ (.B(net292),
    .Y(_20608_),
    .A(\tholin_riscv.regs[3][14] ));
 sky130_as_sc_hs__or2_2 _27110_ (.A(net292),
    .B(\tholin_riscv.regs[2][14] ),
    .Y(_20609_));
 sky130_as_sc_hs__nand3_2 _27111_ (.A(net282),
    .B(_20608_),
    .C(_20609_),
    .Y(_20610_));
 sky130_as_sc_hs__nand3_2 _27112_ (.A(net157),
    .B(_20607_),
    .C(_20610_),
    .Y(_20611_));
 sky130_as_sc_hs__nand2b_2 _27113_ (.B(net283),
    .Y(_20612_),
    .A(\tholin_riscv.regs[7][14] ));
 sky130_as_sc_hs__or2_2 _27114_ (.A(net284),
    .B(\tholin_riscv.regs[6][14] ),
    .Y(_20613_));
 sky130_as_sc_hs__nand3_2 _27115_ (.A(net263),
    .B(_20612_),
    .C(_20613_),
    .Y(_20614_));
 sky130_as_sc_hs__nand2b_2 _27116_ (.B(net292),
    .Y(_20615_),
    .A(\tholin_riscv.regs[5][14] ));
 sky130_as_sc_hs__or2_2 _27117_ (.A(net292),
    .B(\tholin_riscv.regs[4][14] ),
    .Y(_20616_));
 sky130_as_sc_hs__nand3_2 _27118_ (.A(net173),
    .B(_20615_),
    .C(_20616_),
    .Y(_20617_));
 sky130_as_sc_hs__nand3_2 _27119_ (.A(net256),
    .B(_20614_),
    .C(_20617_),
    .Y(_20618_));
 sky130_as_sc_hs__nand3_2 _27120_ (.A(net153),
    .B(_20611_),
    .C(_20618_),
    .Y(_20619_));
 sky130_as_sc_hs__nand3_2 _27121_ (.A(net250),
    .B(_20597_),
    .C(_20604_),
    .Y(_20620_));
 sky130_as_sc_hs__nand3_2 _27122_ (.A(net151),
    .B(_20619_),
    .C(_20620_),
    .Y(_20621_));
 sky130_as_sc_hs__and2_2 _27123_ (.A(_20590_),
    .B(_20621_),
    .Y(_20622_));
 sky130_as_sc_hs__or2_2 _27124_ (.A(_19754_),
    .B(_20622_),
    .Y(_20623_));
 sky130_as_sc_hs__or2_2 _27125_ (.A(net8),
    .B(_19755_),
    .Y(_20624_));
 sky130_as_sc_hs__nand3_2 _27126_ (.A(_19759_),
    .B(_20623_),
    .C(_20624_),
    .Y(_20625_));
 sky130_as_sc_hs__or2_2 _27127_ (.A(net411),
    .B(_20021_),
    .Y(_20626_));
 sky130_as_sc_hs__nand3_2 _27128_ (.A(_20021_),
    .B(_20559_),
    .C(_20625_),
    .Y(_20627_));
 sky130_as_sc_hs__and2_2 _27129_ (.A(net497),
    .B(_20627_),
    .Y(_20628_));
 sky130_as_sc_hs__and2_2 _27130_ (.A(_20626_),
    .B(_20628_),
    .Y(_00011_));
 sky130_as_sc_hs__nand3_2 _27140_ (.A(_20630_),
    .B(_20632_),
    .C(_20635_),
    .Y(_20638_));
 sky130_as_sc_hs__nand3_2 _27141_ (.A(_20633_),
    .B(_20634_),
    .C(_20636_),
    .Y(_20639_));
 sky130_as_sc_hs__or2_2 _27142_ (.A(_20637_),
    .B(_20639_),
    .Y(_20640_));
 sky130_as_sc_hs__nor2_2 _27143_ (.A(_20638_),
    .B(_20640_),
    .Y(_20641_));
 sky130_as_sc_hs__or2_2 _27144_ (.A(_19502_),
    .B(_20039_),
    .Y(_20642_));
 sky130_as_sc_hs__nand2b_2 _27147_ (.B(net285),
    .Y(_20645_),
    .A(\tholin_riscv.regs[25][15] ));
 sky130_as_sc_hs__or2_2 _27148_ (.A(net285),
    .B(\tholin_riscv.regs[24][15] ),
    .Y(_20646_));
 sky130_as_sc_hs__nand3_2 _27149_ (.A(net166),
    .B(_20645_),
    .C(_20646_),
    .Y(_20647_));
 sky130_as_sc_hs__nand2b_2 _27150_ (.B(net285),
    .Y(_20648_),
    .A(\tholin_riscv.regs[27][15] ));
 sky130_as_sc_hs__or2_2 _27151_ (.A(net285),
    .B(\tholin_riscv.regs[26][15] ),
    .Y(_20649_));
 sky130_as_sc_hs__nand3_2 _27152_ (.A(net263),
    .B(_20648_),
    .C(_20649_),
    .Y(_20650_));
 sky130_as_sc_hs__nand3_2 _27153_ (.A(net157),
    .B(_20647_),
    .C(_20650_),
    .Y(_20651_));
 sky130_as_sc_hs__nand2b_2 _27154_ (.B(net285),
    .Y(_20652_),
    .A(\tholin_riscv.regs[29][15] ));
 sky130_as_sc_hs__or2_2 _27155_ (.A(net285),
    .B(\tholin_riscv.regs[28][15] ),
    .Y(_20653_));
 sky130_as_sc_hs__nand3_2 _27156_ (.A(net166),
    .B(_20652_),
    .C(_20653_),
    .Y(_20654_));
 sky130_as_sc_hs__nand2b_2 _27157_ (.B(net285),
    .Y(_20655_),
    .A(\tholin_riscv.regs[31][15] ));
 sky130_as_sc_hs__or2_2 _27158_ (.A(net285),
    .B(\tholin_riscv.regs[30][15] ),
    .Y(_20656_));
 sky130_as_sc_hs__nand3_2 _27159_ (.A(net263),
    .B(_20655_),
    .C(_20656_),
    .Y(_20657_));
 sky130_as_sc_hs__nand3_2 _27160_ (.A(net256),
    .B(_20654_),
    .C(_20657_),
    .Y(_20658_));
 sky130_as_sc_hs__nand2b_2 _27161_ (.B(net285),
    .Y(_20659_),
    .A(\tholin_riscv.regs[17][15] ));
 sky130_as_sc_hs__or2_2 _27162_ (.A(net285),
    .B(\tholin_riscv.regs[16][15] ),
    .Y(_20660_));
 sky130_as_sc_hs__nand3_2 _27163_ (.A(net166),
    .B(_20659_),
    .C(_20660_),
    .Y(_20661_));
 sky130_as_sc_hs__nand2b_2 _27164_ (.B(net285),
    .Y(_20662_),
    .A(\tholin_riscv.regs[19][15] ));
 sky130_as_sc_hs__or2_2 _27165_ (.A(net285),
    .B(\tholin_riscv.regs[18][15] ),
    .Y(_20663_));
 sky130_as_sc_hs__nand3_2 _27166_ (.A(net263),
    .B(_20662_),
    .C(_20663_),
    .Y(_20664_));
 sky130_as_sc_hs__nand3_2 _27167_ (.A(net157),
    .B(_20661_),
    .C(_20664_),
    .Y(_20665_));
 sky130_as_sc_hs__nand2b_2 _27168_ (.B(net285),
    .Y(_20666_),
    .A(\tholin_riscv.regs[23][15] ));
 sky130_as_sc_hs__or2_2 _27169_ (.A(net285),
    .B(\tholin_riscv.regs[22][15] ),
    .Y(_20667_));
 sky130_as_sc_hs__nand3_2 _27170_ (.A(net263),
    .B(_20666_),
    .C(_20667_),
    .Y(_20668_));
 sky130_as_sc_hs__nand2b_2 _27171_ (.B(net285),
    .Y(_20669_),
    .A(\tholin_riscv.regs[21][15] ));
 sky130_as_sc_hs__or2_2 _27172_ (.A(net285),
    .B(\tholin_riscv.regs[20][15] ),
    .Y(_20670_));
 sky130_as_sc_hs__nand3_2 _27173_ (.A(net166),
    .B(_20669_),
    .C(_20670_),
    .Y(_20671_));
 sky130_as_sc_hs__nand3_2 _27174_ (.A(net256),
    .B(_20668_),
    .C(_20671_),
    .Y(_20672_));
 sky130_as_sc_hs__nand3_2 _27175_ (.A(net153),
    .B(_20665_),
    .C(_20672_),
    .Y(_20673_));
 sky130_as_sc_hs__nand3_2 _27176_ (.A(net250),
    .B(_20651_),
    .C(_20658_),
    .Y(_20674_));
 sky130_as_sc_hs__nand3_2 _27177_ (.A(net248),
    .B(_20673_),
    .C(_20674_),
    .Y(_20675_));
 sky130_as_sc_hs__nand2b_2 _27178_ (.B(net291),
    .Y(_20676_),
    .A(\tholin_riscv.regs[9][15] ));
 sky130_as_sc_hs__or2_2 _27179_ (.A(net286),
    .B(\tholin_riscv.regs[8][15] ),
    .Y(_20677_));
 sky130_as_sc_hs__nand3_2 _27180_ (.A(net166),
    .B(_20676_),
    .C(_20677_),
    .Y(_20678_));
 sky130_as_sc_hs__nand2b_2 _27181_ (.B(net286),
    .Y(_20679_),
    .A(\tholin_riscv.regs[11][15] ));
 sky130_as_sc_hs__or2_2 _27182_ (.A(net286),
    .B(\tholin_riscv.regs[10][15] ),
    .Y(_20680_));
 sky130_as_sc_hs__nand3_2 _27183_ (.A(net263),
    .B(_20679_),
    .C(_20680_),
    .Y(_20681_));
 sky130_as_sc_hs__nand3_2 _27184_ (.A(net157),
    .B(_20678_),
    .C(_20681_),
    .Y(_20682_));
 sky130_as_sc_hs__nand2b_2 _27185_ (.B(net311),
    .Y(_20683_),
    .A(\tholin_riscv.regs[13][15] ));
 sky130_as_sc_hs__or2_2 _27186_ (.A(net311),
    .B(\tholin_riscv.regs[12][15] ),
    .Y(_20684_));
 sky130_as_sc_hs__nand3_2 _27187_ (.A(net166),
    .B(_20683_),
    .C(_20684_),
    .Y(_20685_));
 sky130_as_sc_hs__nand2b_2 _27188_ (.B(net311),
    .Y(_20686_),
    .A(\tholin_riscv.regs[15][15] ));
 sky130_as_sc_hs__or2_2 _27189_ (.A(net311),
    .B(\tholin_riscv.regs[14][15] ),
    .Y(_20687_));
 sky130_as_sc_hs__nand3_2 _27190_ (.A(net270),
    .B(_20686_),
    .C(_20687_),
    .Y(_20688_));
 sky130_as_sc_hs__nand3_2 _27191_ (.A(net257),
    .B(_20685_),
    .C(_20688_),
    .Y(_20689_));
 sky130_as_sc_hs__nand2b_2 _27192_ (.B(net286),
    .Y(_20690_),
    .A(\tholin_riscv.regs[1][15] ));
 sky130_as_sc_hs__or2_2 _27193_ (.A(net286),
    .B(\tholin_riscv.regs[0][15] ),
    .Y(_20691_));
 sky130_as_sc_hs__nand3_2 _27194_ (.A(net166),
    .B(_20690_),
    .C(_20691_),
    .Y(_20692_));
 sky130_as_sc_hs__nand2b_2 _27195_ (.B(net286),
    .Y(_20693_),
    .A(\tholin_riscv.regs[3][15] ));
 sky130_as_sc_hs__or2_2 _27196_ (.A(net286),
    .B(\tholin_riscv.regs[2][15] ),
    .Y(_20694_));
 sky130_as_sc_hs__nand3_2 _27197_ (.A(net263),
    .B(_20693_),
    .C(_20694_),
    .Y(_20695_));
 sky130_as_sc_hs__nand3_2 _27198_ (.A(net157),
    .B(_20692_),
    .C(_20695_),
    .Y(_20696_));
 sky130_as_sc_hs__nand2b_2 _27199_ (.B(net286),
    .Y(_20697_),
    .A(\tholin_riscv.regs[7][15] ));
 sky130_as_sc_hs__or2_2 _27200_ (.A(net286),
    .B(\tholin_riscv.regs[6][15] ),
    .Y(_20698_));
 sky130_as_sc_hs__nand3_2 _27201_ (.A(net263),
    .B(_20697_),
    .C(_20698_),
    .Y(_20699_));
 sky130_as_sc_hs__nand2b_2 _27202_ (.B(net286),
    .Y(_20700_),
    .A(\tholin_riscv.regs[5][15] ));
 sky130_as_sc_hs__or2_2 _27203_ (.A(net286),
    .B(\tholin_riscv.regs[4][15] ),
    .Y(_20701_));
 sky130_as_sc_hs__nand3_2 _27204_ (.A(net167),
    .B(_20700_),
    .C(_20701_),
    .Y(_20702_));
 sky130_as_sc_hs__nand3_2 _27205_ (.A(net256),
    .B(_20699_),
    .C(_20702_),
    .Y(_20703_));
 sky130_as_sc_hs__nand3_2 _27206_ (.A(net153),
    .B(_20696_),
    .C(_20703_),
    .Y(_20704_));
 sky130_as_sc_hs__nand3_2 _27207_ (.A(net250),
    .B(_20682_),
    .C(_20689_),
    .Y(_20705_));
 sky130_as_sc_hs__nand3_2 _27208_ (.A(net151),
    .B(_20704_),
    .C(_20705_),
    .Y(_20706_));
 sky130_as_sc_hs__and2_2 _27209_ (.A(_20675_),
    .B(_20706_),
    .Y(_20707_));
 sky130_as_sc_hs__or2_2 _27210_ (.A(_19754_),
    .B(_20707_),
    .Y(_20708_));
 sky130_as_sc_hs__or2_2 _27211_ (.A(net9),
    .B(_19755_),
    .Y(_20709_));
 sky130_as_sc_hs__nand3_2 _27212_ (.A(_19759_),
    .B(_20708_),
    .C(_20709_),
    .Y(_20710_));
 sky130_as_sc_hs__or2_2 _27213_ (.A(net373),
    .B(_20021_),
    .Y(_20711_));
 sky130_as_sc_hs__nand3_2 _27214_ (.A(_20021_),
    .B(_20644_),
    .C(_20710_),
    .Y(_20712_));
 sky130_as_sc_hs__and2_2 _27215_ (.A(net497),
    .B(_20712_),
    .Y(_20713_));
 sky130_as_sc_hs__and2_2 _27216_ (.A(_20711_),
    .B(_20713_),
    .Y(_00012_));
 sky130_as_sc_hs__nor2_2 _27217_ (.A(_19905_),
    .B(_19919_),
    .Y(_20714_));
 sky130_as_sc_hs__or2_2 _27218_ (.A(_19924_),
    .B(_20714_),
    .Y(_20715_));
 sky130_as_sc_hs__and2_2 _27220_ (.A(_20019_),
    .B(_20716_),
    .Y(_20717_));
 sky130_as_sc_hs__and2_2 _27221_ (.A(_20018_),
    .B(_20717_),
    .Y(_20718_));
 sky130_as_sc_hs__or2_2 _27222_ (.A(_19907_),
    .B(_19911_),
    .Y(_20719_));
 sky130_as_sc_hs__or2_2 _27223_ (.A(_20714_),
    .B(_20719_),
    .Y(_20720_));
 sky130_as_sc_hs__nor2_2 _27224_ (.A(_19999_),
    .B(_20720_),
    .Y(_20721_));
 sky130_as_sc_hs__and2_2 _27226_ (.A(_19908_),
    .B(_19911_),
    .Y(_20723_));
 sky130_as_sc_hs__and2_2 _27228_ (.A(_19911_),
    .B(_19916_),
    .Y(_20725_));
 sky130_as_sc_hs__and2_2 _27230_ (.A(_19911_),
    .B(_19919_),
    .Y(_20727_));
 sky130_as_sc_hs__and2_2 _27232_ (.A(_20726_),
    .B(_20728_),
    .Y(_20729_));
 sky130_as_sc_hs__nand3_2 _27233_ (.A(_20722_),
    .B(_20724_),
    .C(_20729_),
    .Y(_20730_));
 sky130_as_sc_hs__and2_2 _27234_ (.A(_19904_),
    .B(_19916_),
    .Y(_20731_));
 sky130_as_sc_hs__and2_2 _27236_ (.A(_19904_),
    .B(_19912_),
    .Y(_20733_));
 sky130_as_sc_hs__and2_2 _27238_ (.A(_20732_),
    .B(_20734_),
    .Y(_20735_));
 sky130_as_sc_hs__and2_2 _27239_ (.A(_19911_),
    .B(_19912_),
    .Y(_20736_));
 sky130_as_sc_hs__and2_2 _27241_ (.A(_19904_),
    .B(_19908_),
    .Y(_20738_));
 sky130_as_sc_hs__nand3_2 _27243_ (.A(_20735_),
    .B(_20737_),
    .C(_20739_),
    .Y(_20740_));
 sky130_as_sc_hs__or2_2 _27244_ (.A(_20730_),
    .B(_20740_),
    .Y(_20741_));
 sky130_as_sc_hs__nor2_2 _27245_ (.A(_20721_),
    .B(_20741_),
    .Y(_20742_));
 sky130_as_sc_hs__and2_2 _27250_ (.A(_20745_),
    .B(_20746_),
    .Y(_20747_));
 sky130_as_sc_hs__nand3_2 _27251_ (.A(_20743_),
    .B(_20744_),
    .C(_20747_),
    .Y(_20748_));
 sky130_as_sc_hs__nand3_2 _27257_ (.A(_19993_),
    .B(_20752_),
    .C(_20753_),
    .Y(_20754_));
 sky130_as_sc_hs__or2_2 _27258_ (.A(_20751_),
    .B(_20754_),
    .Y(_20755_));
 sky130_as_sc_hs__nor2_2 _27259_ (.A(_20748_),
    .B(_20755_),
    .Y(_20756_));
 sky130_as_sc_hs__and2_2 _27263_ (.A(_20758_),
    .B(_20759_),
    .Y(_20760_));
 sky130_as_sc_hs__nand3_2 _27265_ (.A(net137),
    .B(_20757_),
    .C(_20761_),
    .Y(_20762_));
 sky130_as_sc_hs__nand2b_2 _27266_ (.B(net294),
    .Y(_20763_),
    .A(\tholin_riscv.regs[25][0] ));
 sky130_as_sc_hs__or2_2 _27267_ (.A(net295),
    .B(\tholin_riscv.regs[24][0] ),
    .Y(_20764_));
 sky130_as_sc_hs__nand3_2 _27268_ (.A(net168),
    .B(_20763_),
    .C(_20764_),
    .Y(_20765_));
 sky130_as_sc_hs__nand2b_2 _27269_ (.B(net295),
    .Y(_20766_),
    .A(\tholin_riscv.regs[27][0] ));
 sky130_as_sc_hs__or2_2 _27270_ (.A(net295),
    .B(\tholin_riscv.regs[26][0] ),
    .Y(_20767_));
 sky130_as_sc_hs__nand3_2 _27271_ (.A(net266),
    .B(_20766_),
    .C(_20767_),
    .Y(_20768_));
 sky130_as_sc_hs__nand3_2 _27272_ (.A(net162),
    .B(_20765_),
    .C(_20768_),
    .Y(_20769_));
 sky130_as_sc_hs__nand2b_2 _27273_ (.B(net295),
    .Y(_20770_),
    .A(\tholin_riscv.regs[29][0] ));
 sky130_as_sc_hs__or2_2 _27274_ (.A(net295),
    .B(\tholin_riscv.regs[28][0] ),
    .Y(_20771_));
 sky130_as_sc_hs__nand3_2 _27275_ (.A(net168),
    .B(_20770_),
    .C(_20771_),
    .Y(_20772_));
 sky130_as_sc_hs__nand2b_2 _27276_ (.B(net295),
    .Y(_20773_),
    .A(\tholin_riscv.regs[31][0] ));
 sky130_as_sc_hs__or2_2 _27277_ (.A(net295),
    .B(\tholin_riscv.regs[30][0] ),
    .Y(_20774_));
 sky130_as_sc_hs__nand3_2 _27278_ (.A(net265),
    .B(_20773_),
    .C(_20774_),
    .Y(_20775_));
 sky130_as_sc_hs__nand3_2 _27279_ (.A(net255),
    .B(_20772_),
    .C(_20775_),
    .Y(_20776_));
 sky130_as_sc_hs__nand2b_2 _27280_ (.B(net295),
    .Y(_20777_),
    .A(\tholin_riscv.regs[17][0] ));
 sky130_as_sc_hs__or2_2 _27281_ (.A(net295),
    .B(\tholin_riscv.regs[16][0] ),
    .Y(_20778_));
 sky130_as_sc_hs__nand3_2 _27282_ (.A(net168),
    .B(_20777_),
    .C(_20778_),
    .Y(_20779_));
 sky130_as_sc_hs__nand2b_2 _27283_ (.B(net295),
    .Y(_20780_),
    .A(\tholin_riscv.regs[19][0] ));
 sky130_as_sc_hs__or2_2 _27284_ (.A(net295),
    .B(\tholin_riscv.regs[18][0] ),
    .Y(_20781_));
 sky130_as_sc_hs__nand3_2 _27285_ (.A(net265),
    .B(_20780_),
    .C(_20781_),
    .Y(_20782_));
 sky130_as_sc_hs__nand3_2 _27286_ (.A(net161),
    .B(_20779_),
    .C(_20782_),
    .Y(_20783_));
 sky130_as_sc_hs__nand2b_2 _27287_ (.B(net295),
    .Y(_20784_),
    .A(\tholin_riscv.regs[23][0] ));
 sky130_as_sc_hs__or2_2 _27288_ (.A(net295),
    .B(\tholin_riscv.regs[22][0] ),
    .Y(_20785_));
 sky130_as_sc_hs__nand3_2 _27289_ (.A(net265),
    .B(_20784_),
    .C(_20785_),
    .Y(_20786_));
 sky130_as_sc_hs__nand2b_2 _27290_ (.B(net295),
    .Y(_20787_),
    .A(\tholin_riscv.regs[21][0] ));
 sky130_as_sc_hs__or2_2 _27291_ (.A(net295),
    .B(\tholin_riscv.regs[20][0] ),
    .Y(_20788_));
 sky130_as_sc_hs__nand3_2 _27292_ (.A(net168),
    .B(_20787_),
    .C(_20788_),
    .Y(_20789_));
 sky130_as_sc_hs__nand3_2 _27293_ (.A(net255),
    .B(_20786_),
    .C(_20789_),
    .Y(_20790_));
 sky130_as_sc_hs__nand3_2 _27294_ (.A(net154),
    .B(_20783_),
    .C(_20790_),
    .Y(_20791_));
 sky130_as_sc_hs__nand3_2 _27295_ (.A(net253),
    .B(_20769_),
    .C(_20776_),
    .Y(_20792_));
 sky130_as_sc_hs__nand3_2 _27296_ (.A(net247),
    .B(_20791_),
    .C(_20792_),
    .Y(_20793_));
 sky130_as_sc_hs__nand2b_2 _27297_ (.B(net298),
    .Y(_20794_),
    .A(\tholin_riscv.regs[9][0] ));
 sky130_as_sc_hs__or2_2 _27298_ (.A(net296),
    .B(\tholin_riscv.regs[8][0] ),
    .Y(_20795_));
 sky130_as_sc_hs__nand3_2 _27299_ (.A(net169),
    .B(_20794_),
    .C(_20795_),
    .Y(_20796_));
 sky130_as_sc_hs__nand2b_2 _27300_ (.B(net296),
    .Y(_20797_),
    .A(\tholin_riscv.regs[11][0] ));
 sky130_as_sc_hs__or2_2 _27301_ (.A(net296),
    .B(\tholin_riscv.regs[10][0] ),
    .Y(_20798_));
 sky130_as_sc_hs__nand3_2 _27302_ (.A(net266),
    .B(_20797_),
    .C(_20798_),
    .Y(_20799_));
 sky130_as_sc_hs__nand3_2 _27303_ (.A(net162),
    .B(_20796_),
    .C(_20799_),
    .Y(_20800_));
 sky130_as_sc_hs__nand2b_2 _27304_ (.B(net296),
    .Y(_20801_),
    .A(\tholin_riscv.regs[13][0] ));
 sky130_as_sc_hs__or2_2 _27305_ (.A(net296),
    .B(\tholin_riscv.regs[12][0] ),
    .Y(_20802_));
 sky130_as_sc_hs__nand3_2 _27306_ (.A(net169),
    .B(_20801_),
    .C(_20802_),
    .Y(_20803_));
 sky130_as_sc_hs__nand2b_2 _27307_ (.B(net296),
    .Y(_20804_),
    .A(\tholin_riscv.regs[15][0] ));
 sky130_as_sc_hs__or2_2 _27308_ (.A(net296),
    .B(\tholin_riscv.regs[14][0] ),
    .Y(_20805_));
 sky130_as_sc_hs__nand3_2 _27309_ (.A(net266),
    .B(_20804_),
    .C(_20805_),
    .Y(_20806_));
 sky130_as_sc_hs__nand3_2 _27310_ (.A(net255),
    .B(_20803_),
    .C(_20806_),
    .Y(_20807_));
 sky130_as_sc_hs__nand2b_2 _27311_ (.B(net296),
    .Y(_20808_),
    .A(\tholin_riscv.regs[1][0] ));
 sky130_as_sc_hs__or2_2 _27312_ (.A(net296),
    .B(\tholin_riscv.regs[0][0] ),
    .Y(_20809_));
 sky130_as_sc_hs__nand3_2 _27313_ (.A(net169),
    .B(_20808_),
    .C(_20809_),
    .Y(_20810_));
 sky130_as_sc_hs__nand2b_2 _27314_ (.B(net297),
    .Y(_20811_),
    .A(\tholin_riscv.regs[3][0] ));
 sky130_as_sc_hs__or2_2 _27315_ (.A(net307),
    .B(\tholin_riscv.regs[2][0] ),
    .Y(_20812_));
 sky130_as_sc_hs__nand3_2 _27316_ (.A(net266),
    .B(_20811_),
    .C(_20812_),
    .Y(_20813_));
 sky130_as_sc_hs__nand3_2 _27317_ (.A(net162),
    .B(_20810_),
    .C(_20813_),
    .Y(_20814_));
 sky130_as_sc_hs__nand2b_2 _27318_ (.B(net296),
    .Y(_20815_),
    .A(\tholin_riscv.regs[7][0] ));
 sky130_as_sc_hs__or2_2 _27319_ (.A(net307),
    .B(\tholin_riscv.regs[6][0] ),
    .Y(_20816_));
 sky130_as_sc_hs__nand3_2 _27320_ (.A(net266),
    .B(_20815_),
    .C(_20816_),
    .Y(_20817_));
 sky130_as_sc_hs__nand2b_2 _27321_ (.B(net296),
    .Y(_20818_),
    .A(\tholin_riscv.regs[5][0] ));
 sky130_as_sc_hs__or2_2 _27322_ (.A(net307),
    .B(\tholin_riscv.regs[4][0] ),
    .Y(_20819_));
 sky130_as_sc_hs__nand3_2 _27323_ (.A(net169),
    .B(_20818_),
    .C(_20819_),
    .Y(_20820_));
 sky130_as_sc_hs__nand3_2 _27324_ (.A(net255),
    .B(_20817_),
    .C(_20820_),
    .Y(_20821_));
 sky130_as_sc_hs__nand3_2 _27325_ (.A(net154),
    .B(_20814_),
    .C(_20821_),
    .Y(_20822_));
 sky130_as_sc_hs__nand3_2 _27326_ (.A(net251),
    .B(_20800_),
    .C(_20807_),
    .Y(_20823_));
 sky130_as_sc_hs__nand3_2 _27327_ (.A(net151),
    .B(_20822_),
    .C(_20823_),
    .Y(_20824_));
 sky130_as_sc_hs__and2_2 _27328_ (.A(_20793_),
    .B(_20824_),
    .Y(_20825_));
 sky130_as_sc_hs__nand3_2 _27333_ (.A(_19754_),
    .B(_20828_),
    .C(_20829_),
    .Y(_20830_));
 sky130_as_sc_hs__nand3_2 _27334_ (.A(_19759_),
    .B(_20827_),
    .C(_20830_),
    .Y(_20831_));
 sky130_as_sc_hs__nand3_2 _27335_ (.A(_20718_),
    .B(_20762_),
    .C(_20831_),
    .Y(_20832_));
 sky130_as_sc_hs__or2_2 _27336_ (.A(\tholin_riscv.instr[0] ),
    .B(_20718_),
    .Y(_20833_));
 sky130_as_sc_hs__and2_2 _27337_ (.A(net500),
    .B(_20832_),
    .Y(_20834_));
 sky130_as_sc_hs__and2_2 _27338_ (.A(_20833_),
    .B(_20834_),
    .Y(_00013_));
 sky130_as_sc_hs__and2_2 _27343_ (.A(_20837_),
    .B(_20838_),
    .Y(_20839_));
 sky130_as_sc_hs__nand3_2 _27344_ (.A(_20835_),
    .B(_20836_),
    .C(_20839_),
    .Y(_20840_));
 sky130_as_sc_hs__and2_2 _27349_ (.A(_20843_),
    .B(_20844_),
    .Y(_20845_));
 sky130_as_sc_hs__nand3_2 _27350_ (.A(_20841_),
    .B(_20842_),
    .C(_20845_),
    .Y(_20846_));
 sky130_as_sc_hs__or2_2 _27351_ (.A(_20840_),
    .B(_20846_),
    .Y(_20847_));
 sky130_as_sc_hs__nor2_2 _27352_ (.A(_20721_),
    .B(_20847_),
    .Y(_20848_));
 sky130_as_sc_hs__and2_2 _27355_ (.A(_20849_),
    .B(_20850_),
    .Y(_20851_));
 sky130_as_sc_hs__nand3_2 _27358_ (.A(_20851_),
    .B(_20852_),
    .C(_20853_),
    .Y(_20854_));
 sky130_as_sc_hs__nand3_2 _27364_ (.A(_19993_),
    .B(_20858_),
    .C(_20859_),
    .Y(_20860_));
 sky130_as_sc_hs__or2_2 _27365_ (.A(_20857_),
    .B(_20860_),
    .Y(_20861_));
 sky130_as_sc_hs__nor2_2 _27366_ (.A(_20854_),
    .B(_20861_),
    .Y(_20862_));
 sky130_as_sc_hs__and2_2 _27370_ (.A(_20864_),
    .B(_20865_),
    .Y(_20866_));
 sky130_as_sc_hs__nand3_2 _27372_ (.A(_19758_),
    .B(_20863_),
    .C(_20867_),
    .Y(_20868_));
 sky130_as_sc_hs__nand2b_2 _27373_ (.B(net297),
    .Y(_20869_),
    .A(\tholin_riscv.regs[25][1] ));
 sky130_as_sc_hs__or2_2 _27374_ (.A(net296),
    .B(\tholin_riscv.regs[24][1] ),
    .Y(_20870_));
 sky130_as_sc_hs__nand3_2 _27375_ (.A(net169),
    .B(_20869_),
    .C(_20870_),
    .Y(_20871_));
 sky130_as_sc_hs__nand2b_2 _27376_ (.B(net296),
    .Y(_20872_),
    .A(\tholin_riscv.regs[27][1] ));
 sky130_as_sc_hs__or2_2 _27377_ (.A(net296),
    .B(\tholin_riscv.regs[26][1] ),
    .Y(_20873_));
 sky130_as_sc_hs__nand3_2 _27378_ (.A(net265),
    .B(_20872_),
    .C(_20873_),
    .Y(_20874_));
 sky130_as_sc_hs__nand3_2 _27379_ (.A(net162),
    .B(_20871_),
    .C(_20874_),
    .Y(_20875_));
 sky130_as_sc_hs__nand2b_2 _27380_ (.B(net296),
    .Y(_20876_),
    .A(\tholin_riscv.regs[29][1] ));
 sky130_as_sc_hs__or2_2 _27381_ (.A(net296),
    .B(\tholin_riscv.regs[28][1] ),
    .Y(_20877_));
 sky130_as_sc_hs__nand3_2 _27382_ (.A(net169),
    .B(_20876_),
    .C(_20877_),
    .Y(_20878_));
 sky130_as_sc_hs__nand2b_2 _27383_ (.B(net297),
    .Y(_20879_),
    .A(\tholin_riscv.regs[31][1] ));
 sky130_as_sc_hs__or2_2 _27384_ (.A(net297),
    .B(\tholin_riscv.regs[30][1] ),
    .Y(_20880_));
 sky130_as_sc_hs__nand3_2 _27385_ (.A(net265),
    .B(_20879_),
    .C(_20880_),
    .Y(_20881_));
 sky130_as_sc_hs__nand3_2 _27386_ (.A(net255),
    .B(_20878_),
    .C(_20881_),
    .Y(_20882_));
 sky130_as_sc_hs__nand2b_2 _27387_ (.B(net297),
    .Y(_20883_),
    .A(\tholin_riscv.regs[17][1] ));
 sky130_as_sc_hs__or2_2 _27388_ (.A(net297),
    .B(\tholin_riscv.regs[16][1] ),
    .Y(_20884_));
 sky130_as_sc_hs__nand3_2 _27389_ (.A(net169),
    .B(_20883_),
    .C(_20884_),
    .Y(_20885_));
 sky130_as_sc_hs__nand2b_2 _27390_ (.B(net297),
    .Y(_20886_),
    .A(\tholin_riscv.regs[19][1] ));
 sky130_as_sc_hs__or2_2 _27391_ (.A(net297),
    .B(\tholin_riscv.regs[18][1] ),
    .Y(_20887_));
 sky130_as_sc_hs__nand3_2 _27392_ (.A(net265),
    .B(_20886_),
    .C(_20887_),
    .Y(_20888_));
 sky130_as_sc_hs__nand3_2 _27393_ (.A(net162),
    .B(_20885_),
    .C(_20888_),
    .Y(_20889_));
 sky130_as_sc_hs__nand2b_2 _27394_ (.B(net297),
    .Y(_20890_),
    .A(\tholin_riscv.regs[23][1] ));
 sky130_as_sc_hs__or2_2 _27395_ (.A(net297),
    .B(\tholin_riscv.regs[22][1] ),
    .Y(_20891_));
 sky130_as_sc_hs__nand3_2 _27396_ (.A(net266),
    .B(_20890_),
    .C(_20891_),
    .Y(_20892_));
 sky130_as_sc_hs__nand2b_2 _27397_ (.B(net297),
    .Y(_20893_),
    .A(\tholin_riscv.regs[21][1] ));
 sky130_as_sc_hs__or2_2 _27398_ (.A(net297),
    .B(\tholin_riscv.regs[20][1] ),
    .Y(_20894_));
 sky130_as_sc_hs__nand3_2 _27399_ (.A(net169),
    .B(_20893_),
    .C(_20894_),
    .Y(_20895_));
 sky130_as_sc_hs__nand3_2 _27400_ (.A(net255),
    .B(_20892_),
    .C(_20895_),
    .Y(_20896_));
 sky130_as_sc_hs__nand3_2 _27401_ (.A(net154),
    .B(_20889_),
    .C(_20896_),
    .Y(_20897_));
 sky130_as_sc_hs__nand3_2 _27402_ (.A(net251),
    .B(_20875_),
    .C(_20882_),
    .Y(_20898_));
 sky130_as_sc_hs__nand3_2 _27403_ (.A(net247),
    .B(_20897_),
    .C(_20898_),
    .Y(_20899_));
 sky130_as_sc_hs__nand2b_2 _27404_ (.B(net304),
    .Y(_20900_),
    .A(\tholin_riscv.regs[9][1] ));
 sky130_as_sc_hs__or2_2 _27405_ (.A(net303),
    .B(\tholin_riscv.regs[8][1] ),
    .Y(_20901_));
 sky130_as_sc_hs__nand3_2 _27406_ (.A(net169),
    .B(_20900_),
    .C(_20901_),
    .Y(_20902_));
 sky130_as_sc_hs__nand2b_2 _27407_ (.B(net304),
    .Y(_20903_),
    .A(\tholin_riscv.regs[11][1] ));
 sky130_as_sc_hs__or2_2 _27408_ (.A(net304),
    .B(\tholin_riscv.regs[10][1] ),
    .Y(_20904_));
 sky130_as_sc_hs__nand3_2 _27409_ (.A(net268),
    .B(_20903_),
    .C(_20904_),
    .Y(_20905_));
 sky130_as_sc_hs__nand3_2 _27410_ (.A(net162),
    .B(_20902_),
    .C(_20905_),
    .Y(_20906_));
 sky130_as_sc_hs__nand2b_2 _27411_ (.B(net298),
    .Y(_20907_),
    .A(\tholin_riscv.regs[13][1] ));
 sky130_as_sc_hs__or2_2 _27412_ (.A(net298),
    .B(\tholin_riscv.regs[12][1] ),
    .Y(_20908_));
 sky130_as_sc_hs__nand3_2 _27413_ (.A(net169),
    .B(_20907_),
    .C(_20908_),
    .Y(_20909_));
 sky130_as_sc_hs__nand2b_2 _27414_ (.B(net297),
    .Y(_20910_),
    .A(\tholin_riscv.regs[15][1] ));
 sky130_as_sc_hs__or2_2 _27415_ (.A(net297),
    .B(\tholin_riscv.regs[14][1] ),
    .Y(_20911_));
 sky130_as_sc_hs__nand3_2 _27416_ (.A(net266),
    .B(_20910_),
    .C(_20911_),
    .Y(_20912_));
 sky130_as_sc_hs__nand3_2 _27417_ (.A(net255),
    .B(_20909_),
    .C(_20912_),
    .Y(_20913_));
 sky130_as_sc_hs__nand2b_2 _27418_ (.B(net298),
    .Y(_20914_),
    .A(\tholin_riscv.regs[1][1] ));
 sky130_as_sc_hs__or2_2 _27419_ (.A(net298),
    .B(\tholin_riscv.regs[0][1] ),
    .Y(_20915_));
 sky130_as_sc_hs__nand3_2 _27420_ (.A(net169),
    .B(_20914_),
    .C(_20915_),
    .Y(_20916_));
 sky130_as_sc_hs__nand2b_2 _27421_ (.B(net298),
    .Y(_20917_),
    .A(\tholin_riscv.regs[3][1] ));
 sky130_as_sc_hs__or2_2 _27422_ (.A(net298),
    .B(\tholin_riscv.regs[2][1] ),
    .Y(_20918_));
 sky130_as_sc_hs__nand3_2 _27423_ (.A(net266),
    .B(_20917_),
    .C(_20918_),
    .Y(_20919_));
 sky130_as_sc_hs__nand3_2 _27424_ (.A(net162),
    .B(_20916_),
    .C(_20919_),
    .Y(_20920_));
 sky130_as_sc_hs__nand2b_2 _27425_ (.B(net303),
    .Y(_20921_),
    .A(\tholin_riscv.regs[7][1] ));
 sky130_as_sc_hs__or2_2 _27426_ (.A(net303),
    .B(\tholin_riscv.regs[6][1] ),
    .Y(_20922_));
 sky130_as_sc_hs__nand3_2 _27427_ (.A(net268),
    .B(_20921_),
    .C(_20922_),
    .Y(_20923_));
 sky130_as_sc_hs__nand2b_2 _27428_ (.B(net303),
    .Y(_20924_),
    .A(\tholin_riscv.regs[5][1] ));
 sky130_as_sc_hs__or2_2 _27429_ (.A(net303),
    .B(\tholin_riscv.regs[4][1] ),
    .Y(_20925_));
 sky130_as_sc_hs__nand3_2 _27430_ (.A(net171),
    .B(_20924_),
    .C(_20925_),
    .Y(_20926_));
 sky130_as_sc_hs__nand3_2 _27431_ (.A(net254),
    .B(_20923_),
    .C(_20926_),
    .Y(_20927_));
 sky130_as_sc_hs__nand3_2 _27432_ (.A(net154),
    .B(_20920_),
    .C(_20927_),
    .Y(_20928_));
 sky130_as_sc_hs__nand3_2 _27433_ (.A(net251),
    .B(_20906_),
    .C(_20913_),
    .Y(_20929_));
 sky130_as_sc_hs__nand3_2 _27434_ (.A(net151),
    .B(_20928_),
    .C(_20929_),
    .Y(_20930_));
 sky130_as_sc_hs__and2_2 _27435_ (.A(_20899_),
    .B(_20930_),
    .Y(_20931_));
 sky130_as_sc_hs__nand3_2 _27440_ (.A(_19754_),
    .B(_20934_),
    .C(_20935_),
    .Y(_20936_));
 sky130_as_sc_hs__nand3_2 _27441_ (.A(_19759_),
    .B(_20933_),
    .C(_20936_),
    .Y(_20937_));
 sky130_as_sc_hs__nand3_2 _27442_ (.A(_20718_),
    .B(_20868_),
    .C(_20937_),
    .Y(_20938_));
 sky130_as_sc_hs__or2_2 _27443_ (.A(net1684),
    .B(_20718_),
    .Y(_20939_));
 sky130_as_sc_hs__and2_2 _27444_ (.A(net500),
    .B(_20938_),
    .Y(_20940_));
 sky130_as_sc_hs__and2_2 _27445_ (.A(_20939_),
    .B(_20940_),
    .Y(_00014_));
 sky130_as_sc_hs__and2_2 _27455_ (.A(_20948_),
    .B(_20949_),
    .Y(_20950_));
 sky130_as_sc_hs__nand3_2 _27464_ (.A(_20942_),
    .B(_20946_),
    .C(_20956_),
    .Y(_20959_));
 sky130_as_sc_hs__and2_2 _27465_ (.A(_20941_),
    .B(_20944_),
    .Y(_20960_));
 sky130_as_sc_hs__nand3_2 _27466_ (.A(_20945_),
    .B(_20957_),
    .C(_20960_),
    .Y(_20961_));
 sky130_as_sc_hs__or2_2 _27467_ (.A(_20959_),
    .B(_20961_),
    .Y(_20962_));
 sky130_as_sc_hs__nor2_2 _27468_ (.A(_20721_),
    .B(_20962_),
    .Y(_20963_));
 sky130_as_sc_hs__nand3_2 _27469_ (.A(_20950_),
    .B(_20953_),
    .C(_20954_),
    .Y(_20964_));
 sky130_as_sc_hs__nand3_2 _27470_ (.A(_20943_),
    .B(_20947_),
    .C(_20952_),
    .Y(_20965_));
 sky130_as_sc_hs__or2_2 _27471_ (.A(_20958_),
    .B(_20965_),
    .Y(_20966_));
 sky130_as_sc_hs__nor2_2 _27472_ (.A(_20964_),
    .B(_20966_),
    .Y(_20967_));
 sky130_as_sc_hs__and2_2 _27476_ (.A(_20969_),
    .B(_20970_),
    .Y(_20971_));
 sky130_as_sc_hs__nand3_2 _27478_ (.A(_19758_),
    .B(_20968_),
    .C(_20972_),
    .Y(_20973_));
 sky130_as_sc_hs__nand2b_2 _27479_ (.B(net292),
    .Y(_20974_),
    .A(\tholin_riscv.regs[25][2] ));
 sky130_as_sc_hs__or2_2 _27480_ (.A(net292),
    .B(\tholin_riscv.regs[24][2] ),
    .Y(_20975_));
 sky130_as_sc_hs__nand3_2 _27481_ (.A(net173),
    .B(_20974_),
    .C(_20975_),
    .Y(_20976_));
 sky130_as_sc_hs__nand2b_2 _27482_ (.B(net299),
    .Y(_20977_),
    .A(\tholin_riscv.regs[27][2] ));
 sky130_as_sc_hs__or2_2 _27483_ (.A(net288),
    .B(\tholin_riscv.regs[26][2] ),
    .Y(_20978_));
 sky130_as_sc_hs__nand3_2 _27484_ (.A(net267),
    .B(_20977_),
    .C(_20978_),
    .Y(_20979_));
 sky130_as_sc_hs__nand3_2 _27485_ (.A(net161),
    .B(_20976_),
    .C(_20979_),
    .Y(_20980_));
 sky130_as_sc_hs__nand2b_2 _27486_ (.B(net299),
    .Y(_20981_),
    .A(\tholin_riscv.regs[29][2] ));
 sky130_as_sc_hs__or2_2 _27487_ (.A(net299),
    .B(\tholin_riscv.regs[28][2] ),
    .Y(_20982_));
 sky130_as_sc_hs__nand3_2 _27488_ (.A(net168),
    .B(_20981_),
    .C(_20982_),
    .Y(_20983_));
 sky130_as_sc_hs__nand2b_2 _27489_ (.B(net293),
    .Y(_20984_),
    .A(\tholin_riscv.regs[31][2] ));
 sky130_as_sc_hs__or2_2 _27490_ (.A(net293),
    .B(\tholin_riscv.regs[30][2] ),
    .Y(_20985_));
 sky130_as_sc_hs__nand3_2 _27491_ (.A(net265),
    .B(_20984_),
    .C(_20985_),
    .Y(_20986_));
 sky130_as_sc_hs__nand3_2 _27492_ (.A(net255),
    .B(_20983_),
    .C(_20986_),
    .Y(_20987_));
 sky130_as_sc_hs__nand2b_2 _27493_ (.B(net292),
    .Y(_20988_),
    .A(\tholin_riscv.regs[17][2] ));
 sky130_as_sc_hs__or2_2 _27494_ (.A(net292),
    .B(\tholin_riscv.regs[16][2] ),
    .Y(_20989_));
 sky130_as_sc_hs__nand3_2 _27495_ (.A(net168),
    .B(_20988_),
    .C(_20989_),
    .Y(_20990_));
 sky130_as_sc_hs__nand2b_2 _27496_ (.B(net293),
    .Y(_20991_),
    .A(\tholin_riscv.regs[19][2] ));
 sky130_as_sc_hs__or2_2 _27497_ (.A(net293),
    .B(\tholin_riscv.regs[18][2] ),
    .Y(_20992_));
 sky130_as_sc_hs__nand3_2 _27498_ (.A(net265),
    .B(_20991_),
    .C(_20992_),
    .Y(_20993_));
 sky130_as_sc_hs__nand3_2 _27499_ (.A(net161),
    .B(_20990_),
    .C(_20993_),
    .Y(_20994_));
 sky130_as_sc_hs__nand2b_2 _27500_ (.B(net293),
    .Y(_20995_),
    .A(\tholin_riscv.regs[23][2] ));
 sky130_as_sc_hs__or2_2 _27501_ (.A(net293),
    .B(\tholin_riscv.regs[22][2] ),
    .Y(_20996_));
 sky130_as_sc_hs__nand3_2 _27502_ (.A(net265),
    .B(_20995_),
    .C(_20996_),
    .Y(_20997_));
 sky130_as_sc_hs__nand2b_2 _27503_ (.B(net293),
    .Y(_20998_),
    .A(\tholin_riscv.regs[21][2] ));
 sky130_as_sc_hs__or2_2 _27504_ (.A(net293),
    .B(\tholin_riscv.regs[20][2] ),
    .Y(_20999_));
 sky130_as_sc_hs__nand3_2 _27505_ (.A(net168),
    .B(_20998_),
    .C(_20999_),
    .Y(_21000_));
 sky130_as_sc_hs__nand3_2 _27506_ (.A(net255),
    .B(_20997_),
    .C(_21000_),
    .Y(_21001_));
 sky130_as_sc_hs__nand3_2 _27507_ (.A(net154),
    .B(_20994_),
    .C(_21001_),
    .Y(_21002_));
 sky130_as_sc_hs__nand3_2 _27508_ (.A(net251),
    .B(_20980_),
    .C(_20987_),
    .Y(_21003_));
 sky130_as_sc_hs__nand3_2 _27509_ (.A(net247),
    .B(_21002_),
    .C(_21003_),
    .Y(_21004_));
 sky130_as_sc_hs__nand2b_2 _27510_ (.B(net300),
    .Y(_21005_),
    .A(\tholin_riscv.regs[9][2] ));
 sky130_as_sc_hs__or2_2 _27511_ (.A(net300),
    .B(\tholin_riscv.regs[8][2] ),
    .Y(_21006_));
 sky130_as_sc_hs__nand3_2 _27512_ (.A(net168),
    .B(_21005_),
    .C(_21006_),
    .Y(_21007_));
 sky130_as_sc_hs__nand2b_2 _27513_ (.B(net293),
    .Y(_21008_),
    .A(\tholin_riscv.regs[11][2] ));
 sky130_as_sc_hs__or2_2 _27514_ (.A(net294),
    .B(\tholin_riscv.regs[10][2] ),
    .Y(_21009_));
 sky130_as_sc_hs__nand3_2 _27515_ (.A(net265),
    .B(_21008_),
    .C(_21009_),
    .Y(_21010_));
 sky130_as_sc_hs__nand3_2 _27516_ (.A(net161),
    .B(_21007_),
    .C(_21010_),
    .Y(_21011_));
 sky130_as_sc_hs__nand2b_2 _27517_ (.B(net293),
    .Y(_21012_),
    .A(\tholin_riscv.regs[13][2] ));
 sky130_as_sc_hs__or2_2 _27518_ (.A(net299),
    .B(\tholin_riscv.regs[12][2] ),
    .Y(_21013_));
 sky130_as_sc_hs__nand3_2 _27519_ (.A(net168),
    .B(_21012_),
    .C(_21013_),
    .Y(_21014_));
 sky130_as_sc_hs__nand2b_2 _27520_ (.B(net293),
    .Y(_21015_),
    .A(\tholin_riscv.regs[15][2] ));
 sky130_as_sc_hs__or2_2 _27521_ (.A(net293),
    .B(\tholin_riscv.regs[14][2] ),
    .Y(_21016_));
 sky130_as_sc_hs__nand3_2 _27522_ (.A(net265),
    .B(_21015_),
    .C(_21016_),
    .Y(_21017_));
 sky130_as_sc_hs__nand3_2 _27523_ (.A(net255),
    .B(_21014_),
    .C(_21017_),
    .Y(_21018_));
 sky130_as_sc_hs__nand2b_2 _27524_ (.B(net294),
    .Y(_21019_),
    .A(\tholin_riscv.regs[1][2] ));
 sky130_as_sc_hs__or2_2 _27525_ (.A(net294),
    .B(\tholin_riscv.regs[0][2] ),
    .Y(_21020_));
 sky130_as_sc_hs__nand3_2 _27526_ (.A(net168),
    .B(_21019_),
    .C(_21020_),
    .Y(_21021_));
 sky130_as_sc_hs__nand2b_2 _27527_ (.B(net294),
    .Y(_21022_),
    .A(\tholin_riscv.regs[3][2] ));
 sky130_as_sc_hs__or2_2 _27528_ (.A(net294),
    .B(\tholin_riscv.regs[2][2] ),
    .Y(_21023_));
 sky130_as_sc_hs__nand3_2 _27529_ (.A(net265),
    .B(_21022_),
    .C(_21023_),
    .Y(_21024_));
 sky130_as_sc_hs__nand3_2 _27530_ (.A(net161),
    .B(_21021_),
    .C(_21024_),
    .Y(_21025_));
 sky130_as_sc_hs__nand2b_2 _27531_ (.B(net293),
    .Y(_21026_),
    .A(\tholin_riscv.regs[7][2] ));
 sky130_as_sc_hs__or2_2 _27532_ (.A(net293),
    .B(\tholin_riscv.regs[6][2] ),
    .Y(_21027_));
 sky130_as_sc_hs__nand3_2 _27533_ (.A(net265),
    .B(_21026_),
    .C(_21027_),
    .Y(_21028_));
 sky130_as_sc_hs__nand2b_2 _27534_ (.B(net293),
    .Y(_21029_),
    .A(\tholin_riscv.regs[5][2] ));
 sky130_as_sc_hs__or2_2 _27535_ (.A(net293),
    .B(\tholin_riscv.regs[4][2] ),
    .Y(_21030_));
 sky130_as_sc_hs__nand3_2 _27536_ (.A(net168),
    .B(_21029_),
    .C(_21030_),
    .Y(_21031_));
 sky130_as_sc_hs__nand3_2 _27537_ (.A(net255),
    .B(_21028_),
    .C(_21031_),
    .Y(_21032_));
 sky130_as_sc_hs__nand3_2 _27538_ (.A(net154),
    .B(_21025_),
    .C(_21032_),
    .Y(_21033_));
 sky130_as_sc_hs__nand3_2 _27539_ (.A(net251),
    .B(_21011_),
    .C(_21018_),
    .Y(_21034_));
 sky130_as_sc_hs__nand3_2 _27540_ (.A(net151),
    .B(_21033_),
    .C(_21034_),
    .Y(_21035_));
 sky130_as_sc_hs__and2_2 _27541_ (.A(_21004_),
    .B(_21035_),
    .Y(_21036_));
 sky130_as_sc_hs__nand3_2 _27546_ (.A(_19754_),
    .B(_21039_),
    .C(_21040_),
    .Y(_21041_));
 sky130_as_sc_hs__nand3_2 _27547_ (.A(_19759_),
    .B(_21038_),
    .C(_21041_),
    .Y(_21042_));
 sky130_as_sc_hs__nand3_2 _27548_ (.A(_20718_),
    .B(_20973_),
    .C(_21042_),
    .Y(_21043_));
 sky130_as_sc_hs__or2_2 _27549_ (.A(net1640),
    .B(_20718_),
    .Y(_21044_));
 sky130_as_sc_hs__and2_2 _27550_ (.A(net500),
    .B(_21043_),
    .Y(_21045_));
 sky130_as_sc_hs__and2_2 _27551_ (.A(net1641),
    .B(_21045_),
    .Y(_00015_));
 sky130_as_sc_hs__and2_2 _27554_ (.A(_21046_),
    .B(_21047_),
    .Y(_21048_));
 sky130_as_sc_hs__and2_2 _27557_ (.A(_21049_),
    .B(_21050_),
    .Y(_21051_));
 sky130_as_sc_hs__and2_2 _27558_ (.A(_21048_),
    .B(_21051_),
    .Y(_21052_));
 sky130_as_sc_hs__and2_2 _27561_ (.A(_21053_),
    .B(_21054_),
    .Y(_21055_));
 sky130_as_sc_hs__nand3_2 _27564_ (.A(_21055_),
    .B(_21056_),
    .C(_21057_),
    .Y(_21058_));
 sky130_as_sc_hs__nor2_2 _27565_ (.A(_20721_),
    .B(_21058_),
    .Y(_21059_));
 sky130_as_sc_hs__and2_2 _27573_ (.A(_21064_),
    .B(_21066_),
    .Y(_21067_));
 sky130_as_sc_hs__nand3_2 _27574_ (.A(_21063_),
    .B(_21065_),
    .C(_21067_),
    .Y(_21068_));
 sky130_as_sc_hs__nor2_2 _27575_ (.A(_21062_),
    .B(_21068_),
    .Y(_21069_));
 sky130_as_sc_hs__nand3_2 _27576_ (.A(_21052_),
    .B(_21059_),
    .C(_21069_),
    .Y(_21070_));
 sky130_as_sc_hs__and2_2 _27579_ (.A(_21071_),
    .B(_21072_),
    .Y(_21073_));
 sky130_as_sc_hs__nand3_2 _27581_ (.A(net137),
    .B(_21070_),
    .C(_21074_),
    .Y(_21075_));
 sky130_as_sc_hs__nand2b_2 _27582_ (.B(net287),
    .Y(_21076_),
    .A(\tholin_riscv.regs[25][3] ));
 sky130_as_sc_hs__or2_2 _27583_ (.A(net287),
    .B(\tholin_riscv.regs[24][3] ),
    .Y(_21077_));
 sky130_as_sc_hs__nand3_2 _27584_ (.A(net167),
    .B(_21076_),
    .C(_21077_),
    .Y(_21078_));
 sky130_as_sc_hs__nand2b_2 _27585_ (.B(net287),
    .Y(_21079_),
    .A(\tholin_riscv.regs[27][3] ));
 sky130_as_sc_hs__or2_2 _27586_ (.A(net287),
    .B(\tholin_riscv.regs[26][3] ),
    .Y(_21080_));
 sky130_as_sc_hs__nand3_2 _27587_ (.A(net264),
    .B(_21079_),
    .C(_21080_),
    .Y(_21081_));
 sky130_as_sc_hs__nand3_2 _27588_ (.A(net157),
    .B(_21078_),
    .C(_21081_),
    .Y(_21082_));
 sky130_as_sc_hs__nand2b_2 _27589_ (.B(net288),
    .Y(_21083_),
    .A(\tholin_riscv.regs[29][3] ));
 sky130_as_sc_hs__or2_2 _27590_ (.A(net288),
    .B(\tholin_riscv.regs[28][3] ),
    .Y(_21084_));
 sky130_as_sc_hs__nand3_2 _27591_ (.A(net167),
    .B(_21083_),
    .C(_21084_),
    .Y(_21085_));
 sky130_as_sc_hs__nand2b_2 _27592_ (.B(net288),
    .Y(_21086_),
    .A(\tholin_riscv.regs[31][3] ));
 sky130_as_sc_hs__or2_2 _27593_ (.A(net288),
    .B(\tholin_riscv.regs[30][3] ),
    .Y(_21087_));
 sky130_as_sc_hs__nand3_2 _27594_ (.A(net264),
    .B(_21086_),
    .C(_21087_),
    .Y(_21088_));
 sky130_as_sc_hs__nand3_2 _27595_ (.A(net256),
    .B(_21085_),
    .C(_21088_),
    .Y(_21089_));
 sky130_as_sc_hs__nand2b_2 _27596_ (.B(net287),
    .Y(_21090_),
    .A(\tholin_riscv.regs[17][3] ));
 sky130_as_sc_hs__or2_2 _27597_ (.A(net287),
    .B(\tholin_riscv.regs[16][3] ),
    .Y(_21091_));
 sky130_as_sc_hs__nand3_2 _27598_ (.A(net173),
    .B(_21090_),
    .C(_21091_),
    .Y(_21092_));
 sky130_as_sc_hs__nand2b_2 _27599_ (.B(net287),
    .Y(_21093_),
    .A(\tholin_riscv.regs[19][3] ));
 sky130_as_sc_hs__or2_2 _27600_ (.A(net287),
    .B(\tholin_riscv.regs[18][3] ),
    .Y(_21094_));
 sky130_as_sc_hs__nand3_2 _27601_ (.A(net264),
    .B(_21093_),
    .C(_21094_),
    .Y(_21095_));
 sky130_as_sc_hs__nand3_2 _27602_ (.A(net157),
    .B(_21092_),
    .C(_21095_),
    .Y(_21096_));
 sky130_as_sc_hs__nand2b_2 _27603_ (.B(net292),
    .Y(_21097_),
    .A(\tholin_riscv.regs[23][3] ));
 sky130_as_sc_hs__or2_2 _27604_ (.A(net292),
    .B(\tholin_riscv.regs[22][3] ),
    .Y(_21098_));
 sky130_as_sc_hs__nand3_2 _27605_ (.A(net282),
    .B(_21097_),
    .C(_21098_),
    .Y(_21099_));
 sky130_as_sc_hs__nand2b_2 _27606_ (.B(net292),
    .Y(_21100_),
    .A(\tholin_riscv.regs[21][3] ));
 sky130_as_sc_hs__or2_2 _27607_ (.A(net292),
    .B(\tholin_riscv.regs[20][3] ),
    .Y(_21101_));
 sky130_as_sc_hs__nand3_2 _27608_ (.A(net173),
    .B(_21100_),
    .C(_21101_),
    .Y(_21102_));
 sky130_as_sc_hs__nand3_2 _27609_ (.A(net256),
    .B(_21099_),
    .C(_21102_),
    .Y(_21103_));
 sky130_as_sc_hs__nand3_2 _27610_ (.A(net153),
    .B(_21096_),
    .C(_21103_),
    .Y(_21104_));
 sky130_as_sc_hs__nand3_2 _27611_ (.A(net250),
    .B(_21082_),
    .C(_21089_),
    .Y(_21105_));
 sky130_as_sc_hs__and2_2 _27612_ (.A(_21104_),
    .B(_21105_),
    .Y(_21106_));
 sky130_as_sc_hs__and2_2 _27613_ (.A(net248),
    .B(_21106_),
    .Y(_21107_));
 sky130_as_sc_hs__nand2b_2 _27614_ (.B(net287),
    .Y(_21108_),
    .A(\tholin_riscv.regs[9][3] ));
 sky130_as_sc_hs__or2_2 _27615_ (.A(net287),
    .B(\tholin_riscv.regs[8][3] ),
    .Y(_21109_));
 sky130_as_sc_hs__nand3_2 _27616_ (.A(net167),
    .B(_21108_),
    .C(_21109_),
    .Y(_21110_));
 sky130_as_sc_hs__nand2b_2 _27617_ (.B(net289),
    .Y(_21111_),
    .A(\tholin_riscv.regs[11][3] ));
 sky130_as_sc_hs__or2_2 _27618_ (.A(net289),
    .B(\tholin_riscv.regs[10][3] ),
    .Y(_21112_));
 sky130_as_sc_hs__nand3_2 _27619_ (.A(net264),
    .B(_21111_),
    .C(_21112_),
    .Y(_21113_));
 sky130_as_sc_hs__nand3_2 _27620_ (.A(net160),
    .B(_21110_),
    .C(_21113_),
    .Y(_21114_));
 sky130_as_sc_hs__nand2b_2 _27621_ (.B(net287),
    .Y(_21115_),
    .A(\tholin_riscv.regs[13][3] ));
 sky130_as_sc_hs__or2_2 _27622_ (.A(net288),
    .B(\tholin_riscv.regs[12][3] ),
    .Y(_21116_));
 sky130_as_sc_hs__nand3_2 _27623_ (.A(net167),
    .B(_21115_),
    .C(_21116_),
    .Y(_21117_));
 sky130_as_sc_hs__nand2b_2 _27624_ (.B(net288),
    .Y(_21118_),
    .A(\tholin_riscv.regs[15][3] ));
 sky130_as_sc_hs__or2_2 _27625_ (.A(net288),
    .B(\tholin_riscv.regs[14][3] ),
    .Y(_21119_));
 sky130_as_sc_hs__nand3_2 _27626_ (.A(net264),
    .B(_21118_),
    .C(_21119_),
    .Y(_21120_));
 sky130_as_sc_hs__nand3_2 _27627_ (.A(net256),
    .B(_21117_),
    .C(_21120_),
    .Y(_21121_));
 sky130_as_sc_hs__nand2b_2 _27628_ (.B(net287),
    .Y(_21122_),
    .A(\tholin_riscv.regs[1][3] ));
 sky130_as_sc_hs__or2_2 _27629_ (.A(net287),
    .B(\tholin_riscv.regs[0][3] ),
    .Y(_21123_));
 sky130_as_sc_hs__nand3_2 _27630_ (.A(net167),
    .B(_21122_),
    .C(_21123_),
    .Y(_21124_));
 sky130_as_sc_hs__nand2b_2 _27631_ (.B(net287),
    .Y(_21125_),
    .A(\tholin_riscv.regs[3][3] ));
 sky130_as_sc_hs__or2_2 _27632_ (.A(net287),
    .B(\tholin_riscv.regs[2][3] ),
    .Y(_21126_));
 sky130_as_sc_hs__nand3_2 _27633_ (.A(net264),
    .B(_21125_),
    .C(_21126_),
    .Y(_21127_));
 sky130_as_sc_hs__nand3_2 _27634_ (.A(net160),
    .B(_21124_),
    .C(_21127_),
    .Y(_21128_));
 sky130_as_sc_hs__nand2b_2 _27635_ (.B(net289),
    .Y(_21129_),
    .A(\tholin_riscv.regs[7][3] ));
 sky130_as_sc_hs__or2_2 _27636_ (.A(net289),
    .B(\tholin_riscv.regs[6][3] ),
    .Y(_21130_));
 sky130_as_sc_hs__nand3_2 _27637_ (.A(net264),
    .B(_21129_),
    .C(_21130_),
    .Y(_21131_));
 sky130_as_sc_hs__nand2b_2 _27638_ (.B(net289),
    .Y(_21132_),
    .A(\tholin_riscv.regs[5][3] ));
 sky130_as_sc_hs__or2_2 _27639_ (.A(net289),
    .B(\tholin_riscv.regs[4][3] ),
    .Y(_21133_));
 sky130_as_sc_hs__nand3_2 _27640_ (.A(net167),
    .B(_21132_),
    .C(_21133_),
    .Y(_21134_));
 sky130_as_sc_hs__nand3_2 _27641_ (.A(net256),
    .B(_21131_),
    .C(_21134_),
    .Y(_21135_));
 sky130_as_sc_hs__nand3_2 _27642_ (.A(net153),
    .B(_21128_),
    .C(_21135_),
    .Y(_21136_));
 sky130_as_sc_hs__nand3_2 _27643_ (.A(net250),
    .B(_21114_),
    .C(_21121_),
    .Y(_21137_));
 sky130_as_sc_hs__and2_2 _27644_ (.A(_21136_),
    .B(_21137_),
    .Y(_21138_));
 sky130_as_sc_hs__and2_2 _27645_ (.A(net151),
    .B(_21138_),
    .Y(_21139_));
 sky130_as_sc_hs__nor2_2 _27646_ (.A(_21107_),
    .B(_21139_),
    .Y(_21140_));
 sky130_as_sc_hs__or2_2 _27647_ (.A(_21107_),
    .B(_21139_),
    .Y(_21141_));
 sky130_as_sc_hs__nand3_2 _27651_ (.A(_19754_),
    .B(_21143_),
    .C(_21144_),
    .Y(_21145_));
 sky130_as_sc_hs__nand3_2 _27652_ (.A(_19759_),
    .B(_21142_),
    .C(_21145_),
    .Y(_21146_));
 sky130_as_sc_hs__nand3_2 _27653_ (.A(_20718_),
    .B(_21075_),
    .C(_21146_),
    .Y(_21147_));
 sky130_as_sc_hs__or2_2 _27654_ (.A(net1628),
    .B(_20718_),
    .Y(_21148_));
 sky130_as_sc_hs__and2_2 _27655_ (.A(net500),
    .B(_21147_),
    .Y(_21149_));
 sky130_as_sc_hs__and2_2 _27656_ (.A(net1629),
    .B(_21149_),
    .Y(_00016_));
 sky130_as_sc_hs__nand3_2 _27660_ (.A(_21150_),
    .B(_21151_),
    .C(_21152_),
    .Y(_21153_));
 sky130_as_sc_hs__and2_2 _27663_ (.A(_21154_),
    .B(_21155_),
    .Y(_21156_));
 sky130_as_sc_hs__nand3_2 _27666_ (.A(_21156_),
    .B(_21157_),
    .C(_21158_),
    .Y(_21159_));
 sky130_as_sc_hs__or2_2 _27667_ (.A(_21153_),
    .B(_21159_),
    .Y(_21160_));
 sky130_as_sc_hs__nor2_2 _27668_ (.A(_20721_),
    .B(_21160_),
    .Y(_21161_));
 sky130_as_sc_hs__nand3_2 _27676_ (.A(_21162_),
    .B(_21165_),
    .C(_21168_),
    .Y(_21169_));
 sky130_as_sc_hs__nand3_2 _27678_ (.A(_19920_),
    .B(_21163_),
    .C(_21166_),
    .Y(_21171_));
 sky130_as_sc_hs__or2_2 _27679_ (.A(_21170_),
    .B(_21171_),
    .Y(_21172_));
 sky130_as_sc_hs__nor2_2 _27680_ (.A(_21169_),
    .B(_21172_),
    .Y(_21173_));
 sky130_as_sc_hs__and2_2 _27684_ (.A(_21175_),
    .B(_21176_),
    .Y(_21177_));
 sky130_as_sc_hs__nand3_2 _27686_ (.A(net137),
    .B(_21174_),
    .C(_21178_),
    .Y(_21179_));
 sky130_as_sc_hs__or2_2 _27688_ (.A(net301),
    .B(\tholin_riscv.regs[24][4] ),
    .Y(_21181_));
 sky130_as_sc_hs__nand3_2 _27689_ (.A(net170),
    .B(_21180_),
    .C(_21181_),
    .Y(_21182_));
 sky130_as_sc_hs__or2_2 _27691_ (.A(net302),
    .B(\tholin_riscv.regs[26][4] ),
    .Y(_21184_));
 sky130_as_sc_hs__nand3_2 _27692_ (.A(net269),
    .B(_21183_),
    .C(_21184_),
    .Y(_21185_));
 sky130_as_sc_hs__nand3_2 _27693_ (.A(net161),
    .B(_21182_),
    .C(_21185_),
    .Y(_21186_));
 sky130_as_sc_hs__or2_2 _27695_ (.A(net302),
    .B(\tholin_riscv.regs[28][4] ),
    .Y(_21188_));
 sky130_as_sc_hs__nand3_2 _27696_ (.A(net170),
    .B(_21187_),
    .C(_21188_),
    .Y(_21189_));
 sky130_as_sc_hs__or2_2 _27698_ (.A(net300),
    .B(\tholin_riscv.regs[30][4] ),
    .Y(_21191_));
 sky130_as_sc_hs__nand3_2 _27699_ (.A(net267),
    .B(_21190_),
    .C(_21191_),
    .Y(_21192_));
 sky130_as_sc_hs__nand3_2 _27700_ (.A(net254),
    .B(_21189_),
    .C(_21192_),
    .Y(_21193_));
 sky130_as_sc_hs__or2_2 _27702_ (.A(net300),
    .B(\tholin_riscv.regs[16][4] ),
    .Y(_21195_));
 sky130_as_sc_hs__nand3_2 _27703_ (.A(net170),
    .B(_21194_),
    .C(_21195_),
    .Y(_21196_));
 sky130_as_sc_hs__or2_2 _27705_ (.A(net300),
    .B(\tholin_riscv.regs[18][4] ),
    .Y(_21198_));
 sky130_as_sc_hs__nand3_2 _27706_ (.A(net267),
    .B(_21197_),
    .C(_21198_),
    .Y(_21199_));
 sky130_as_sc_hs__nand3_2 _27707_ (.A(net161),
    .B(_21196_),
    .C(_21199_),
    .Y(_21200_));
 sky130_as_sc_hs__or2_2 _27709_ (.A(net300),
    .B(\tholin_riscv.regs[22][4] ),
    .Y(_21202_));
 sky130_as_sc_hs__nand3_2 _27710_ (.A(net267),
    .B(_21201_),
    .C(_21202_),
    .Y(_21203_));
 sky130_as_sc_hs__or2_2 _27712_ (.A(net300),
    .B(\tholin_riscv.regs[20][4] ),
    .Y(_21205_));
 sky130_as_sc_hs__nand3_2 _27713_ (.A(net170),
    .B(_21204_),
    .C(_21205_),
    .Y(_21206_));
 sky130_as_sc_hs__nand3_2 _27714_ (.A(net254),
    .B(_21203_),
    .C(_21206_),
    .Y(_21207_));
 sky130_as_sc_hs__nand3_2 _27715_ (.A(net154),
    .B(_21200_),
    .C(_21207_),
    .Y(_21208_));
 sky130_as_sc_hs__nand3_2 _27716_ (.A(net251),
    .B(_21186_),
    .C(_21193_),
    .Y(_21209_));
 sky130_as_sc_hs__nand3_2 _27717_ (.A(net247),
    .B(_21208_),
    .C(_21209_),
    .Y(_21210_));
 sky130_as_sc_hs__or2_2 _27719_ (.A(net302),
    .B(\tholin_riscv.regs[8][4] ),
    .Y(_21212_));
 sky130_as_sc_hs__nand3_2 _27720_ (.A(net170),
    .B(_21211_),
    .C(_21212_),
    .Y(_21213_));
 sky130_as_sc_hs__or2_2 _27722_ (.A(net302),
    .B(\tholin_riscv.regs[10][4] ),
    .Y(_21215_));
 sky130_as_sc_hs__nand3_2 _27723_ (.A(net269),
    .B(_21214_),
    .C(_21215_),
    .Y(_21216_));
 sky130_as_sc_hs__nand3_2 _27724_ (.A(net161),
    .B(_21213_),
    .C(_21216_),
    .Y(_21217_));
 sky130_as_sc_hs__or2_2 _27726_ (.A(net302),
    .B(\tholin_riscv.regs[12][4] ),
    .Y(_21219_));
 sky130_as_sc_hs__nand3_2 _27727_ (.A(net170),
    .B(_21218_),
    .C(_21219_),
    .Y(_21220_));
 sky130_as_sc_hs__or2_2 _27729_ (.A(net302),
    .B(\tholin_riscv.regs[14][4] ),
    .Y(_21222_));
 sky130_as_sc_hs__nand3_2 _27730_ (.A(net269),
    .B(_21221_),
    .C(_21222_),
    .Y(_21223_));
 sky130_as_sc_hs__nand3_2 _27731_ (.A(net254),
    .B(_21220_),
    .C(_21223_),
    .Y(_21224_));
 sky130_as_sc_hs__or2_2 _27733_ (.A(net301),
    .B(\tholin_riscv.regs[0][4] ),
    .Y(_21226_));
 sky130_as_sc_hs__nand3_2 _27734_ (.A(net170),
    .B(_21225_),
    .C(_21226_),
    .Y(_21227_));
 sky130_as_sc_hs__or2_2 _27736_ (.A(net322),
    .B(\tholin_riscv.regs[2][4] ),
    .Y(_21229_));
 sky130_as_sc_hs__nand3_2 _27737_ (.A(net267),
    .B(_21228_),
    .C(_21229_),
    .Y(_21230_));
 sky130_as_sc_hs__nand3_2 _27738_ (.A(net161),
    .B(_21227_),
    .C(_21230_),
    .Y(_21231_));
 sky130_as_sc_hs__or2_2 _27740_ (.A(net302),
    .B(\tholin_riscv.regs[6][4] ),
    .Y(_21233_));
 sky130_as_sc_hs__nand3_2 _27741_ (.A(net267),
    .B(_21232_),
    .C(_21233_),
    .Y(_21234_));
 sky130_as_sc_hs__or2_2 _27743_ (.A(net302),
    .B(\tholin_riscv.regs[4][4] ),
    .Y(_21236_));
 sky130_as_sc_hs__nand3_2 _27744_ (.A(net172),
    .B(_21235_),
    .C(_21236_),
    .Y(_21237_));
 sky130_as_sc_hs__nand3_2 _27745_ (.A(net254),
    .B(_21234_),
    .C(_21237_),
    .Y(_21238_));
 sky130_as_sc_hs__nand3_2 _27746_ (.A(net154),
    .B(_21231_),
    .C(_21238_),
    .Y(_21239_));
 sky130_as_sc_hs__nand3_2 _27747_ (.A(net251),
    .B(_21217_),
    .C(_21224_),
    .Y(_21240_));
 sky130_as_sc_hs__nand3_2 _27748_ (.A(net151),
    .B(_21239_),
    .C(_21240_),
    .Y(_21241_));
 sky130_as_sc_hs__nand3_2 _27753_ (.A(_19754_),
    .B(_21244_),
    .C(_21245_),
    .Y(_21246_));
 sky130_as_sc_hs__nand3_2 _27754_ (.A(_19759_),
    .B(_21243_),
    .C(_21246_),
    .Y(_21247_));
 sky130_as_sc_hs__nand3_2 _27755_ (.A(_20718_),
    .B(_21179_),
    .C(_21247_),
    .Y(_21248_));
 sky130_as_sc_hs__or2_2 _27756_ (.A(net1634),
    .B(_20718_),
    .Y(_21249_));
 sky130_as_sc_hs__and2_2 _27757_ (.A(net500),
    .B(_21248_),
    .Y(_21250_));
 sky130_as_sc_hs__and2_2 _27758_ (.A(net1635),
    .B(_21250_),
    .Y(_00017_));
 sky130_as_sc_hs__and2_2 _27761_ (.A(_21251_),
    .B(_21252_),
    .Y(_21253_));
 sky130_as_sc_hs__and2_2 _27764_ (.A(_21254_),
    .B(_21255_),
    .Y(_21256_));
 sky130_as_sc_hs__and2_2 _27765_ (.A(_21253_),
    .B(_21256_),
    .Y(_21257_));
 sky130_as_sc_hs__and2_2 _27768_ (.A(_21258_),
    .B(_21259_),
    .Y(_21260_));
 sky130_as_sc_hs__nand3_2 _27771_ (.A(_21260_),
    .B(_21261_),
    .C(_21262_),
    .Y(_21263_));
 sky130_as_sc_hs__nor2_2 _27772_ (.A(_20721_),
    .B(_21263_),
    .Y(_21264_));
 sky130_as_sc_hs__and2_2 _27780_ (.A(_21269_),
    .B(_21271_),
    .Y(_21272_));
 sky130_as_sc_hs__nand3_2 _27781_ (.A(_21268_),
    .B(_21270_),
    .C(_21272_),
    .Y(_21273_));
 sky130_as_sc_hs__nor2_2 _27782_ (.A(_21267_),
    .B(_21273_),
    .Y(_21274_));
 sky130_as_sc_hs__nand3_2 _27783_ (.A(_21257_),
    .B(_21264_),
    .C(_21274_),
    .Y(_21275_));
 sky130_as_sc_hs__and2_2 _27786_ (.A(_21276_),
    .B(_21277_),
    .Y(_21278_));
 sky130_as_sc_hs__nand3_2 _27788_ (.A(_19758_),
    .B(_21275_),
    .C(_21279_),
    .Y(_21280_));
 sky130_as_sc_hs__nand2b_2 _27789_ (.B(net289),
    .Y(_21281_),
    .A(\tholin_riscv.regs[25][5] ));
 sky130_as_sc_hs__or2_2 _27790_ (.A(net289),
    .B(\tholin_riscv.regs[24][5] ),
    .Y(_21282_));
 sky130_as_sc_hs__nand3_2 _27791_ (.A(net167),
    .B(_21281_),
    .C(_21282_),
    .Y(_21283_));
 sky130_as_sc_hs__nand2b_2 _27792_ (.B(net312),
    .Y(_21284_),
    .A(\tholin_riscv.regs[27][5] ));
 sky130_as_sc_hs__or2_2 _27793_ (.A(net312),
    .B(\tholin_riscv.regs[26][5] ),
    .Y(_21285_));
 sky130_as_sc_hs__nand3_2 _27794_ (.A(net264),
    .B(_21284_),
    .C(_21285_),
    .Y(_21286_));
 sky130_as_sc_hs__nand3_2 _27795_ (.A(net157),
    .B(_21283_),
    .C(_21286_),
    .Y(_21287_));
 sky130_as_sc_hs__nand2b_2 _27796_ (.B(net289),
    .Y(_21288_),
    .A(\tholin_riscv.regs[29][5] ));
 sky130_as_sc_hs__or2_2 _27797_ (.A(net289),
    .B(\tholin_riscv.regs[28][5] ),
    .Y(_21289_));
 sky130_as_sc_hs__nand3_2 _27798_ (.A(net167),
    .B(_21288_),
    .C(_21289_),
    .Y(_21290_));
 sky130_as_sc_hs__nand2b_2 _27799_ (.B(net289),
    .Y(_21291_),
    .A(\tholin_riscv.regs[31][5] ));
 sky130_as_sc_hs__or2_2 _27800_ (.A(net289),
    .B(\tholin_riscv.regs[30][5] ),
    .Y(_21292_));
 sky130_as_sc_hs__nand3_2 _27801_ (.A(net264),
    .B(_21291_),
    .C(_21292_),
    .Y(_21293_));
 sky130_as_sc_hs__nand3_2 _27802_ (.A(net256),
    .B(_21290_),
    .C(_21293_),
    .Y(_21294_));
 sky130_as_sc_hs__nand2b_2 _27803_ (.B(net290),
    .Y(_21295_),
    .A(\tholin_riscv.regs[17][5] ));
 sky130_as_sc_hs__or2_2 _27804_ (.A(net290),
    .B(\tholin_riscv.regs[16][5] ),
    .Y(_21296_));
 sky130_as_sc_hs__nand3_2 _27805_ (.A(net167),
    .B(_21295_),
    .C(_21296_),
    .Y(_21297_));
 sky130_as_sc_hs__nand2b_2 _27806_ (.B(net289),
    .Y(_21298_),
    .A(\tholin_riscv.regs[19][5] ));
 sky130_as_sc_hs__or2_2 _27807_ (.A(net289),
    .B(\tholin_riscv.regs[18][5] ),
    .Y(_21299_));
 sky130_as_sc_hs__nand3_2 _27808_ (.A(net264),
    .B(_21298_),
    .C(_21299_),
    .Y(_21300_));
 sky130_as_sc_hs__nand3_2 _27809_ (.A(net157),
    .B(_21297_),
    .C(_21300_),
    .Y(_21301_));
 sky130_as_sc_hs__nand2b_2 _27810_ (.B(net290),
    .Y(_21302_),
    .A(\tholin_riscv.regs[23][5] ));
 sky130_as_sc_hs__or2_2 _27811_ (.A(net290),
    .B(\tholin_riscv.regs[22][5] ),
    .Y(_21303_));
 sky130_as_sc_hs__nand3_2 _27812_ (.A(net264),
    .B(_21302_),
    .C(_21303_),
    .Y(_21304_));
 sky130_as_sc_hs__nand2b_2 _27813_ (.B(net290),
    .Y(_21305_),
    .A(\tholin_riscv.regs[21][5] ));
 sky130_as_sc_hs__or2_2 _27814_ (.A(net290),
    .B(\tholin_riscv.regs[20][5] ),
    .Y(_21306_));
 sky130_as_sc_hs__nand3_2 _27815_ (.A(net167),
    .B(_21305_),
    .C(_21306_),
    .Y(_21307_));
 sky130_as_sc_hs__nand3_2 _27816_ (.A(net256),
    .B(_21304_),
    .C(_21307_),
    .Y(_21308_));
 sky130_as_sc_hs__nand3_2 _27817_ (.A(net153),
    .B(_21301_),
    .C(_21308_),
    .Y(_21309_));
 sky130_as_sc_hs__nand3_2 _27818_ (.A(net250),
    .B(_21287_),
    .C(_21294_),
    .Y(_21310_));
 sky130_as_sc_hs__nand3_2 _27819_ (.A(net248),
    .B(_21309_),
    .C(_21310_),
    .Y(_21311_));
 sky130_as_sc_hs__nand2b_2 _27820_ (.B(net321),
    .Y(_21312_),
    .A(\tholin_riscv.regs[9][5] ));
 sky130_as_sc_hs__or2_2 _27821_ (.A(net321),
    .B(\tholin_riscv.regs[8][5] ),
    .Y(_21313_));
 sky130_as_sc_hs__nand3_2 _27822_ (.A(net172),
    .B(_21312_),
    .C(_21313_),
    .Y(_21314_));
 sky130_as_sc_hs__nand2b_2 _27823_ (.B(net321),
    .Y(_21315_),
    .A(\tholin_riscv.regs[11][5] ));
 sky130_as_sc_hs__or2_2 _27824_ (.A(net321),
    .B(\tholin_riscv.regs[10][5] ),
    .Y(_21316_));
 sky130_as_sc_hs__nand3_2 _27825_ (.A(net277),
    .B(_21315_),
    .C(_21316_),
    .Y(_21317_));
 sky130_as_sc_hs__nand3_2 _27826_ (.A(net161),
    .B(_21314_),
    .C(_21317_),
    .Y(_21318_));
 sky130_as_sc_hs__nand2b_2 _27827_ (.B(net321),
    .Y(_21319_),
    .A(\tholin_riscv.regs[13][5] ));
 sky130_as_sc_hs__or2_2 _27828_ (.A(net312),
    .B(\tholin_riscv.regs[12][5] ),
    .Y(_21320_));
 sky130_as_sc_hs__nand3_2 _27829_ (.A(net182),
    .B(_21319_),
    .C(_21320_),
    .Y(_21321_));
 sky130_as_sc_hs__nand2b_2 _27830_ (.B(net321),
    .Y(_21322_),
    .A(\tholin_riscv.regs[15][5] ));
 sky130_as_sc_hs__or2_2 _27831_ (.A(net321),
    .B(\tholin_riscv.regs[14][5] ),
    .Y(_21323_));
 sky130_as_sc_hs__nand3_2 _27832_ (.A(net277),
    .B(_21322_),
    .C(_21323_),
    .Y(_21324_));
 sky130_as_sc_hs__nand3_2 _27833_ (.A(net260),
    .B(_21321_),
    .C(_21324_),
    .Y(_21325_));
 sky130_as_sc_hs__nand2b_2 _27834_ (.B(net290),
    .Y(_21326_),
    .A(\tholin_riscv.regs[1][5] ));
 sky130_as_sc_hs__or2_2 _27835_ (.A(net290),
    .B(\tholin_riscv.regs[0][5] ),
    .Y(_21327_));
 sky130_as_sc_hs__nand3_2 _27836_ (.A(net172),
    .B(_21326_),
    .C(_21327_),
    .Y(_21328_));
 sky130_as_sc_hs__nand2b_2 _27837_ (.B(net301),
    .Y(_21329_),
    .A(\tholin_riscv.regs[3][5] ));
 sky130_as_sc_hs__or2_2 _27838_ (.A(net301),
    .B(\tholin_riscv.regs[2][5] ),
    .Y(_21330_));
 sky130_as_sc_hs__nand3_2 _27839_ (.A(net269),
    .B(_21329_),
    .C(_21330_),
    .Y(_21331_));
 sky130_as_sc_hs__nand3_2 _27840_ (.A(net165),
    .B(_21328_),
    .C(_21331_),
    .Y(_21332_));
 sky130_as_sc_hs__nand2b_2 _27841_ (.B(net312),
    .Y(_21333_),
    .A(\tholin_riscv.regs[7][5] ));
 sky130_as_sc_hs__or2_2 _27842_ (.A(net312),
    .B(\tholin_riscv.regs[6][5] ),
    .Y(_21334_));
 sky130_as_sc_hs__nand3_2 _27843_ (.A(net271),
    .B(_21333_),
    .C(_21334_),
    .Y(_21335_));
 sky130_as_sc_hs__nand2b_2 _27844_ (.B(net312),
    .Y(_21336_),
    .A(\tholin_riscv.regs[5][5] ));
 sky130_as_sc_hs__or2_2 _27845_ (.A(net312),
    .B(\tholin_riscv.regs[4][5] ),
    .Y(_21337_));
 sky130_as_sc_hs__nand3_2 _27846_ (.A(net175),
    .B(_21336_),
    .C(_21337_),
    .Y(_21338_));
 sky130_as_sc_hs__nand3_2 _27847_ (.A(net257),
    .B(_21335_),
    .C(_21338_),
    .Y(_21339_));
 sky130_as_sc_hs__nand3_2 _27848_ (.A(net154),
    .B(_21332_),
    .C(_21339_),
    .Y(_21340_));
 sky130_as_sc_hs__nand3_2 _27849_ (.A(net251),
    .B(_21318_),
    .C(_21325_),
    .Y(_21341_));
 sky130_as_sc_hs__nand3_2 _27850_ (.A(net151),
    .B(_21340_),
    .C(_21341_),
    .Y(_21342_));
 sky130_as_sc_hs__and2_2 _27851_ (.A(_21311_),
    .B(_21342_),
    .Y(_21343_));
 sky130_as_sc_hs__nand3_2 _27856_ (.A(_19754_),
    .B(_21346_),
    .C(_21347_),
    .Y(_21348_));
 sky130_as_sc_hs__nand3_2 _27857_ (.A(_19759_),
    .B(_21345_),
    .C(_21348_),
    .Y(_21349_));
 sky130_as_sc_hs__nand3_2 _27858_ (.A(_20718_),
    .B(_21280_),
    .C(_21349_),
    .Y(_21350_));
 sky130_as_sc_hs__or2_2 _27859_ (.A(net1654),
    .B(_20718_),
    .Y(_21351_));
 sky130_as_sc_hs__and2_2 _27860_ (.A(net500),
    .B(_21350_),
    .Y(_21352_));
 sky130_as_sc_hs__and2_2 _27861_ (.A(_21351_),
    .B(_21352_),
    .Y(_00018_));
 sky130_as_sc_hs__and2_2 _27869_ (.A(_21358_),
    .B(_21359_),
    .Y(_21360_));
 sky130_as_sc_hs__nand3_2 _27870_ (.A(_21356_),
    .B(_21357_),
    .C(_21360_),
    .Y(_21361_));
 sky130_as_sc_hs__nor2_2 _27871_ (.A(_20721_),
    .B(_21361_),
    .Y(_21362_));
 sky130_as_sc_hs__and2_2 _27876_ (.A(_21353_),
    .B(_21355_),
    .Y(_21367_));
 sky130_as_sc_hs__and2_2 _27877_ (.A(_21366_),
    .B(_21367_),
    .Y(_21368_));
 sky130_as_sc_hs__nand3_2 _27879_ (.A(_19998_),
    .B(_21364_),
    .C(_21365_),
    .Y(_21370_));
 sky130_as_sc_hs__nor2_2 _27880_ (.A(_21369_),
    .B(_21370_),
    .Y(_21371_));
 sky130_as_sc_hs__nand3_2 _27881_ (.A(_21362_),
    .B(_21368_),
    .C(_21371_),
    .Y(_21372_));
 sky130_as_sc_hs__and2_2 _27884_ (.A(_21373_),
    .B(_21374_),
    .Y(_21375_));
 sky130_as_sc_hs__nand3_2 _27886_ (.A(_19758_),
    .B(_21372_),
    .C(_21376_),
    .Y(_21377_));
 sky130_as_sc_hs__nand2b_2 _27887_ (.B(net299),
    .Y(_21378_),
    .A(\tholin_riscv.regs[25][6] ));
 sky130_as_sc_hs__or2_2 _27888_ (.A(net288),
    .B(\tholin_riscv.regs[24][6] ),
    .Y(_21379_));
 sky130_as_sc_hs__nand3_2 _27889_ (.A(net170),
    .B(_21378_),
    .C(_21379_),
    .Y(_21380_));
 sky130_as_sc_hs__nand2b_2 _27890_ (.B(net299),
    .Y(_21381_),
    .A(\tholin_riscv.regs[27][6] ));
 sky130_as_sc_hs__or2_2 _27891_ (.A(net299),
    .B(\tholin_riscv.regs[26][6] ),
    .Y(_21382_));
 sky130_as_sc_hs__nand3_2 _27892_ (.A(net267),
    .B(_21381_),
    .C(_21382_),
    .Y(_21383_));
 sky130_as_sc_hs__nand3_2 _27893_ (.A(net161),
    .B(_21380_),
    .C(_21383_),
    .Y(_21384_));
 sky130_as_sc_hs__nand2b_2 _27894_ (.B(net299),
    .Y(_21385_),
    .A(\tholin_riscv.regs[29][6] ));
 sky130_as_sc_hs__or2_2 _27895_ (.A(net299),
    .B(\tholin_riscv.regs[28][6] ),
    .Y(_21386_));
 sky130_as_sc_hs__nand3_2 _27896_ (.A(net170),
    .B(_21385_),
    .C(_21386_),
    .Y(_21387_));
 sky130_as_sc_hs__nand2b_2 _27897_ (.B(net299),
    .Y(_21388_),
    .A(\tholin_riscv.regs[31][6] ));
 sky130_as_sc_hs__or2_2 _27898_ (.A(net299),
    .B(\tholin_riscv.regs[30][6] ),
    .Y(_21389_));
 sky130_as_sc_hs__nand3_2 _27899_ (.A(net267),
    .B(_21388_),
    .C(_21389_),
    .Y(_21390_));
 sky130_as_sc_hs__nand3_2 _27900_ (.A(net254),
    .B(_21387_),
    .C(_21390_),
    .Y(_21391_));
 sky130_as_sc_hs__nand2b_2 _27901_ (.B(net288),
    .Y(_21392_),
    .A(\tholin_riscv.regs[17][6] ));
 sky130_as_sc_hs__or2_2 _27902_ (.A(net288),
    .B(\tholin_riscv.regs[16][6] ),
    .Y(_21393_));
 sky130_as_sc_hs__nand3_2 _27903_ (.A(net167),
    .B(_21392_),
    .C(_21393_),
    .Y(_21394_));
 sky130_as_sc_hs__nand2b_2 _27904_ (.B(net289),
    .Y(_21395_),
    .A(\tholin_riscv.regs[19][6] ));
 sky130_as_sc_hs__or2_2 _27905_ (.A(net290),
    .B(\tholin_riscv.regs[18][6] ),
    .Y(_21396_));
 sky130_as_sc_hs__nand3_2 _27906_ (.A(net264),
    .B(_21395_),
    .C(_21396_),
    .Y(_21397_));
 sky130_as_sc_hs__nand3_2 _27907_ (.A(net157),
    .B(_21394_),
    .C(_21397_),
    .Y(_21398_));
 sky130_as_sc_hs__nand2b_2 _27908_ (.B(net301),
    .Y(_21399_),
    .A(\tholin_riscv.regs[23][6] ));
 sky130_as_sc_hs__or2_2 _27909_ (.A(net301),
    .B(\tholin_riscv.regs[22][6] ),
    .Y(_21400_));
 sky130_as_sc_hs__nand3_2 _27910_ (.A(net267),
    .B(_21399_),
    .C(_21400_),
    .Y(_21401_));
 sky130_as_sc_hs__nand2b_2 _27911_ (.B(net301),
    .Y(_21402_),
    .A(\tholin_riscv.regs[21][6] ));
 sky130_as_sc_hs__or2_2 _27912_ (.A(net301),
    .B(\tholin_riscv.regs[20][6] ),
    .Y(_21403_));
 sky130_as_sc_hs__nand3_2 _27913_ (.A(net170),
    .B(_21402_),
    .C(_21403_),
    .Y(_21404_));
 sky130_as_sc_hs__nand3_2 _27914_ (.A(net254),
    .B(_21401_),
    .C(_21404_),
    .Y(_21405_));
 sky130_as_sc_hs__nand3_2 _27915_ (.A(net154),
    .B(_21398_),
    .C(_21405_),
    .Y(_21406_));
 sky130_as_sc_hs__nand3_2 _27916_ (.A(net251),
    .B(_21384_),
    .C(_21391_),
    .Y(_21407_));
 sky130_as_sc_hs__nand3_2 _27917_ (.A(net247),
    .B(_21406_),
    .C(_21407_),
    .Y(_21408_));
 sky130_as_sc_hs__nand2b_2 _27918_ (.B(net299),
    .Y(_21409_),
    .A(\tholin_riscv.regs[9][6] ));
 sky130_as_sc_hs__or2_2 _27919_ (.A(net299),
    .B(\tholin_riscv.regs[8][6] ),
    .Y(_21410_));
 sky130_as_sc_hs__nand3_2 _27920_ (.A(net170),
    .B(_21409_),
    .C(_21410_),
    .Y(_21411_));
 sky130_as_sc_hs__nand2b_2 _27921_ (.B(net299),
    .Y(_21412_),
    .A(\tholin_riscv.regs[11][6] ));
 sky130_as_sc_hs__or2_2 _27922_ (.A(net299),
    .B(\tholin_riscv.regs[10][6] ),
    .Y(_21413_));
 sky130_as_sc_hs__nand3_2 _27923_ (.A(net267),
    .B(_21412_),
    .C(_21413_),
    .Y(_21414_));
 sky130_as_sc_hs__nand3_2 _27924_ (.A(net161),
    .B(_21411_),
    .C(_21414_),
    .Y(_21415_));
 sky130_as_sc_hs__nand2b_2 _27925_ (.B(net301),
    .Y(_21416_),
    .A(\tholin_riscv.regs[13][6] ));
 sky130_as_sc_hs__or2_2 _27926_ (.A(net301),
    .B(\tholin_riscv.regs[12][6] ),
    .Y(_21417_));
 sky130_as_sc_hs__nand3_2 _27927_ (.A(net170),
    .B(_21416_),
    .C(_21417_),
    .Y(_21418_));
 sky130_as_sc_hs__nand2b_2 _27928_ (.B(net302),
    .Y(_21419_),
    .A(\tholin_riscv.regs[15][6] ));
 sky130_as_sc_hs__or2_2 _27929_ (.A(net302),
    .B(\tholin_riscv.regs[14][6] ),
    .Y(_21420_));
 sky130_as_sc_hs__nand3_2 _27930_ (.A(net267),
    .B(_21419_),
    .C(_21420_),
    .Y(_21421_));
 sky130_as_sc_hs__nand3_2 _27931_ (.A(net254),
    .B(_21418_),
    .C(_21421_),
    .Y(_21422_));
 sky130_as_sc_hs__nand2b_2 _27932_ (.B(net301),
    .Y(_21423_),
    .A(\tholin_riscv.regs[1][6] ));
 sky130_as_sc_hs__or2_2 _27933_ (.A(net301),
    .B(\tholin_riscv.regs[0][6] ),
    .Y(_21424_));
 sky130_as_sc_hs__nand3_2 _27934_ (.A(net170),
    .B(_21423_),
    .C(_21424_),
    .Y(_21425_));
 sky130_as_sc_hs__nand2b_2 _27935_ (.B(net301),
    .Y(_21426_),
    .A(\tholin_riscv.regs[3][6] ));
 sky130_as_sc_hs__or2_2 _27936_ (.A(net301),
    .B(\tholin_riscv.regs[2][6] ),
    .Y(_21427_));
 sky130_as_sc_hs__nand3_2 _27937_ (.A(net267),
    .B(_21426_),
    .C(_21427_),
    .Y(_21428_));
 sky130_as_sc_hs__nand3_2 _27938_ (.A(net161),
    .B(_21425_),
    .C(_21428_),
    .Y(_21429_));
 sky130_as_sc_hs__nand2b_2 _27939_ (.B(net301),
    .Y(_21430_),
    .A(\tholin_riscv.regs[7][6] ));
 sky130_as_sc_hs__or2_2 _27940_ (.A(net301),
    .B(\tholin_riscv.regs[6][6] ),
    .Y(_21431_));
 sky130_as_sc_hs__nand3_2 _27941_ (.A(net267),
    .B(_21430_),
    .C(_21431_),
    .Y(_21432_));
 sky130_as_sc_hs__nand2b_2 _27942_ (.B(net321),
    .Y(_21433_),
    .A(\tholin_riscv.regs[5][6] ));
 sky130_as_sc_hs__or2_2 _27943_ (.A(net321),
    .B(\tholin_riscv.regs[4][6] ),
    .Y(_21434_));
 sky130_as_sc_hs__nand3_2 _27944_ (.A(net170),
    .B(_21433_),
    .C(_21434_),
    .Y(_21435_));
 sky130_as_sc_hs__nand3_2 _27945_ (.A(net254),
    .B(_21432_),
    .C(_21435_),
    .Y(_21436_));
 sky130_as_sc_hs__nand3_2 _27946_ (.A(net154),
    .B(_21429_),
    .C(_21436_),
    .Y(_21437_));
 sky130_as_sc_hs__nand3_2 _27947_ (.A(net251),
    .B(_21415_),
    .C(_21422_),
    .Y(_21438_));
 sky130_as_sc_hs__nand3_2 _27948_ (.A(net151),
    .B(_21437_),
    .C(_21438_),
    .Y(_21439_));
 sky130_as_sc_hs__and2_2 _27949_ (.A(_21408_),
    .B(_21439_),
    .Y(_21440_));
 sky130_as_sc_hs__or2_2 _27950_ (.A(_19754_),
    .B(_21440_),
    .Y(_21441_));
 sky130_as_sc_hs__nand3_2 _27953_ (.A(_19754_),
    .B(_21442_),
    .C(_21443_),
    .Y(_21444_));
 sky130_as_sc_hs__nand3_2 _27954_ (.A(_19759_),
    .B(_21441_),
    .C(_21444_),
    .Y(_21445_));
 sky130_as_sc_hs__nand3_2 _27955_ (.A(_20718_),
    .B(_21377_),
    .C(_21445_),
    .Y(_21446_));
 sky130_as_sc_hs__or2_2 _27956_ (.A(net1428),
    .B(_20718_),
    .Y(_21447_));
 sky130_as_sc_hs__and2_2 _27957_ (.A(net502),
    .B(_21446_),
    .Y(_21448_));
 sky130_as_sc_hs__and2_2 _27958_ (.A(net1429),
    .B(_21448_),
    .Y(_00019_));
 sky130_as_sc_hs__nand3_2 _27965_ (.A(_21452_),
    .B(_21453_),
    .C(_21454_),
    .Y(_21455_));
 sky130_as_sc_hs__nor2_2 _27966_ (.A(_20721_),
    .B(_21455_),
    .Y(_21456_));
 sky130_as_sc_hs__and2_2 _27972_ (.A(_21451_),
    .B(_21460_),
    .Y(_21462_));
 sky130_as_sc_hs__and2_2 _27973_ (.A(_21461_),
    .B(_21462_),
    .Y(_21463_));
 sky130_as_sc_hs__nand3_2 _27974_ (.A(_21449_),
    .B(_21458_),
    .C(_21459_),
    .Y(_21464_));
 sky130_as_sc_hs__nor2_2 _27976_ (.A(_21464_),
    .B(_21465_),
    .Y(_21466_));
 sky130_as_sc_hs__nand3_2 _27977_ (.A(_21456_),
    .B(_21463_),
    .C(_21466_),
    .Y(_21467_));
 sky130_as_sc_hs__nand3_2 _27980_ (.A(_20721_),
    .B(_21468_),
    .C(_21469_),
    .Y(_21470_));
 sky130_as_sc_hs__nand3_2 _27981_ (.A(_19758_),
    .B(_21467_),
    .C(_21470_),
    .Y(_21471_));
 sky130_as_sc_hs__or2_2 _27982_ (.A(net188),
    .B(\tholin_riscv.regs[25][7] ),
    .Y(_21472_));
 sky130_as_sc_hs__or2_2 _27983_ (.A(net312),
    .B(\tholin_riscv.regs[24][7] ),
    .Y(_21473_));
 sky130_as_sc_hs__nand3_2 _27984_ (.A(net167),
    .B(_21472_),
    .C(_21473_),
    .Y(_21474_));
 sky130_as_sc_hs__or2_2 _27985_ (.A(net188),
    .B(\tholin_riscv.regs[27][7] ),
    .Y(_21475_));
 sky130_as_sc_hs__or2_2 _27986_ (.A(net312),
    .B(\tholin_riscv.regs[26][7] ),
    .Y(_21476_));
 sky130_as_sc_hs__nand3_2 _27987_ (.A(net271),
    .B(_21475_),
    .C(_21476_),
    .Y(_21477_));
 sky130_as_sc_hs__nand3_2 _27988_ (.A(net160),
    .B(_21474_),
    .C(_21477_),
    .Y(_21478_));
 sky130_as_sc_hs__or2_2 _27989_ (.A(net188),
    .B(\tholin_riscv.regs[29][7] ),
    .Y(_21479_));
 sky130_as_sc_hs__or2_2 _27990_ (.A(net308),
    .B(\tholin_riscv.regs[28][7] ),
    .Y(_21480_));
 sky130_as_sc_hs__nand3_2 _27991_ (.A(net174),
    .B(_21479_),
    .C(_21480_),
    .Y(_21481_));
 sky130_as_sc_hs__or2_2 _27992_ (.A(net188),
    .B(\tholin_riscv.regs[31][7] ),
    .Y(_21482_));
 sky130_as_sc_hs__or2_2 _27993_ (.A(net312),
    .B(\tholin_riscv.regs[30][7] ),
    .Y(_21483_));
 sky130_as_sc_hs__nand3_2 _27994_ (.A(net271),
    .B(_21482_),
    .C(_21483_),
    .Y(_21484_));
 sky130_as_sc_hs__nand3_2 _27995_ (.A(net257),
    .B(_21481_),
    .C(_21484_),
    .Y(_21485_));
 sky130_as_sc_hs__or2_2 _27996_ (.A(net187),
    .B(\tholin_riscv.regs[17][7] ),
    .Y(_21486_));
 sky130_as_sc_hs__or2_2 _27997_ (.A(net286),
    .B(\tholin_riscv.regs[16][7] ),
    .Y(_21487_));
 sky130_as_sc_hs__nand3_2 _27998_ (.A(net167),
    .B(_21486_),
    .C(_21487_),
    .Y(_21488_));
 sky130_as_sc_hs__or2_2 _27999_ (.A(net188),
    .B(\tholin_riscv.regs[19][7] ),
    .Y(_21489_));
 sky130_as_sc_hs__or2_2 _28000_ (.A(net289),
    .B(\tholin_riscv.regs[18][7] ),
    .Y(_21490_));
 sky130_as_sc_hs__nand3_2 _28001_ (.A(net264),
    .B(_21489_),
    .C(_21490_),
    .Y(_21491_));
 sky130_as_sc_hs__nand3_2 _28002_ (.A(net157),
    .B(_21488_),
    .C(_21491_),
    .Y(_21492_));
 sky130_as_sc_hs__or2_2 _28003_ (.A(net187),
    .B(\tholin_riscv.regs[23][7] ),
    .Y(_21493_));
 sky130_as_sc_hs__or2_2 _28004_ (.A(net311),
    .B(\tholin_riscv.regs[22][7] ),
    .Y(_21494_));
 sky130_as_sc_hs__nand3_2 _28005_ (.A(net270),
    .B(_21493_),
    .C(_21494_),
    .Y(_21495_));
 sky130_as_sc_hs__or2_2 _28006_ (.A(net187),
    .B(\tholin_riscv.regs[21][7] ),
    .Y(_21496_));
 sky130_as_sc_hs__or2_2 _28007_ (.A(net311),
    .B(\tholin_riscv.regs[20][7] ),
    .Y(_21497_));
 sky130_as_sc_hs__nand3_2 _28008_ (.A(net174),
    .B(_21496_),
    .C(_21497_),
    .Y(_21498_));
 sky130_as_sc_hs__nand3_2 _28009_ (.A(net257),
    .B(_21495_),
    .C(_21498_),
    .Y(_21499_));
 sky130_as_sc_hs__nand3_2 _28010_ (.A(net153),
    .B(_21492_),
    .C(_21499_),
    .Y(_21500_));
 sky130_as_sc_hs__nand3_2 _28011_ (.A(net250),
    .B(_21478_),
    .C(_21485_),
    .Y(_21501_));
 sky130_as_sc_hs__nand3_2 _28012_ (.A(net248),
    .B(_21500_),
    .C(_21501_),
    .Y(_21502_));
 sky130_as_sc_hs__or2_2 _28013_ (.A(net188),
    .B(\tholin_riscv.regs[9][7] ),
    .Y(_21503_));
 sky130_as_sc_hs__or2_2 _28014_ (.A(net312),
    .B(\tholin_riscv.regs[8][7] ),
    .Y(_21504_));
 sky130_as_sc_hs__nand3_2 _28015_ (.A(net175),
    .B(_21503_),
    .C(_21504_),
    .Y(_21505_));
 sky130_as_sc_hs__or2_2 _28016_ (.A(net188),
    .B(\tholin_riscv.regs[11][7] ),
    .Y(_21506_));
 sky130_as_sc_hs__or2_2 _28017_ (.A(net313),
    .B(\tholin_riscv.regs[10][7] ),
    .Y(_21507_));
 sky130_as_sc_hs__nand3_2 _28018_ (.A(net271),
    .B(_21506_),
    .C(_21507_),
    .Y(_21508_));
 sky130_as_sc_hs__nand3_2 _28019_ (.A(net159),
    .B(_21505_),
    .C(_21508_),
    .Y(_21509_));
 sky130_as_sc_hs__or2_2 _28020_ (.A(net189),
    .B(\tholin_riscv.regs[13][7] ),
    .Y(_21510_));
 sky130_as_sc_hs__or2_2 _28021_ (.A(net313),
    .B(\tholin_riscv.regs[12][7] ),
    .Y(_21511_));
 sky130_as_sc_hs__nand3_2 _28022_ (.A(net175),
    .B(_21510_),
    .C(_21511_),
    .Y(_21512_));
 sky130_as_sc_hs__or2_2 _28023_ (.A(net188),
    .B(\tholin_riscv.regs[15][7] ),
    .Y(_21513_));
 sky130_as_sc_hs__or2_2 _28024_ (.A(net312),
    .B(\tholin_riscv.regs[14][7] ),
    .Y(_21514_));
 sky130_as_sc_hs__nand3_2 _28025_ (.A(net271),
    .B(_21513_),
    .C(_21514_),
    .Y(_21515_));
 sky130_as_sc_hs__nand3_2 _28026_ (.A(net257),
    .B(_21512_),
    .C(_21515_),
    .Y(_21516_));
 sky130_as_sc_hs__or2_2 _28027_ (.A(net188),
    .B(\tholin_riscv.regs[1][7] ),
    .Y(_21517_));
 sky130_as_sc_hs__or2_2 _28028_ (.A(net312),
    .B(\tholin_riscv.regs[0][7] ),
    .Y(_21518_));
 sky130_as_sc_hs__nand3_2 _28029_ (.A(net175),
    .B(_21517_),
    .C(_21518_),
    .Y(_21519_));
 sky130_as_sc_hs__or2_2 _28030_ (.A(net188),
    .B(\tholin_riscv.regs[3][7] ),
    .Y(_21520_));
 sky130_as_sc_hs__or2_2 _28031_ (.A(net312),
    .B(\tholin_riscv.regs[2][7] ),
    .Y(_21521_));
 sky130_as_sc_hs__nand3_2 _28032_ (.A(net271),
    .B(_21520_),
    .C(_21521_),
    .Y(_21522_));
 sky130_as_sc_hs__nand3_2 _28033_ (.A(net159),
    .B(_21519_),
    .C(_21522_),
    .Y(_21523_));
 sky130_as_sc_hs__or2_2 _28034_ (.A(net189),
    .B(\tholin_riscv.regs[7][7] ),
    .Y(_21524_));
 sky130_as_sc_hs__or2_2 _28035_ (.A(net313),
    .B(\tholin_riscv.regs[6][7] ),
    .Y(_21525_));
 sky130_as_sc_hs__nand3_2 _28036_ (.A(net271),
    .B(_21524_),
    .C(_21525_),
    .Y(_21526_));
 sky130_as_sc_hs__or2_2 _28037_ (.A(net189),
    .B(\tholin_riscv.regs[5][7] ),
    .Y(_21527_));
 sky130_as_sc_hs__or2_2 _28038_ (.A(net312),
    .B(\tholin_riscv.regs[4][7] ),
    .Y(_21528_));
 sky130_as_sc_hs__nand3_2 _28039_ (.A(net175),
    .B(_21527_),
    .C(_21528_),
    .Y(_21529_));
 sky130_as_sc_hs__nand3_2 _28040_ (.A(net257),
    .B(_21526_),
    .C(_21529_),
    .Y(_21530_));
 sky130_as_sc_hs__nand3_2 _28041_ (.A(net152),
    .B(_21523_),
    .C(_21530_),
    .Y(_21531_));
 sky130_as_sc_hs__nand3_2 _28042_ (.A(net249),
    .B(_21509_),
    .C(_21516_),
    .Y(_21532_));
 sky130_as_sc_hs__nand3_2 _28043_ (.A(net150),
    .B(_21531_),
    .C(_21532_),
    .Y(_21533_));
 sky130_as_sc_hs__inv_2 _28045_ (.Y(_21535_),
    .A(_21534_));
 sky130_as_sc_hs__nand3_2 _28049_ (.A(_19754_),
    .B(_21537_),
    .C(_21538_),
    .Y(_21539_));
 sky130_as_sc_hs__nand3_2 _28050_ (.A(_19759_),
    .B(_21536_),
    .C(_21539_),
    .Y(_21540_));
 sky130_as_sc_hs__nand3_2 _28051_ (.A(_20718_),
    .B(_21471_),
    .C(_21540_),
    .Y(_21541_));
 sky130_as_sc_hs__or2_2 _28052_ (.A(\tholin_riscv.Bimm[11] ),
    .B(_20718_),
    .Y(_21542_));
 sky130_as_sc_hs__and2_2 _28053_ (.A(net500),
    .B(_21541_),
    .Y(_21543_));
 sky130_as_sc_hs__and2_2 _28054_ (.A(_21542_),
    .B(_21543_),
    .Y(_00020_));
 sky130_as_sc_hs__and2_2 _28055_ (.A(net494),
    .B(_19748_),
    .Y(_21544_));
 sky130_as_sc_hs__and2_2 _28056_ (.A(_19752_),
    .B(_21544_),
    .Y(_21545_));
 sky130_as_sc_hs__or2_2 _28058_ (.A(\tholin_riscv.load_dest[4] ),
    .B(_21546_),
    .Y(_21547_));
 sky130_as_sc_hs__or2_2 _28059_ (.A(\tholin_riscv.Bimm[4] ),
    .B(_21545_),
    .Y(_21548_));
 sky130_as_sc_hs__and2_2 _28060_ (.A(_21547_),
    .B(_21548_),
    .Y(_21549_));
 sky130_as_sc_hs__or2_2 _28062_ (.A(\tholin_riscv.load_dest[3] ),
    .B(_21546_),
    .Y(_21551_));
 sky130_as_sc_hs__or2_2 _28063_ (.A(\tholin_riscv.Bimm[3] ),
    .B(_21545_),
    .Y(_21552_));
 sky130_as_sc_hs__and2_2 _28064_ (.A(_21551_),
    .B(_21552_),
    .Y(_21553_));
 sky130_as_sc_hs__and2_2 _28066_ (.A(_21549_),
    .B(_21553_),
    .Y(_21555_));
 sky130_as_sc_hs__or2_2 _28067_ (.A(\tholin_riscv.load_dest[2] ),
    .B(_21546_),
    .Y(_21556_));
 sky130_as_sc_hs__or2_2 _28068_ (.A(\tholin_riscv.Bimm[2] ),
    .B(_21545_),
    .Y(_21557_));
 sky130_as_sc_hs__and2_2 _28069_ (.A(_21556_),
    .B(_21557_),
    .Y(_21558_));
 sky130_as_sc_hs__and2_2 _28071_ (.A(_21555_),
    .B(_21558_),
    .Y(_21560_));
 sky130_as_sc_hs__and2_2 _28072_ (.A(\tholin_riscv.cycle[3] ),
    .B(_19497_),
    .Y(_21561_));
 sky130_as_sc_hs__or2_2 _28073_ (.A(\tholin_riscv.cycle[1] ),
    .B(\tholin_riscv.mul_delay ),
    .Y(_21562_));
 sky130_as_sc_hs__and2_2 _28074_ (.A(_19498_),
    .B(_21562_),
    .Y(_21563_));
 sky130_as_sc_hs__nand3_2 _28077_ (.A(net145),
    .B(_19978_),
    .C(_19988_),
    .Y(_21566_));
 sky130_as_sc_hs__and2_2 _28079_ (.A(net497),
    .B(_21567_),
    .Y(_21568_));
 sky130_as_sc_hs__and2_2 _28081_ (.A(net502),
    .B(net145),
    .Y(_21570_));
 sky130_as_sc_hs__nor2_2 _28082_ (.A(_19475_),
    .B(_19977_),
    .Y(_21571_));
 sky130_as_sc_hs__and2_2 _28083_ (.A(_21570_),
    .B(_21571_),
    .Y(_21572_));
 sky130_as_sc_hs__nand2b_2 _28085_ (.B(_21570_),
    .Y(_21574_),
    .A(_19948_));
 sky130_as_sc_hs__nand3_2 _28086_ (.A(_21546_),
    .B(_21573_),
    .C(_21574_),
    .Y(_21575_));
 sky130_as_sc_hs__or2_2 _28087_ (.A(net413),
    .B(_21575_),
    .Y(_21576_));
 sky130_as_sc_hs__or2_2 _28088_ (.A(\tholin_riscv.load_dest[1] ),
    .B(_21546_),
    .Y(_21577_));
 sky130_as_sc_hs__or2_2 _28089_ (.A(\tholin_riscv.Bimm[1] ),
    .B(_21545_),
    .Y(_21578_));
 sky130_as_sc_hs__nor2b_2 _28091_ (.A(_21579_),
    .Y(_21580_),
    .B(_21576_));
 sky130_as_sc_hs__or2_2 _28092_ (.A(\tholin_riscv.load_dest[0] ),
    .B(_21546_),
    .Y(_21581_));
 sky130_as_sc_hs__or2_2 _28093_ (.A(\tholin_riscv.Bimm[11] ),
    .B(_21545_),
    .Y(_21582_));
 sky130_as_sc_hs__and2_2 _28094_ (.A(_21581_),
    .B(_21582_),
    .Y(_21583_));
 sky130_as_sc_hs__and2_2 _28096_ (.A(_21580_),
    .B(_21583_),
    .Y(_21585_));
 sky130_as_sc_hs__and2_2 _28097_ (.A(_21560_),
    .B(_21585_),
    .Y(_21586_));
 sky130_as_sc_hs__or2_2 _28099_ (.A(\tholin_riscv.instr[0] ),
    .B(_21546_),
    .Y(_21588_));
 sky130_as_sc_hs__and2_2 _28100_ (.A(\tholin_riscv.instr[5] ),
    .B(_21572_),
    .Y(_21589_));
 sky130_as_sc_hs__nand3_2 _28106_ (.A(net226),
    .B(_21593_),
    .C(_21594_),
    .Y(_21595_));
 sky130_as_sc_hs__nand3_2 _28109_ (.A(net365),
    .B(_21596_),
    .C(_21597_),
    .Y(_21598_));
 sky130_as_sc_hs__nand3_2 _28110_ (.A(net237),
    .B(_21595_),
    .C(_21598_),
    .Y(_21599_));
 sky130_as_sc_hs__nand3_2 _28113_ (.A(net226),
    .B(_21600_),
    .C(_21601_),
    .Y(_21602_));
 sky130_as_sc_hs__nand3_2 _28116_ (.A(net365),
    .B(_21603_),
    .C(_21604_),
    .Y(_21605_));
 sky130_as_sc_hs__nand3_2 _28117_ (.A(net348),
    .B(_21602_),
    .C(_21605_),
    .Y(_21606_));
 sky130_as_sc_hs__nand3_2 _28120_ (.A(net225),
    .B(_21607_),
    .C(_21608_),
    .Y(_21609_));
 sky130_as_sc_hs__nand3_2 _28123_ (.A(net364),
    .B(_21610_),
    .C(_21611_),
    .Y(_21612_));
 sky130_as_sc_hs__nand3_2 _28124_ (.A(net237),
    .B(_21609_),
    .C(_21612_),
    .Y(_21613_));
 sky130_as_sc_hs__nand3_2 _28127_ (.A(net364),
    .B(_21614_),
    .C(_21615_),
    .Y(_21616_));
 sky130_as_sc_hs__nand3_2 _28130_ (.A(net225),
    .B(_21617_),
    .C(_21618_),
    .Y(_21619_));
 sky130_as_sc_hs__nand3_2 _28131_ (.A(net348),
    .B(_21616_),
    .C(_21619_),
    .Y(_21620_));
 sky130_as_sc_hs__nand3_2 _28132_ (.A(net243),
    .B(_21613_),
    .C(_21620_),
    .Y(_21621_));
 sky130_as_sc_hs__nand3_2 _28133_ (.A(net339),
    .B(_21599_),
    .C(_21606_),
    .Y(_21622_));
 sky130_as_sc_hs__nand3_2 _28134_ (.A(\tholin_riscv.Jimm[19] ),
    .B(_21621_),
    .C(_21622_),
    .Y(_21623_));
 sky130_as_sc_hs__nand3_2 _28137_ (.A(net225),
    .B(_21624_),
    .C(_21625_),
    .Y(_21626_));
 sky130_as_sc_hs__nand3_2 _28140_ (.A(net365),
    .B(_21627_),
    .C(_21628_),
    .Y(_21629_));
 sky130_as_sc_hs__nand3_2 _28141_ (.A(net237),
    .B(_21626_),
    .C(_21629_),
    .Y(_21630_));
 sky130_as_sc_hs__nand3_2 _28144_ (.A(net226),
    .B(_21631_),
    .C(_21632_),
    .Y(_21633_));
 sky130_as_sc_hs__nand3_2 _28147_ (.A(net365),
    .B(_21634_),
    .C(_21635_),
    .Y(_21636_));
 sky130_as_sc_hs__nand3_2 _28148_ (.A(net348),
    .B(_21633_),
    .C(_21636_),
    .Y(_21637_));
 sky130_as_sc_hs__nand3_2 _28151_ (.A(net225),
    .B(_21638_),
    .C(_21639_),
    .Y(_21640_));
 sky130_as_sc_hs__nand3_2 _28154_ (.A(net365),
    .B(_21641_),
    .C(_21642_),
    .Y(_21643_));
 sky130_as_sc_hs__nand3_2 _28155_ (.A(net237),
    .B(_21640_),
    .C(_21643_),
    .Y(_21644_));
 sky130_as_sc_hs__nand3_2 _28158_ (.A(net364),
    .B(_21645_),
    .C(_21646_),
    .Y(_21647_));
 sky130_as_sc_hs__nand3_2 _28161_ (.A(net225),
    .B(_21648_),
    .C(_21649_),
    .Y(_21650_));
 sky130_as_sc_hs__nand3_2 _28162_ (.A(net348),
    .B(_21647_),
    .C(_21650_),
    .Y(_21651_));
 sky130_as_sc_hs__nand3_2 _28163_ (.A(net243),
    .B(_21644_),
    .C(_21651_),
    .Y(_21652_));
 sky130_as_sc_hs__nand3_2 _28164_ (.A(net339),
    .B(_21630_),
    .C(_21637_),
    .Y(_21653_));
 sky130_as_sc_hs__nand3_2 _28165_ (.A(net245),
    .B(_21652_),
    .C(_21653_),
    .Y(_21654_));
 sky130_as_sc_hs__and2_2 _28167_ (.A(\tholin_riscv.Jimm[13] ),
    .B(\tholin_riscv.Jimm[12] ),
    .Y(_21656_));
 sky130_as_sc_hs__nor2_2 _28169_ (.A(net411),
    .B(_21656_),
    .Y(_21658_));
 sky130_as_sc_hs__and2_2 _28170_ (.A(_21655_),
    .B(_21658_),
    .Y(_21659_));
 sky130_as_sc_hs__nand3_2 _28174_ (.A(net222),
    .B(_21661_),
    .C(_21662_),
    .Y(_21663_));
 sky130_as_sc_hs__nand3_2 _28177_ (.A(net362),
    .B(_21664_),
    .C(_21665_),
    .Y(_21666_));
 sky130_as_sc_hs__nand3_2 _28178_ (.A(net235),
    .B(_21663_),
    .C(_21666_),
    .Y(_21667_));
 sky130_as_sc_hs__nand3_2 _28181_ (.A(net224),
    .B(_21668_),
    .C(_21669_),
    .Y(_21670_));
 sky130_as_sc_hs__nand3_2 _28184_ (.A(net362),
    .B(_21671_),
    .C(_21672_),
    .Y(_21673_));
 sky130_as_sc_hs__nand3_2 _28185_ (.A(net346),
    .B(_21670_),
    .C(_21673_),
    .Y(_21674_));
 sky130_as_sc_hs__nand3_2 _28188_ (.A(net222),
    .B(_21675_),
    .C(_21676_),
    .Y(_21677_));
 sky130_as_sc_hs__nand3_2 _28191_ (.A(net362),
    .B(_21678_),
    .C(_21679_),
    .Y(_21680_));
 sky130_as_sc_hs__nand3_2 _28192_ (.A(net235),
    .B(_21677_),
    .C(_21680_),
    .Y(_21681_));
 sky130_as_sc_hs__nand3_2 _28195_ (.A(net362),
    .B(_21682_),
    .C(_21683_),
    .Y(_21684_));
 sky130_as_sc_hs__nand3_2 _28198_ (.A(net222),
    .B(_21685_),
    .C(_21686_),
    .Y(_21687_));
 sky130_as_sc_hs__nand3_2 _28199_ (.A(net346),
    .B(_21684_),
    .C(_21687_),
    .Y(_21688_));
 sky130_as_sc_hs__nand3_2 _28200_ (.A(net242),
    .B(_21681_),
    .C(_21688_),
    .Y(_21689_));
 sky130_as_sc_hs__nand3_2 _28201_ (.A(net340),
    .B(_21667_),
    .C(_21674_),
    .Y(_21690_));
 sky130_as_sc_hs__nand3_2 _28202_ (.A(net335),
    .B(_21689_),
    .C(_21690_),
    .Y(_21691_));
 sky130_as_sc_hs__nand3_2 _28205_ (.A(net225),
    .B(_21692_),
    .C(_21693_),
    .Y(_21694_));
 sky130_as_sc_hs__nand3_2 _28208_ (.A(net365),
    .B(_21695_),
    .C(_21696_),
    .Y(_21697_));
 sky130_as_sc_hs__nand3_2 _28209_ (.A(net237),
    .B(_21694_),
    .C(_21697_),
    .Y(_21698_));
 sky130_as_sc_hs__nand3_2 _28212_ (.A(net225),
    .B(_21699_),
    .C(_21700_),
    .Y(_21701_));
 sky130_as_sc_hs__nand3_2 _28215_ (.A(net365),
    .B(_21702_),
    .C(_21703_),
    .Y(_21704_));
 sky130_as_sc_hs__nand3_2 _28216_ (.A(net348),
    .B(_21701_),
    .C(_21704_),
    .Y(_21705_));
 sky130_as_sc_hs__nand3_2 _28219_ (.A(net225),
    .B(_21706_),
    .C(_21707_),
    .Y(_21708_));
 sky130_as_sc_hs__nand3_2 _28222_ (.A(net365),
    .B(_21709_),
    .C(_21710_),
    .Y(_21711_));
 sky130_as_sc_hs__nand3_2 _28223_ (.A(net237),
    .B(_21708_),
    .C(_21711_),
    .Y(_21712_));
 sky130_as_sc_hs__nand3_2 _28226_ (.A(net364),
    .B(_21713_),
    .C(_21714_),
    .Y(_21715_));
 sky130_as_sc_hs__nand3_2 _28229_ (.A(net226),
    .B(_21716_),
    .C(_21717_),
    .Y(_21718_));
 sky130_as_sc_hs__nand3_2 _28230_ (.A(net348),
    .B(_21715_),
    .C(_21718_),
    .Y(_21719_));
 sky130_as_sc_hs__nand3_2 _28231_ (.A(net243),
    .B(_21712_),
    .C(_21719_),
    .Y(_21720_));
 sky130_as_sc_hs__nand3_2 _28232_ (.A(net339),
    .B(_21698_),
    .C(_21705_),
    .Y(_21721_));
 sky130_as_sc_hs__nand3_2 _28233_ (.A(net245),
    .B(_21720_),
    .C(_21721_),
    .Y(_21722_));
 sky130_as_sc_hs__or2_2 _28235_ (.A(net400),
    .B(\tholin_riscv.regs[24][19] ),
    .Y(_21724_));
 sky130_as_sc_hs__nand3_2 _28237_ (.A(net224),
    .B(_21724_),
    .C(_21725_),
    .Y(_21726_));
 sky130_as_sc_hs__or2_2 _28238_ (.A(net400),
    .B(\tholin_riscv.regs[26][19] ),
    .Y(_21727_));
 sky130_as_sc_hs__nand3_2 _28240_ (.A(net368),
    .B(_21727_),
    .C(_21728_),
    .Y(_21729_));
 sky130_as_sc_hs__nand3_2 _28241_ (.A(net235),
    .B(_21726_),
    .C(_21729_),
    .Y(_21730_));
 sky130_as_sc_hs__or2_2 _28242_ (.A(net400),
    .B(\tholin_riscv.regs[28][19] ),
    .Y(_21731_));
 sky130_as_sc_hs__nand3_2 _28244_ (.A(net224),
    .B(_21731_),
    .C(_21732_),
    .Y(_21733_));
 sky130_as_sc_hs__or2_2 _28245_ (.A(net400),
    .B(\tholin_riscv.regs[30][19] ),
    .Y(_21734_));
 sky130_as_sc_hs__nand3_2 _28247_ (.A(net368),
    .B(_21734_),
    .C(_21735_),
    .Y(_21736_));
 sky130_as_sc_hs__nand3_2 _28248_ (.A(net349),
    .B(_21733_),
    .C(_21736_),
    .Y(_21737_));
 sky130_as_sc_hs__or2_2 _28249_ (.A(net399),
    .B(\tholin_riscv.regs[16][19] ),
    .Y(_21738_));
 sky130_as_sc_hs__nand3_2 _28251_ (.A(net229),
    .B(_21738_),
    .C(_21739_),
    .Y(_21740_));
 sky130_as_sc_hs__or2_2 _28252_ (.A(net399),
    .B(\tholin_riscv.regs[18][19] ),
    .Y(_21741_));
 sky130_as_sc_hs__nand3_2 _28254_ (.A(net368),
    .B(_21741_),
    .C(_21742_),
    .Y(_21743_));
 sky130_as_sc_hs__nand3_2 _28255_ (.A(net239),
    .B(_21740_),
    .C(_21743_),
    .Y(_21744_));
 sky130_as_sc_hs__or2_2 _28256_ (.A(net398),
    .B(\tholin_riscv.regs[22][19] ),
    .Y(_21745_));
 sky130_as_sc_hs__nand3_2 _28258_ (.A(net368),
    .B(_21745_),
    .C(_21746_),
    .Y(_21747_));
 sky130_as_sc_hs__or2_2 _28259_ (.A(net398),
    .B(\tholin_riscv.regs[20][19] ),
    .Y(_21748_));
 sky130_as_sc_hs__nand3_2 _28261_ (.A(net229),
    .B(_21748_),
    .C(_21749_),
    .Y(_21750_));
 sky130_as_sc_hs__nand3_2 _28262_ (.A(net349),
    .B(_21747_),
    .C(_21750_),
    .Y(_21751_));
 sky130_as_sc_hs__nand3_2 _28263_ (.A(net243),
    .B(_21744_),
    .C(_21751_),
    .Y(_21752_));
 sky130_as_sc_hs__nand3_2 _28264_ (.A(net339),
    .B(_21730_),
    .C(_21737_),
    .Y(_21753_));
 sky130_as_sc_hs__nand3_2 _28265_ (.A(net335),
    .B(_21752_),
    .C(_21753_),
    .Y(_21754_));
 sky130_as_sc_hs__or2_2 _28266_ (.A(net401),
    .B(\tholin_riscv.regs[8][19] ),
    .Y(_21755_));
 sky130_as_sc_hs__nand3_2 _28268_ (.A(net225),
    .B(_21755_),
    .C(_21756_),
    .Y(_21757_));
 sky130_as_sc_hs__or2_2 _28269_ (.A(net409),
    .B(\tholin_riscv.regs[10][19] ),
    .Y(_21758_));
 sky130_as_sc_hs__nand3_2 _28271_ (.A(net365),
    .B(_21758_),
    .C(_21759_),
    .Y(_21760_));
 sky130_as_sc_hs__nand3_2 _28272_ (.A(net237),
    .B(_21757_),
    .C(_21760_),
    .Y(_21761_));
 sky130_as_sc_hs__or2_2 _28273_ (.A(net409),
    .B(\tholin_riscv.regs[12][19] ),
    .Y(_21762_));
 sky130_as_sc_hs__nand3_2 _28275_ (.A(net225),
    .B(_21762_),
    .C(_21763_),
    .Y(_21764_));
 sky130_as_sc_hs__or2_2 _28276_ (.A(net409),
    .B(\tholin_riscv.regs[14][19] ),
    .Y(_21765_));
 sky130_as_sc_hs__nand3_2 _28278_ (.A(net365),
    .B(_21765_),
    .C(_21766_),
    .Y(_21767_));
 sky130_as_sc_hs__nand3_2 _28279_ (.A(net348),
    .B(_21764_),
    .C(_21767_),
    .Y(_21768_));
 sky130_as_sc_hs__or2_2 _28280_ (.A(net401),
    .B(\tholin_riscv.regs[0][19] ),
    .Y(_21769_));
 sky130_as_sc_hs__nand3_2 _28282_ (.A(net225),
    .B(_21769_),
    .C(_21770_),
    .Y(_21771_));
 sky130_as_sc_hs__or2_2 _28283_ (.A(net401),
    .B(\tholin_riscv.regs[2][19] ),
    .Y(_21772_));
 sky130_as_sc_hs__nand3_2 _28285_ (.A(net365),
    .B(_21772_),
    .C(_21773_),
    .Y(_21774_));
 sky130_as_sc_hs__nand3_2 _28286_ (.A(net237),
    .B(_21771_),
    .C(_21774_),
    .Y(_21775_));
 sky130_as_sc_hs__or2_2 _28287_ (.A(net401),
    .B(\tholin_riscv.regs[6][19] ),
    .Y(_21776_));
 sky130_as_sc_hs__nand3_2 _28289_ (.A(net366),
    .B(_21776_),
    .C(_21777_),
    .Y(_21778_));
 sky130_as_sc_hs__or2_2 _28290_ (.A(net401),
    .B(\tholin_riscv.regs[4][19] ),
    .Y(_21779_));
 sky130_as_sc_hs__nand3_2 _28292_ (.A(net225),
    .B(_21779_),
    .C(_21780_),
    .Y(_21781_));
 sky130_as_sc_hs__nand3_2 _28293_ (.A(net350),
    .B(_21778_),
    .C(_21781_),
    .Y(_21782_));
 sky130_as_sc_hs__nand3_2 _28294_ (.A(net243),
    .B(_21775_),
    .C(_21782_),
    .Y(_21783_));
 sky130_as_sc_hs__nand3_2 _28295_ (.A(net339),
    .B(_21761_),
    .C(_21768_),
    .Y(_21784_));
 sky130_as_sc_hs__nand3_2 _28296_ (.A(net245),
    .B(_21783_),
    .C(_21784_),
    .Y(_21785_));
 sky130_as_sc_hs__inv_2 _28298_ (.Y(_21787_),
    .A(_21786_));
 sky130_as_sc_hs__or2_2 _28299_ (.A(net406),
    .B(\tholin_riscv.regs[24][17] ),
    .Y(_21788_));
 sky130_as_sc_hs__nand3_2 _28301_ (.A(net230),
    .B(_21788_),
    .C(_21789_),
    .Y(_21790_));
 sky130_as_sc_hs__or2_2 _28302_ (.A(net406),
    .B(\tholin_riscv.regs[26][17] ),
    .Y(_21791_));
 sky130_as_sc_hs__nand3_2 _28304_ (.A(net369),
    .B(_21791_),
    .C(_21792_),
    .Y(_21793_));
 sky130_as_sc_hs__nand3_2 _28305_ (.A(net238),
    .B(_21790_),
    .C(_21793_),
    .Y(_21794_));
 sky130_as_sc_hs__or2_2 _28306_ (.A(net406),
    .B(\tholin_riscv.regs[28][17] ),
    .Y(_21795_));
 sky130_as_sc_hs__nand3_2 _28308_ (.A(net230),
    .B(_21795_),
    .C(_21796_),
    .Y(_21797_));
 sky130_as_sc_hs__or2_2 _28309_ (.A(net406),
    .B(\tholin_riscv.regs[30][17] ),
    .Y(_21798_));
 sky130_as_sc_hs__nand3_2 _28311_ (.A(net369),
    .B(_21798_),
    .C(_21799_),
    .Y(_21800_));
 sky130_as_sc_hs__nand3_2 _28312_ (.A(net349),
    .B(_21797_),
    .C(_21800_),
    .Y(_21801_));
 sky130_as_sc_hs__or2_2 _28313_ (.A(net405),
    .B(\tholin_riscv.regs[16][17] ),
    .Y(_21802_));
 sky130_as_sc_hs__nand3_2 _28315_ (.A(net228),
    .B(_21802_),
    .C(_21803_),
    .Y(_21804_));
 sky130_as_sc_hs__or2_2 _28316_ (.A(net405),
    .B(\tholin_riscv.regs[18][17] ),
    .Y(_21805_));
 sky130_as_sc_hs__nand3_2 _28318_ (.A(net367),
    .B(_21805_),
    .C(_21806_),
    .Y(_21807_));
 sky130_as_sc_hs__nand3_2 _28319_ (.A(net238),
    .B(_21804_),
    .C(_21807_),
    .Y(_21808_));
 sky130_as_sc_hs__or2_2 _28320_ (.A(net405),
    .B(\tholin_riscv.regs[22][17] ),
    .Y(_21809_));
 sky130_as_sc_hs__nand3_2 _28322_ (.A(net367),
    .B(_21809_),
    .C(_21810_),
    .Y(_21811_));
 sky130_as_sc_hs__or2_2 _28323_ (.A(net406),
    .B(\tholin_riscv.regs[20][17] ),
    .Y(_21812_));
 sky130_as_sc_hs__nand3_2 _28325_ (.A(net228),
    .B(_21812_),
    .C(_21813_),
    .Y(_21814_));
 sky130_as_sc_hs__nand3_2 _28326_ (.A(net350),
    .B(_21811_),
    .C(_21814_),
    .Y(_21815_));
 sky130_as_sc_hs__nand3_2 _28327_ (.A(net244),
    .B(_21808_),
    .C(_21815_),
    .Y(_21816_));
 sky130_as_sc_hs__nand3_2 _28328_ (.A(net339),
    .B(_21794_),
    .C(_21801_),
    .Y(_21817_));
 sky130_as_sc_hs__nand3_2 _28329_ (.A(net335),
    .B(_21816_),
    .C(_21817_),
    .Y(_21818_));
 sky130_as_sc_hs__or2_2 _28330_ (.A(net403),
    .B(\tholin_riscv.regs[8][17] ),
    .Y(_21819_));
 sky130_as_sc_hs__nand3_2 _28332_ (.A(net227),
    .B(_21819_),
    .C(_21820_),
    .Y(_21821_));
 sky130_as_sc_hs__or2_2 _28333_ (.A(net404),
    .B(\tholin_riscv.regs[10][17] ),
    .Y(_21822_));
 sky130_as_sc_hs__nand3_2 _28335_ (.A(net366),
    .B(_21822_),
    .C(_21823_),
    .Y(_21824_));
 sky130_as_sc_hs__nand3_2 _28336_ (.A(net238),
    .B(_21821_),
    .C(_21824_),
    .Y(_21825_));
 sky130_as_sc_hs__or2_2 _28337_ (.A(net403),
    .B(\tholin_riscv.regs[12][17] ),
    .Y(_21826_));
 sky130_as_sc_hs__nand3_2 _28339_ (.A(net227),
    .B(_21826_),
    .C(_21827_),
    .Y(_21828_));
 sky130_as_sc_hs__or2_2 _28340_ (.A(net403),
    .B(\tholin_riscv.regs[14][17] ),
    .Y(_21829_));
 sky130_as_sc_hs__nand3_2 _28342_ (.A(net366),
    .B(_21829_),
    .C(_21830_),
    .Y(_21831_));
 sky130_as_sc_hs__nand3_2 _28343_ (.A(net350),
    .B(_21828_),
    .C(_21831_),
    .Y(_21832_));
 sky130_as_sc_hs__or2_2 _28344_ (.A(net404),
    .B(\tholin_riscv.regs[0][17] ),
    .Y(_21833_));
 sky130_as_sc_hs__nand3_2 _28346_ (.A(net227),
    .B(_21833_),
    .C(_21834_),
    .Y(_21835_));
 sky130_as_sc_hs__or2_2 _28347_ (.A(net403),
    .B(\tholin_riscv.regs[2][17] ),
    .Y(_21836_));
 sky130_as_sc_hs__nand3_2 _28349_ (.A(net366),
    .B(_21836_),
    .C(_21837_),
    .Y(_21838_));
 sky130_as_sc_hs__nand3_2 _28350_ (.A(net238),
    .B(_21835_),
    .C(_21838_),
    .Y(_21839_));
 sky130_as_sc_hs__or2_2 _28351_ (.A(net403),
    .B(\tholin_riscv.regs[6][17] ),
    .Y(_21840_));
 sky130_as_sc_hs__nand3_2 _28353_ (.A(net366),
    .B(_21840_),
    .C(_21841_),
    .Y(_21842_));
 sky130_as_sc_hs__or2_2 _28354_ (.A(net403),
    .B(\tholin_riscv.regs[4][17] ),
    .Y(_21843_));
 sky130_as_sc_hs__nand3_2 _28356_ (.A(net227),
    .B(_21843_),
    .C(_21844_),
    .Y(_21845_));
 sky130_as_sc_hs__nand3_2 _28357_ (.A(net350),
    .B(_21842_),
    .C(_21845_),
    .Y(_21846_));
 sky130_as_sc_hs__nand3_2 _28358_ (.A(net243),
    .B(_21839_),
    .C(_21846_),
    .Y(_21847_));
 sky130_as_sc_hs__nand3_2 _28359_ (.A(net339),
    .B(_21825_),
    .C(_21832_),
    .Y(_21848_));
 sky130_as_sc_hs__nand3_2 _28360_ (.A(net245),
    .B(_21847_),
    .C(_21848_),
    .Y(_21849_));
 sky130_as_sc_hs__inv_2 _28362_ (.Y(_21851_),
    .A(_21850_));
 sky130_as_sc_hs__or2_2 _28363_ (.A(net385),
    .B(\tholin_riscv.regs[24][5] ),
    .Y(_21852_));
 sky130_as_sc_hs__or2_2 _28364_ (.A(net205),
    .B(\tholin_riscv.regs[25][5] ),
    .Y(_21853_));
 sky130_as_sc_hs__nand3_2 _28365_ (.A(net217),
    .B(_21852_),
    .C(_21853_),
    .Y(_21854_));
 sky130_as_sc_hs__or2_2 _28366_ (.A(net385),
    .B(\tholin_riscv.regs[26][5] ),
    .Y(_21855_));
 sky130_as_sc_hs__or2_2 _28367_ (.A(net205),
    .B(\tholin_riscv.regs[27][5] ),
    .Y(_21856_));
 sky130_as_sc_hs__nand3_2 _28368_ (.A(net358),
    .B(_21855_),
    .C(_21856_),
    .Y(_21857_));
 sky130_as_sc_hs__nand3_2 _28369_ (.A(net233),
    .B(_21854_),
    .C(_21857_),
    .Y(_21858_));
 sky130_as_sc_hs__or2_2 _28370_ (.A(net385),
    .B(\tholin_riscv.regs[28][5] ),
    .Y(_21859_));
 sky130_as_sc_hs__or2_2 _28371_ (.A(net205),
    .B(\tholin_riscv.regs[29][5] ),
    .Y(_21860_));
 sky130_as_sc_hs__nand3_2 _28372_ (.A(net214),
    .B(_21859_),
    .C(_21860_),
    .Y(_21861_));
 sky130_as_sc_hs__or2_2 _28373_ (.A(net386),
    .B(\tholin_riscv.regs[30][5] ),
    .Y(_21862_));
 sky130_as_sc_hs__or2_2 _28374_ (.A(net205),
    .B(\tholin_riscv.regs[31][5] ),
    .Y(_21863_));
 sky130_as_sc_hs__nand3_2 _28375_ (.A(net358),
    .B(_21862_),
    .C(_21863_),
    .Y(_21864_));
 sky130_as_sc_hs__nand3_2 _28376_ (.A(net345),
    .B(_21861_),
    .C(_21864_),
    .Y(_21865_));
 sky130_as_sc_hs__or2_2 _28377_ (.A(net385),
    .B(\tholin_riscv.regs[16][5] ),
    .Y(_21866_));
 sky130_as_sc_hs__or2_2 _28378_ (.A(net205),
    .B(\tholin_riscv.regs[17][5] ),
    .Y(_21867_));
 sky130_as_sc_hs__nand3_2 _28379_ (.A(net217),
    .B(_21866_),
    .C(_21867_),
    .Y(_21868_));
 sky130_as_sc_hs__or2_2 _28380_ (.A(net385),
    .B(\tholin_riscv.regs[18][5] ),
    .Y(_21869_));
 sky130_as_sc_hs__or2_2 _28381_ (.A(net205),
    .B(\tholin_riscv.regs[19][5] ),
    .Y(_21870_));
 sky130_as_sc_hs__nand3_2 _28382_ (.A(net358),
    .B(_21869_),
    .C(_21870_),
    .Y(_21871_));
 sky130_as_sc_hs__nand3_2 _28383_ (.A(net233),
    .B(_21868_),
    .C(_21871_),
    .Y(_21872_));
 sky130_as_sc_hs__or2_2 _28384_ (.A(net386),
    .B(\tholin_riscv.regs[22][5] ),
    .Y(_21873_));
 sky130_as_sc_hs__or2_2 _28385_ (.A(net205),
    .B(\tholin_riscv.regs[23][5] ),
    .Y(_21874_));
 sky130_as_sc_hs__nand3_2 _28386_ (.A(net358),
    .B(_21873_),
    .C(_21874_),
    .Y(_21875_));
 sky130_as_sc_hs__or2_2 _28387_ (.A(net386),
    .B(\tholin_riscv.regs[20][5] ),
    .Y(_21876_));
 sky130_as_sc_hs__or2_2 _28388_ (.A(net205),
    .B(\tholin_riscv.regs[21][5] ),
    .Y(_21877_));
 sky130_as_sc_hs__nand3_2 _28389_ (.A(net214),
    .B(_21876_),
    .C(_21877_),
    .Y(_21878_));
 sky130_as_sc_hs__nand3_2 _28390_ (.A(net345),
    .B(_21875_),
    .C(_21878_),
    .Y(_21879_));
 sky130_as_sc_hs__nand3_2 _28391_ (.A(net241),
    .B(_21872_),
    .C(_21879_),
    .Y(_21880_));
 sky130_as_sc_hs__nand3_2 _28392_ (.A(net338),
    .B(_21858_),
    .C(_21865_),
    .Y(_21881_));
 sky130_as_sc_hs__nand3_2 _28393_ (.A(net336),
    .B(_21880_),
    .C(_21881_),
    .Y(_21882_));
 sky130_as_sc_hs__or2_2 _28394_ (.A(net409),
    .B(\tholin_riscv.regs[8][5] ),
    .Y(_21883_));
 sky130_as_sc_hs__or2_2 _28395_ (.A(net205),
    .B(\tholin_riscv.regs[9][5] ),
    .Y(_21884_));
 sky130_as_sc_hs__nand3_2 _28396_ (.A(net225),
    .B(_21883_),
    .C(_21884_),
    .Y(_21885_));
 sky130_as_sc_hs__or2_2 _28397_ (.A(net409),
    .B(\tholin_riscv.regs[10][5] ),
    .Y(_21886_));
 sky130_as_sc_hs__or2_2 _28398_ (.A(net205),
    .B(\tholin_riscv.regs[11][5] ),
    .Y(_21887_));
 sky130_as_sc_hs__nand3_2 _28399_ (.A(net365),
    .B(_21886_),
    .C(_21887_),
    .Y(_21888_));
 sky130_as_sc_hs__nand3_2 _28400_ (.A(net237),
    .B(_21885_),
    .C(_21888_),
    .Y(_21889_));
 sky130_as_sc_hs__or2_2 _28401_ (.A(net385),
    .B(\tholin_riscv.regs[12][5] ),
    .Y(_21890_));
 sky130_as_sc_hs__or2_2 _28402_ (.A(net209),
    .B(\tholin_riscv.regs[13][5] ),
    .Y(_21891_));
 sky130_as_sc_hs__nand3_2 _28403_ (.A(net217),
    .B(_21890_),
    .C(_21891_),
    .Y(_21892_));
 sky130_as_sc_hs__or2_2 _28404_ (.A(net410),
    .B(\tholin_riscv.regs[14][5] ),
    .Y(_21893_));
 sky130_as_sc_hs__or2_2 _28405_ (.A(net205),
    .B(\tholin_riscv.regs[15][5] ),
    .Y(_21894_));
 sky130_as_sc_hs__nand3_2 _28406_ (.A(net358),
    .B(_21893_),
    .C(_21894_),
    .Y(_21895_));
 sky130_as_sc_hs__nand3_2 _28407_ (.A(net345),
    .B(_21892_),
    .C(_21895_),
    .Y(_21896_));
 sky130_as_sc_hs__or2_2 _28408_ (.A(net410),
    .B(\tholin_riscv.regs[0][5] ),
    .Y(_21897_));
 sky130_as_sc_hs__or2_2 _28409_ (.A(net205),
    .B(\tholin_riscv.regs[1][5] ),
    .Y(_21898_));
 sky130_as_sc_hs__nand3_2 _28410_ (.A(net217),
    .B(_21897_),
    .C(_21898_),
    .Y(_21899_));
 sky130_as_sc_hs__or2_2 _28411_ (.A(net385),
    .B(\tholin_riscv.regs[2][5] ),
    .Y(_21900_));
 sky130_as_sc_hs__or2_2 _28412_ (.A(net205),
    .B(\tholin_riscv.regs[3][5] ),
    .Y(_21901_));
 sky130_as_sc_hs__nand3_2 _28413_ (.A(net358),
    .B(_21900_),
    .C(_21901_),
    .Y(_21902_));
 sky130_as_sc_hs__nand3_2 _28414_ (.A(net234),
    .B(_21899_),
    .C(_21902_),
    .Y(_21903_));
 sky130_as_sc_hs__or2_2 _28415_ (.A(net385),
    .B(\tholin_riscv.regs[6][5] ),
    .Y(_21904_));
 sky130_as_sc_hs__or2_2 _28416_ (.A(net205),
    .B(\tholin_riscv.regs[7][5] ),
    .Y(_21905_));
 sky130_as_sc_hs__nand3_2 _28417_ (.A(net358),
    .B(_21904_),
    .C(_21905_),
    .Y(_21906_));
 sky130_as_sc_hs__or2_2 _28418_ (.A(net385),
    .B(\tholin_riscv.regs[4][5] ),
    .Y(_21907_));
 sky130_as_sc_hs__or2_2 _28419_ (.A(net205),
    .B(\tholin_riscv.regs[5][5] ),
    .Y(_21908_));
 sky130_as_sc_hs__nand3_2 _28420_ (.A(net217),
    .B(_21907_),
    .C(_21908_),
    .Y(_21909_));
 sky130_as_sc_hs__nand3_2 _28421_ (.A(net345),
    .B(_21906_),
    .C(_21909_),
    .Y(_21910_));
 sky130_as_sc_hs__nand3_2 _28422_ (.A(net241),
    .B(_21903_),
    .C(_21910_),
    .Y(_21911_));
 sky130_as_sc_hs__nand3_2 _28423_ (.A(net338),
    .B(_21889_),
    .C(_21896_),
    .Y(_21912_));
 sky130_as_sc_hs__nand3_2 _28424_ (.A(net245),
    .B(_21911_),
    .C(_21912_),
    .Y(_21913_));
 sky130_as_sc_hs__and2_2 _28425_ (.A(_21882_),
    .B(_21913_),
    .Y(_21914_));
 sky130_as_sc_hs__or2_2 _28426_ (.A(net372),
    .B(\tholin_riscv.regs[24][3] ),
    .Y(_21915_));
 sky130_as_sc_hs__or2_2 _28427_ (.A(net204),
    .B(\tholin_riscv.regs[25][3] ),
    .Y(_21916_));
 sky130_as_sc_hs__nand3_2 _28428_ (.A(net214),
    .B(_21915_),
    .C(_21916_),
    .Y(_21917_));
 sky130_as_sc_hs__or2_2 _28429_ (.A(net372),
    .B(\tholin_riscv.regs[26][3] ),
    .Y(_21918_));
 sky130_as_sc_hs__or2_2 _28430_ (.A(net204),
    .B(\tholin_riscv.regs[27][3] ),
    .Y(_21919_));
 sky130_as_sc_hs__nand3_2 _28431_ (.A(net354),
    .B(_21918_),
    .C(_21919_),
    .Y(_21920_));
 sky130_as_sc_hs__nand3_2 _28432_ (.A(net232),
    .B(_21917_),
    .C(_21920_),
    .Y(_21921_));
 sky130_as_sc_hs__or2_2 _28433_ (.A(net386),
    .B(\tholin_riscv.regs[28][3] ),
    .Y(_21922_));
 sky130_as_sc_hs__or2_2 _28434_ (.A(net204),
    .B(\tholin_riscv.regs[29][3] ),
    .Y(_21923_));
 sky130_as_sc_hs__nand3_2 _28435_ (.A(net214),
    .B(_21922_),
    .C(_21923_),
    .Y(_21924_));
 sky130_as_sc_hs__or2_2 _28436_ (.A(net372),
    .B(\tholin_riscv.regs[30][3] ),
    .Y(_21925_));
 sky130_as_sc_hs__or2_2 _28437_ (.A(net204),
    .B(\tholin_riscv.regs[31][3] ),
    .Y(_21926_));
 sky130_as_sc_hs__nand3_2 _28438_ (.A(net354),
    .B(_21925_),
    .C(_21926_),
    .Y(_21927_));
 sky130_as_sc_hs__nand3_2 _28439_ (.A(net343),
    .B(_21924_),
    .C(_21927_),
    .Y(_21928_));
 sky130_as_sc_hs__or2_2 _28440_ (.A(net373),
    .B(\tholin_riscv.regs[16][3] ),
    .Y(_21929_));
 sky130_as_sc_hs__or2_2 _28441_ (.A(net201),
    .B(\tholin_riscv.regs[17][3] ),
    .Y(_21930_));
 sky130_as_sc_hs__nand3_2 _28442_ (.A(net214),
    .B(_21929_),
    .C(_21930_),
    .Y(_21931_));
 sky130_as_sc_hs__or2_2 _28443_ (.A(net373),
    .B(\tholin_riscv.regs[18][3] ),
    .Y(_21932_));
 sky130_as_sc_hs__or2_2 _28444_ (.A(net201),
    .B(\tholin_riscv.regs[19][3] ),
    .Y(_21933_));
 sky130_as_sc_hs__nand3_2 _28445_ (.A(net354),
    .B(_21932_),
    .C(_21933_),
    .Y(_21934_));
 sky130_as_sc_hs__nand3_2 _28446_ (.A(net232),
    .B(_21931_),
    .C(_21934_),
    .Y(_21935_));
 sky130_as_sc_hs__or2_2 _28447_ (.A(net372),
    .B(\tholin_riscv.regs[22][3] ),
    .Y(_21936_));
 sky130_as_sc_hs__or2_2 _28448_ (.A(net201),
    .B(\tholin_riscv.regs[23][3] ),
    .Y(_21937_));
 sky130_as_sc_hs__nand3_2 _28449_ (.A(net354),
    .B(_21936_),
    .C(_21937_),
    .Y(_21938_));
 sky130_as_sc_hs__or2_2 _28450_ (.A(net372),
    .B(\tholin_riscv.regs[20][3] ),
    .Y(_21939_));
 sky130_as_sc_hs__or2_2 _28451_ (.A(net204),
    .B(\tholin_riscv.regs[21][3] ),
    .Y(_21940_));
 sky130_as_sc_hs__nand3_2 _28452_ (.A(net213),
    .B(_21939_),
    .C(_21940_),
    .Y(_21941_));
 sky130_as_sc_hs__nand3_2 _28453_ (.A(net343),
    .B(_21938_),
    .C(_21941_),
    .Y(_21942_));
 sky130_as_sc_hs__nand3_2 _28454_ (.A(net240),
    .B(_21935_),
    .C(_21942_),
    .Y(_21943_));
 sky130_as_sc_hs__nand3_2 _28455_ (.A(net337),
    .B(_21921_),
    .C(_21928_),
    .Y(_21944_));
 sky130_as_sc_hs__nand3_2 _28456_ (.A(net336),
    .B(_21943_),
    .C(_21944_),
    .Y(_21945_));
 sky130_as_sc_hs__or2_2 _28457_ (.A(net386),
    .B(\tholin_riscv.regs[8][3] ),
    .Y(_21946_));
 sky130_as_sc_hs__or2_2 _28458_ (.A(net204),
    .B(\tholin_riscv.regs[9][3] ),
    .Y(_21947_));
 sky130_as_sc_hs__nand3_2 _28459_ (.A(net214),
    .B(_21946_),
    .C(_21947_),
    .Y(_21948_));
 sky130_as_sc_hs__or2_2 _28460_ (.A(net386),
    .B(\tholin_riscv.regs[10][3] ),
    .Y(_21949_));
 sky130_as_sc_hs__or2_2 _28461_ (.A(net204),
    .B(\tholin_riscv.regs[11][3] ),
    .Y(_21950_));
 sky130_as_sc_hs__nand3_2 _28462_ (.A(net354),
    .B(_21949_),
    .C(_21950_),
    .Y(_21951_));
 sky130_as_sc_hs__nand3_2 _28463_ (.A(_19483_),
    .B(_21948_),
    .C(_21951_),
    .Y(_21952_));
 sky130_as_sc_hs__or2_2 _28464_ (.A(net386),
    .B(\tholin_riscv.regs[12][3] ),
    .Y(_21953_));
 sky130_as_sc_hs__or2_2 _28465_ (.A(net204),
    .B(\tholin_riscv.regs[13][3] ),
    .Y(_21954_));
 sky130_as_sc_hs__nand3_2 _28466_ (.A(net214),
    .B(_21953_),
    .C(_21954_),
    .Y(_21955_));
 sky130_as_sc_hs__or2_2 _28467_ (.A(net386),
    .B(\tholin_riscv.regs[14][3] ),
    .Y(_21956_));
 sky130_as_sc_hs__or2_2 _28468_ (.A(net204),
    .B(\tholin_riscv.regs[15][3] ),
    .Y(_21957_));
 sky130_as_sc_hs__nand3_2 _28469_ (.A(net354),
    .B(_21956_),
    .C(_21957_),
    .Y(_21958_));
 sky130_as_sc_hs__nand3_2 _28470_ (.A(net342),
    .B(_21955_),
    .C(_21958_),
    .Y(_21959_));
 sky130_as_sc_hs__or2_2 _28471_ (.A(net386),
    .B(\tholin_riscv.regs[0][3] ),
    .Y(_21960_));
 sky130_as_sc_hs__or2_2 _28472_ (.A(net202),
    .B(\tholin_riscv.regs[1][3] ),
    .Y(_21961_));
 sky130_as_sc_hs__nand3_2 _28473_ (.A(net214),
    .B(_21960_),
    .C(_21961_),
    .Y(_21962_));
 sky130_as_sc_hs__or2_2 _28474_ (.A(net386),
    .B(\tholin_riscv.regs[2][3] ),
    .Y(_21963_));
 sky130_as_sc_hs__or2_2 _28475_ (.A(net202),
    .B(\tholin_riscv.regs[3][3] ),
    .Y(_21964_));
 sky130_as_sc_hs__nand3_2 _28476_ (.A(net354),
    .B(_21963_),
    .C(_21964_),
    .Y(_21965_));
 sky130_as_sc_hs__nand3_2 _28477_ (.A(net232),
    .B(_21962_),
    .C(_21965_),
    .Y(_21966_));
 sky130_as_sc_hs__or2_2 _28478_ (.A(net386),
    .B(\tholin_riscv.regs[6][3] ),
    .Y(_21967_));
 sky130_as_sc_hs__or2_2 _28479_ (.A(net201),
    .B(\tholin_riscv.regs[7][3] ),
    .Y(_21968_));
 sky130_as_sc_hs__nand3_2 _28480_ (.A(net354),
    .B(_21967_),
    .C(_21968_),
    .Y(_21969_));
 sky130_as_sc_hs__or2_2 _28481_ (.A(net386),
    .B(\tholin_riscv.regs[4][3] ),
    .Y(_21970_));
 sky130_as_sc_hs__or2_2 _28482_ (.A(net203),
    .B(\tholin_riscv.regs[5][3] ),
    .Y(_21971_));
 sky130_as_sc_hs__nand3_2 _28483_ (.A(net214),
    .B(_21970_),
    .C(_21971_),
    .Y(_21972_));
 sky130_as_sc_hs__nand3_2 _28484_ (.A(net343),
    .B(_21969_),
    .C(_21972_),
    .Y(_21973_));
 sky130_as_sc_hs__nand3_2 _28485_ (.A(net240),
    .B(_21966_),
    .C(_21973_),
    .Y(_21974_));
 sky130_as_sc_hs__nand3_2 _28486_ (.A(net337),
    .B(_21952_),
    .C(_21959_),
    .Y(_21975_));
 sky130_as_sc_hs__nand3_2 _28487_ (.A(net246),
    .B(_21974_),
    .C(_21975_),
    .Y(_21976_));
 sky130_as_sc_hs__and2_2 _28488_ (.A(_21945_),
    .B(_21976_),
    .Y(_21977_));
 sky130_as_sc_hs__or2_2 _28489_ (.A(net372),
    .B(\tholin_riscv.regs[24][2] ),
    .Y(_21978_));
 sky130_as_sc_hs__nand2b_2 _28490_ (.B(net372),
    .Y(_21979_),
    .A(\tholin_riscv.regs[25][2] ));
 sky130_as_sc_hs__nand3_2 _28491_ (.A(net214),
    .B(_21978_),
    .C(_21979_),
    .Y(_21980_));
 sky130_as_sc_hs__or2_2 _28492_ (.A(net373),
    .B(\tholin_riscv.regs[26][2] ),
    .Y(_21981_));
 sky130_as_sc_hs__nand2b_2 _28493_ (.B(net375),
    .Y(_21982_),
    .A(\tholin_riscv.regs[27][2] ));
 sky130_as_sc_hs__nand3_2 _28494_ (.A(net354),
    .B(_21981_),
    .C(_21982_),
    .Y(_21983_));
 sky130_as_sc_hs__nand3_2 _28495_ (.A(net231),
    .B(_21980_),
    .C(_21983_),
    .Y(_21984_));
 sky130_as_sc_hs__or2_2 _28496_ (.A(net375),
    .B(\tholin_riscv.regs[28][2] ),
    .Y(_21985_));
 sky130_as_sc_hs__nand2b_2 _28497_ (.B(net375),
    .Y(_21986_),
    .A(\tholin_riscv.regs[29][2] ));
 sky130_as_sc_hs__nand3_2 _28498_ (.A(net220),
    .B(_21985_),
    .C(_21986_),
    .Y(_21987_));
 sky130_as_sc_hs__or2_2 _28499_ (.A(net375),
    .B(\tholin_riscv.regs[30][2] ),
    .Y(_21988_));
 sky130_as_sc_hs__nand2b_2 _28500_ (.B(net375),
    .Y(_21989_),
    .A(\tholin_riscv.regs[31][2] ));
 sky130_as_sc_hs__nand3_2 _28501_ (.A(net361),
    .B(_21988_),
    .C(_21989_),
    .Y(_21990_));
 sky130_as_sc_hs__nand3_2 _28502_ (.A(net347),
    .B(_21987_),
    .C(_21990_),
    .Y(_21991_));
 sky130_as_sc_hs__or2_2 _28503_ (.A(net373),
    .B(\tholin_riscv.regs[16][2] ),
    .Y(_21992_));
 sky130_as_sc_hs__nand2b_2 _28504_ (.B(net372),
    .Y(_21993_),
    .A(\tholin_riscv.regs[17][2] ));
 sky130_as_sc_hs__nand3_2 _28505_ (.A(net213),
    .B(_21992_),
    .C(_21993_),
    .Y(_21994_));
 sky130_as_sc_hs__or2_2 _28506_ (.A(net373),
    .B(\tholin_riscv.regs[18][2] ),
    .Y(_21995_));
 sky130_as_sc_hs__nand2b_2 _28507_ (.B(net375),
    .Y(_21996_),
    .A(\tholin_riscv.regs[19][2] ));
 sky130_as_sc_hs__nand3_2 _28508_ (.A(net354),
    .B(_21995_),
    .C(_21996_),
    .Y(_21997_));
 sky130_as_sc_hs__nand3_2 _28509_ (.A(net231),
    .B(_21994_),
    .C(_21997_),
    .Y(_21998_));
 sky130_as_sc_hs__or2_2 _28510_ (.A(net374),
    .B(\tholin_riscv.regs[22][2] ),
    .Y(_21999_));
 sky130_as_sc_hs__nand2b_2 _28511_ (.B(net374),
    .Y(_22000_),
    .A(\tholin_riscv.regs[23][2] ));
 sky130_as_sc_hs__nand3_2 _28512_ (.A(net360),
    .B(_21999_),
    .C(_22000_),
    .Y(_22001_));
 sky130_as_sc_hs__or2_2 _28513_ (.A(net374),
    .B(\tholin_riscv.regs[20][2] ),
    .Y(_22002_));
 sky130_as_sc_hs__nand2b_2 _28514_ (.B(net374),
    .Y(_22003_),
    .A(\tholin_riscv.regs[21][2] ));
 sky130_as_sc_hs__nand3_2 _28515_ (.A(net221),
    .B(_22002_),
    .C(_22003_),
    .Y(_22004_));
 sky130_as_sc_hs__nand3_2 _28516_ (.A(net347),
    .B(_22001_),
    .C(_22004_),
    .Y(_22005_));
 sky130_as_sc_hs__nand3_2 _28517_ (.A(net242),
    .B(_21998_),
    .C(_22005_),
    .Y(_22006_));
 sky130_as_sc_hs__nand3_2 _28518_ (.A(net340),
    .B(_21984_),
    .C(_21991_),
    .Y(_22007_));
 sky130_as_sc_hs__nand3_2 _28519_ (.A(net335),
    .B(_22006_),
    .C(_22007_),
    .Y(_22008_));
 sky130_as_sc_hs__or2_2 _28520_ (.A(net375),
    .B(\tholin_riscv.regs[8][2] ),
    .Y(_22009_));
 sky130_as_sc_hs__nand2b_2 _28521_ (.B(net376),
    .Y(_22010_),
    .A(\tholin_riscv.regs[9][2] ));
 sky130_as_sc_hs__nand3_2 _28522_ (.A(net224),
    .B(_22009_),
    .C(_22010_),
    .Y(_22011_));
 sky130_as_sc_hs__or2_2 _28523_ (.A(net376),
    .B(\tholin_riscv.regs[10][2] ),
    .Y(_22012_));
 sky130_as_sc_hs__nand2b_2 _28524_ (.B(net376),
    .Y(_22013_),
    .A(\tholin_riscv.regs[11][2] ));
 sky130_as_sc_hs__nand3_2 _28525_ (.A(net361),
    .B(_22012_),
    .C(_22013_),
    .Y(_22014_));
 sky130_as_sc_hs__nand3_2 _28526_ (.A(net236),
    .B(_22011_),
    .C(_22014_),
    .Y(_22015_));
 sky130_as_sc_hs__or2_2 _28527_ (.A(net375),
    .B(\tholin_riscv.regs[12][2] ),
    .Y(_22016_));
 sky130_as_sc_hs__nand2b_2 _28528_ (.B(net375),
    .Y(_22017_),
    .A(\tholin_riscv.regs[13][2] ));
 sky130_as_sc_hs__nand3_2 _28529_ (.A(net221),
    .B(_22016_),
    .C(_22017_),
    .Y(_22018_));
 sky130_as_sc_hs__or2_2 _28530_ (.A(net375),
    .B(\tholin_riscv.regs[14][2] ),
    .Y(_22019_));
 sky130_as_sc_hs__nand2b_2 _28531_ (.B(net375),
    .Y(_22020_),
    .A(\tholin_riscv.regs[15][2] ));
 sky130_as_sc_hs__nand3_2 _28532_ (.A(net361),
    .B(_22019_),
    .C(_22020_),
    .Y(_22021_));
 sky130_as_sc_hs__nand3_2 _28533_ (.A(net347),
    .B(_22018_),
    .C(_22021_),
    .Y(_22022_));
 sky130_as_sc_hs__or2_2 _28534_ (.A(net376),
    .B(\tholin_riscv.regs[0][2] ),
    .Y(_22023_));
 sky130_as_sc_hs__nand2b_2 _28535_ (.B(net376),
    .Y(_22024_),
    .A(\tholin_riscv.regs[1][2] ));
 sky130_as_sc_hs__nand3_2 _28536_ (.A(net221),
    .B(_22023_),
    .C(_22024_),
    .Y(_22025_));
 sky130_as_sc_hs__or2_2 _28537_ (.A(net377),
    .B(\tholin_riscv.regs[2][2] ),
    .Y(_22026_));
 sky130_as_sc_hs__nand2b_2 _28538_ (.B(net377),
    .Y(_22027_),
    .A(\tholin_riscv.regs[3][2] ));
 sky130_as_sc_hs__nand3_2 _28539_ (.A(net360),
    .B(_22026_),
    .C(_22027_),
    .Y(_22028_));
 sky130_as_sc_hs__nand3_2 _28540_ (.A(net236),
    .B(_22025_),
    .C(_22028_),
    .Y(_22029_));
 sky130_as_sc_hs__or2_2 _28541_ (.A(net375),
    .B(\tholin_riscv.regs[6][2] ),
    .Y(_22030_));
 sky130_as_sc_hs__nand2b_2 _28542_ (.B(net375),
    .Y(_22031_),
    .A(\tholin_riscv.regs[7][2] ));
 sky130_as_sc_hs__nand3_2 _28543_ (.A(net361),
    .B(_22030_),
    .C(_22031_),
    .Y(_22032_));
 sky130_as_sc_hs__or2_2 _28544_ (.A(net374),
    .B(\tholin_riscv.regs[4][2] ),
    .Y(_22033_));
 sky130_as_sc_hs__nand2b_2 _28545_ (.B(net374),
    .Y(_22034_),
    .A(\tholin_riscv.regs[5][2] ));
 sky130_as_sc_hs__nand3_2 _28546_ (.A(net221),
    .B(_22033_),
    .C(_22034_),
    .Y(_22035_));
 sky130_as_sc_hs__nand3_2 _28547_ (.A(net347),
    .B(_22032_),
    .C(_22035_),
    .Y(_22036_));
 sky130_as_sc_hs__nand3_2 _28548_ (.A(net242),
    .B(_22029_),
    .C(_22036_),
    .Y(_22037_));
 sky130_as_sc_hs__nand3_2 _28549_ (.A(net340),
    .B(_22015_),
    .C(_22022_),
    .Y(_22038_));
 sky130_as_sc_hs__nand3_2 _28550_ (.A(net246),
    .B(_22037_),
    .C(_22038_),
    .Y(_22039_));
 sky130_as_sc_hs__and2_2 _28551_ (.A(_22008_),
    .B(_22039_),
    .Y(_22040_));
 sky130_as_sc_hs__or2_2 _28553_ (.A(net379),
    .B(\tholin_riscv.regs[24][1] ),
    .Y(_22042_));
 sky130_as_sc_hs__nand2b_2 _28554_ (.B(net378),
    .Y(_22043_),
    .A(\tholin_riscv.regs[25][1] ));
 sky130_as_sc_hs__nand3_2 _28555_ (.A(net223),
    .B(_22042_),
    .C(_22043_),
    .Y(_22044_));
 sky130_as_sc_hs__or2_2 _28556_ (.A(net378),
    .B(\tholin_riscv.regs[26][1] ),
    .Y(_22045_));
 sky130_as_sc_hs__nand2b_2 _28557_ (.B(net378),
    .Y(_22046_),
    .A(\tholin_riscv.regs[27][1] ));
 sky130_as_sc_hs__nand3_2 _28558_ (.A(net363),
    .B(_22045_),
    .C(_22046_),
    .Y(_22047_));
 sky130_as_sc_hs__nand3_2 _28559_ (.A(net235),
    .B(_22044_),
    .C(_22047_),
    .Y(_22048_));
 sky130_as_sc_hs__or2_2 _28560_ (.A(net379),
    .B(\tholin_riscv.regs[28][1] ),
    .Y(_22049_));
 sky130_as_sc_hs__nand2b_2 _28561_ (.B(net379),
    .Y(_22050_),
    .A(\tholin_riscv.regs[29][1] ));
 sky130_as_sc_hs__nand3_2 _28562_ (.A(net223),
    .B(_22049_),
    .C(_22050_),
    .Y(_22051_));
 sky130_as_sc_hs__or2_2 _28563_ (.A(net379),
    .B(\tholin_riscv.regs[30][1] ),
    .Y(_22052_));
 sky130_as_sc_hs__nand2b_2 _28564_ (.B(net379),
    .Y(_22053_),
    .A(\tholin_riscv.regs[31][1] ));
 sky130_as_sc_hs__nand3_2 _28565_ (.A(net363),
    .B(_22052_),
    .C(_22053_),
    .Y(_22054_));
 sky130_as_sc_hs__nand3_2 _28566_ (.A(net346),
    .B(_22051_),
    .C(_22054_),
    .Y(_22055_));
 sky130_as_sc_hs__or2_2 _28567_ (.A(net378),
    .B(\tholin_riscv.regs[16][1] ),
    .Y(_22056_));
 sky130_as_sc_hs__nand2b_2 _28568_ (.B(net378),
    .Y(_22057_),
    .A(\tholin_riscv.regs[17][1] ));
 sky130_as_sc_hs__nand3_2 _28569_ (.A(net223),
    .B(_22056_),
    .C(_22057_),
    .Y(_22058_));
 sky130_as_sc_hs__or2_2 _28570_ (.A(net380),
    .B(\tholin_riscv.regs[18][1] ),
    .Y(_22059_));
 sky130_as_sc_hs__nand2b_2 _28571_ (.B(net380),
    .Y(_22060_),
    .A(\tholin_riscv.regs[19][1] ));
 sky130_as_sc_hs__nand3_2 _28572_ (.A(net363),
    .B(_22059_),
    .C(_22060_),
    .Y(_22061_));
 sky130_as_sc_hs__nand3_2 _28573_ (.A(net235),
    .B(_22058_),
    .C(_22061_),
    .Y(_22062_));
 sky130_as_sc_hs__or2_2 _28574_ (.A(net380),
    .B(\tholin_riscv.regs[22][1] ),
    .Y(_22063_));
 sky130_as_sc_hs__nand2b_2 _28575_ (.B(net380),
    .Y(_22064_),
    .A(\tholin_riscv.regs[23][1] ));
 sky130_as_sc_hs__nand3_2 _28576_ (.A(net363),
    .B(_22063_),
    .C(_22064_),
    .Y(_22065_));
 sky130_as_sc_hs__or2_2 _28577_ (.A(net380),
    .B(\tholin_riscv.regs[20][1] ),
    .Y(_22066_));
 sky130_as_sc_hs__nand2b_2 _28578_ (.B(net380),
    .Y(_22067_),
    .A(\tholin_riscv.regs[21][1] ));
 sky130_as_sc_hs__nand3_2 _28579_ (.A(net223),
    .B(_22066_),
    .C(_22067_),
    .Y(_22068_));
 sky130_as_sc_hs__nand3_2 _28580_ (.A(net346),
    .B(_22065_),
    .C(_22068_),
    .Y(_22069_));
 sky130_as_sc_hs__nand3_2 _28581_ (.A(net244),
    .B(_22062_),
    .C(_22069_),
    .Y(_22070_));
 sky130_as_sc_hs__nand3_2 _28582_ (.A(net340),
    .B(_22048_),
    .C(_22055_),
    .Y(_22071_));
 sky130_as_sc_hs__nand3_2 _28583_ (.A(net335),
    .B(_22070_),
    .C(_22071_),
    .Y(_22072_));
 sky130_as_sc_hs__or2_2 _28584_ (.A(net381),
    .B(\tholin_riscv.regs[8][1] ),
    .Y(_22073_));
 sky130_as_sc_hs__nand2b_2 _28585_ (.B(net382),
    .Y(_22074_),
    .A(\tholin_riscv.regs[9][1] ));
 sky130_as_sc_hs__nand3_2 _28586_ (.A(net222),
    .B(_22073_),
    .C(_22074_),
    .Y(_22075_));
 sky130_as_sc_hs__or2_2 _28587_ (.A(net381),
    .B(\tholin_riscv.regs[10][1] ),
    .Y(_22076_));
 sky130_as_sc_hs__nand2b_2 _28588_ (.B(net381),
    .Y(_22077_),
    .A(\tholin_riscv.regs[11][1] ));
 sky130_as_sc_hs__nand3_2 _28589_ (.A(net362),
    .B(_22076_),
    .C(_22077_),
    .Y(_22078_));
 sky130_as_sc_hs__nand3_2 _28590_ (.A(net235),
    .B(_22075_),
    .C(_22078_),
    .Y(_22079_));
 sky130_as_sc_hs__or2_2 _28591_ (.A(net380),
    .B(\tholin_riscv.regs[12][1] ),
    .Y(_22080_));
 sky130_as_sc_hs__nand2b_2 _28592_ (.B(net380),
    .Y(_22081_),
    .A(\tholin_riscv.regs[13][1] ));
 sky130_as_sc_hs__nand3_2 _28593_ (.A(net223),
    .B(_22080_),
    .C(_22081_),
    .Y(_22082_));
 sky130_as_sc_hs__or2_2 _28594_ (.A(net380),
    .B(\tholin_riscv.regs[14][1] ),
    .Y(_22083_));
 sky130_as_sc_hs__nand2b_2 _28595_ (.B(net380),
    .Y(_22084_),
    .A(\tholin_riscv.regs[15][1] ));
 sky130_as_sc_hs__nand3_2 _28596_ (.A(net362),
    .B(_22083_),
    .C(_22084_),
    .Y(_22085_));
 sky130_as_sc_hs__nand3_2 _28597_ (.A(net346),
    .B(_22082_),
    .C(_22085_),
    .Y(_22086_));
 sky130_as_sc_hs__or2_2 _28598_ (.A(net381),
    .B(\tholin_riscv.regs[0][1] ),
    .Y(_22087_));
 sky130_as_sc_hs__nand2b_2 _28599_ (.B(net381),
    .Y(_22088_),
    .A(\tholin_riscv.regs[1][1] ));
 sky130_as_sc_hs__nand3_2 _28600_ (.A(net223),
    .B(_22087_),
    .C(_22088_),
    .Y(_22089_));
 sky130_as_sc_hs__or2_2 _28601_ (.A(net381),
    .B(\tholin_riscv.regs[2][1] ),
    .Y(_22090_));
 sky130_as_sc_hs__nand2b_2 _28602_ (.B(net381),
    .Y(_22091_),
    .A(\tholin_riscv.regs[3][1] ));
 sky130_as_sc_hs__nand3_2 _28603_ (.A(net362),
    .B(_22090_),
    .C(_22091_),
    .Y(_22092_));
 sky130_as_sc_hs__nand3_2 _28604_ (.A(net235),
    .B(_22089_),
    .C(_22092_),
    .Y(_22093_));
 sky130_as_sc_hs__or2_2 _28605_ (.A(net381),
    .B(\tholin_riscv.regs[6][1] ),
    .Y(_22094_));
 sky130_as_sc_hs__nand2b_2 _28606_ (.B(net381),
    .Y(_22095_),
    .A(\tholin_riscv.regs[7][1] ));
 sky130_as_sc_hs__nand3_2 _28607_ (.A(net362),
    .B(_22094_),
    .C(_22095_),
    .Y(_22096_));
 sky130_as_sc_hs__or2_2 _28608_ (.A(net381),
    .B(\tholin_riscv.regs[4][1] ),
    .Y(_22097_));
 sky130_as_sc_hs__nand2b_2 _28609_ (.B(net381),
    .Y(_22098_),
    .A(\tholin_riscv.regs[5][1] ));
 sky130_as_sc_hs__nand3_2 _28610_ (.A(net222),
    .B(_22097_),
    .C(_22098_),
    .Y(_22099_));
 sky130_as_sc_hs__nand3_2 _28611_ (.A(net346),
    .B(_22096_),
    .C(_22099_),
    .Y(_22100_));
 sky130_as_sc_hs__nand3_2 _28612_ (.A(net242),
    .B(_22093_),
    .C(_22100_),
    .Y(_22101_));
 sky130_as_sc_hs__nand3_2 _28613_ (.A(net340),
    .B(_22079_),
    .C(_22086_),
    .Y(_22102_));
 sky130_as_sc_hs__nand3_2 _28614_ (.A(net246),
    .B(_22101_),
    .C(_22102_),
    .Y(_22103_));
 sky130_as_sc_hs__or2_2 _28616_ (.A(net374),
    .B(\tholin_riscv.regs[24][0] ),
    .Y(_22105_));
 sky130_as_sc_hs__nand2b_2 _28617_ (.B(net374),
    .Y(_22106_),
    .A(\tholin_riscv.regs[25][0] ));
 sky130_as_sc_hs__nand3_2 _28618_ (.A(net221),
    .B(_22105_),
    .C(_22106_),
    .Y(_22107_));
 sky130_as_sc_hs__or2_2 _28619_ (.A(net374),
    .B(\tholin_riscv.regs[26][0] ),
    .Y(_22108_));
 sky130_as_sc_hs__nand2b_2 _28620_ (.B(net374),
    .Y(_22109_),
    .A(\tholin_riscv.regs[27][0] ));
 sky130_as_sc_hs__nand3_2 _28621_ (.A(net360),
    .B(_22108_),
    .C(_22109_),
    .Y(_22110_));
 sky130_as_sc_hs__nand3_2 _28622_ (.A(net236),
    .B(_22107_),
    .C(_22110_),
    .Y(_22111_));
 sky130_as_sc_hs__or2_2 _28623_ (.A(net374),
    .B(\tholin_riscv.regs[28][0] ),
    .Y(_22112_));
 sky130_as_sc_hs__nand2b_2 _28624_ (.B(net374),
    .Y(_22113_),
    .A(\tholin_riscv.regs[29][0] ));
 sky130_as_sc_hs__nand3_2 _28625_ (.A(net221),
    .B(_22112_),
    .C(_22113_),
    .Y(_22114_));
 sky130_as_sc_hs__or2_2 _28626_ (.A(net382),
    .B(\tholin_riscv.regs[30][0] ),
    .Y(_22115_));
 sky130_as_sc_hs__nand2b_2 _28627_ (.B(net382),
    .Y(_22116_),
    .A(\tholin_riscv.regs[31][0] ));
 sky130_as_sc_hs__nand3_2 _28628_ (.A(net360),
    .B(_22115_),
    .C(_22116_),
    .Y(_22117_));
 sky130_as_sc_hs__nand3_2 _28629_ (.A(net347),
    .B(_22114_),
    .C(_22117_),
    .Y(_22118_));
 sky130_as_sc_hs__or2_2 _28630_ (.A(net374),
    .B(\tholin_riscv.regs[16][0] ),
    .Y(_22119_));
 sky130_as_sc_hs__nand2b_2 _28631_ (.B(net374),
    .Y(_22120_),
    .A(\tholin_riscv.regs[17][0] ));
 sky130_as_sc_hs__nand3_2 _28632_ (.A(net221),
    .B(_22119_),
    .C(_22120_),
    .Y(_22121_));
 sky130_as_sc_hs__or2_2 _28633_ (.A(net374),
    .B(\tholin_riscv.regs[18][0] ),
    .Y(_22122_));
 sky130_as_sc_hs__nand2b_2 _28634_ (.B(net374),
    .Y(_22123_),
    .A(\tholin_riscv.regs[19][0] ));
 sky130_as_sc_hs__nand3_2 _28635_ (.A(net360),
    .B(_22122_),
    .C(_22123_),
    .Y(_22124_));
 sky130_as_sc_hs__nand3_2 _28636_ (.A(net236),
    .B(_22121_),
    .C(_22124_),
    .Y(_22125_));
 sky130_as_sc_hs__or2_2 _28637_ (.A(net382),
    .B(\tholin_riscv.regs[22][0] ),
    .Y(_22126_));
 sky130_as_sc_hs__nand2b_2 _28638_ (.B(net382),
    .Y(_22127_),
    .A(\tholin_riscv.regs[23][0] ));
 sky130_as_sc_hs__nand3_2 _28639_ (.A(net360),
    .B(_22126_),
    .C(_22127_),
    .Y(_22128_));
 sky130_as_sc_hs__or2_2 _28640_ (.A(net377),
    .B(\tholin_riscv.regs[20][0] ),
    .Y(_22129_));
 sky130_as_sc_hs__nand2b_2 _28641_ (.B(net377),
    .Y(_22130_),
    .A(\tholin_riscv.regs[21][0] ));
 sky130_as_sc_hs__nand3_2 _28642_ (.A(net221),
    .B(_22129_),
    .C(_22130_),
    .Y(_22131_));
 sky130_as_sc_hs__nand3_2 _28643_ (.A(net347),
    .B(_22128_),
    .C(_22131_),
    .Y(_22132_));
 sky130_as_sc_hs__nand3_2 _28644_ (.A(net242),
    .B(_22125_),
    .C(_22132_),
    .Y(_22133_));
 sky130_as_sc_hs__nand3_2 _28645_ (.A(net340),
    .B(_22111_),
    .C(_22118_),
    .Y(_22134_));
 sky130_as_sc_hs__nand3_2 _28646_ (.A(net335),
    .B(_22133_),
    .C(_22134_),
    .Y(_22135_));
 sky130_as_sc_hs__or2_2 _28647_ (.A(net378),
    .B(\tholin_riscv.regs[8][0] ),
    .Y(_22136_));
 sky130_as_sc_hs__nand2b_2 _28648_ (.B(net378),
    .Y(_22137_),
    .A(\tholin_riscv.regs[9][0] ));
 sky130_as_sc_hs__nand3_2 _28649_ (.A(net223),
    .B(_22136_),
    .C(_22137_),
    .Y(_22138_));
 sky130_as_sc_hs__or2_2 _28650_ (.A(net378),
    .B(\tholin_riscv.regs[10][0] ),
    .Y(_22139_));
 sky130_as_sc_hs__nand2b_2 _28651_ (.B(net378),
    .Y(_22140_),
    .A(\tholin_riscv.regs[11][0] ));
 sky130_as_sc_hs__nand3_2 _28652_ (.A(net363),
    .B(_22139_),
    .C(_22140_),
    .Y(_22141_));
 sky130_as_sc_hs__nand3_2 _28653_ (.A(net235),
    .B(_22138_),
    .C(_22141_),
    .Y(_22142_));
 sky130_as_sc_hs__or2_2 _28654_ (.A(net378),
    .B(\tholin_riscv.regs[12][0] ),
    .Y(_22143_));
 sky130_as_sc_hs__nand2b_2 _28655_ (.B(net378),
    .Y(_22144_),
    .A(\tholin_riscv.regs[13][0] ));
 sky130_as_sc_hs__nand3_2 _28656_ (.A(net223),
    .B(_22143_),
    .C(_22144_),
    .Y(_22145_));
 sky130_as_sc_hs__or2_2 _28657_ (.A(net382),
    .B(\tholin_riscv.regs[14][0] ),
    .Y(_22146_));
 sky130_as_sc_hs__nand2b_2 _28658_ (.B(net382),
    .Y(_22147_),
    .A(\tholin_riscv.regs[15][0] ));
 sky130_as_sc_hs__nand3_2 _28659_ (.A(net363),
    .B(_22146_),
    .C(_22147_),
    .Y(_22148_));
 sky130_as_sc_hs__nand3_2 _28660_ (.A(net346),
    .B(_22145_),
    .C(_22148_),
    .Y(_22149_));
 sky130_as_sc_hs__or2_2 _28661_ (.A(net378),
    .B(\tholin_riscv.regs[0][0] ),
    .Y(_22150_));
 sky130_as_sc_hs__nand2b_2 _28662_ (.B(net378),
    .Y(_22151_),
    .A(\tholin_riscv.regs[1][0] ));
 sky130_as_sc_hs__nand3_2 _28663_ (.A(net223),
    .B(_22150_),
    .C(_22151_),
    .Y(_22152_));
 sky130_as_sc_hs__or2_2 _28664_ (.A(net378),
    .B(\tholin_riscv.regs[2][0] ),
    .Y(_22153_));
 sky130_as_sc_hs__nand2b_2 _28665_ (.B(net379),
    .Y(_22154_),
    .A(\tholin_riscv.regs[3][0] ));
 sky130_as_sc_hs__nand3_2 _28666_ (.A(net363),
    .B(_22153_),
    .C(_22154_),
    .Y(_22155_));
 sky130_as_sc_hs__nand3_2 _28667_ (.A(net235),
    .B(_22152_),
    .C(_22155_),
    .Y(_22156_));
 sky130_as_sc_hs__or2_2 _28668_ (.A(net382),
    .B(\tholin_riscv.regs[6][0] ),
    .Y(_22157_));
 sky130_as_sc_hs__nand2b_2 _28669_ (.B(net382),
    .Y(_22158_),
    .A(\tholin_riscv.regs[7][0] ));
 sky130_as_sc_hs__nand3_2 _28670_ (.A(net363),
    .B(_22157_),
    .C(_22158_),
    .Y(_22159_));
 sky130_as_sc_hs__or2_2 _28671_ (.A(net379),
    .B(\tholin_riscv.regs[4][0] ),
    .Y(_22160_));
 sky130_as_sc_hs__nand2b_2 _28672_ (.B(net379),
    .Y(_22161_),
    .A(\tholin_riscv.regs[5][0] ));
 sky130_as_sc_hs__nand3_2 _28673_ (.A(net223),
    .B(_22160_),
    .C(_22161_),
    .Y(_22162_));
 sky130_as_sc_hs__nand3_2 _28674_ (.A(net346),
    .B(_22159_),
    .C(_22162_),
    .Y(_22163_));
 sky130_as_sc_hs__nand3_2 _28675_ (.A(net244),
    .B(_22156_),
    .C(_22163_),
    .Y(_22164_));
 sky130_as_sc_hs__nand3_2 _28676_ (.A(net340),
    .B(_22142_),
    .C(_22149_),
    .Y(_22165_));
 sky130_as_sc_hs__nand3_2 _28677_ (.A(net246),
    .B(_22164_),
    .C(_22165_),
    .Y(_22166_));
 sky130_as_sc_hs__and2_2 _28678_ (.A(_22135_),
    .B(_22166_),
    .Y(_22167_));
 sky130_as_sc_hs__nand3_2 _28681_ (.A(_22041_),
    .B(_22104_),
    .C(_22168_),
    .Y(_22170_));
 sky130_as_sc_hs__nor2_2 _28682_ (.A(_21977_),
    .B(_22170_),
    .Y(_22171_));
 sky130_as_sc_hs__or2_2 _28683_ (.A(net395),
    .B(\tholin_riscv.regs[24][4] ),
    .Y(_22172_));
 sky130_as_sc_hs__nand3_2 _28685_ (.A(net220),
    .B(_22172_),
    .C(_22173_),
    .Y(_22174_));
 sky130_as_sc_hs__or2_2 _28686_ (.A(net395),
    .B(\tholin_riscv.regs[26][4] ),
    .Y(_22175_));
 sky130_as_sc_hs__nand3_2 _28688_ (.A(net361),
    .B(_22175_),
    .C(_22176_),
    .Y(_22177_));
 sky130_as_sc_hs__nand3_2 _28689_ (.A(net236),
    .B(_22174_),
    .C(_22177_),
    .Y(_22178_));
 sky130_as_sc_hs__or2_2 _28690_ (.A(net395),
    .B(\tholin_riscv.regs[28][4] ),
    .Y(_22179_));
 sky130_as_sc_hs__nand3_2 _28692_ (.A(net220),
    .B(_22179_),
    .C(_22180_),
    .Y(_22181_));
 sky130_as_sc_hs__or2_2 _28693_ (.A(net396),
    .B(\tholin_riscv.regs[30][4] ),
    .Y(_22182_));
 sky130_as_sc_hs__nand3_2 _28695_ (.A(net360),
    .B(_22182_),
    .C(_22183_),
    .Y(_22184_));
 sky130_as_sc_hs__nand3_2 _28696_ (.A(net347),
    .B(_22181_),
    .C(_22184_),
    .Y(_22185_));
 sky130_as_sc_hs__or2_2 _28697_ (.A(net395),
    .B(\tholin_riscv.regs[16][4] ),
    .Y(_22186_));
 sky130_as_sc_hs__nand3_2 _28699_ (.A(net220),
    .B(_22186_),
    .C(_22187_),
    .Y(_22188_));
 sky130_as_sc_hs__or2_2 _28700_ (.A(net395),
    .B(\tholin_riscv.regs[18][4] ),
    .Y(_22189_));
 sky130_as_sc_hs__nand3_2 _28702_ (.A(net361),
    .B(_22189_),
    .C(_22190_),
    .Y(_22191_));
 sky130_as_sc_hs__nand3_2 _28703_ (.A(net236),
    .B(_22188_),
    .C(_22191_),
    .Y(_22192_));
 sky130_as_sc_hs__or2_2 _28704_ (.A(net395),
    .B(\tholin_riscv.regs[22][4] ),
    .Y(_22193_));
 sky130_as_sc_hs__nand3_2 _28706_ (.A(net361),
    .B(_22193_),
    .C(_22194_),
    .Y(_22195_));
 sky130_as_sc_hs__or2_2 _28707_ (.A(net375),
    .B(\tholin_riscv.regs[20][4] ),
    .Y(_22196_));
 sky130_as_sc_hs__nand3_2 _28709_ (.A(net220),
    .B(_22196_),
    .C(_22197_),
    .Y(_22198_));
 sky130_as_sc_hs__nand3_2 _28710_ (.A(net347),
    .B(_22195_),
    .C(_22198_),
    .Y(_22199_));
 sky130_as_sc_hs__nand3_2 _28711_ (.A(net242),
    .B(_22192_),
    .C(_22199_),
    .Y(_22200_));
 sky130_as_sc_hs__nand3_2 _28712_ (.A(net340),
    .B(_22178_),
    .C(_22185_),
    .Y(_22201_));
 sky130_as_sc_hs__nand3_2 _28713_ (.A(net335),
    .B(_22200_),
    .C(_22201_),
    .Y(_22202_));
 sky130_as_sc_hs__or2_2 _28714_ (.A(net396),
    .B(\tholin_riscv.regs[8][4] ),
    .Y(_22203_));
 sky130_as_sc_hs__nand3_2 _28716_ (.A(net220),
    .B(_22203_),
    .C(_22204_),
    .Y(_22205_));
 sky130_as_sc_hs__or2_2 _28717_ (.A(net396),
    .B(\tholin_riscv.regs[10][4] ),
    .Y(_22206_));
 sky130_as_sc_hs__nand3_2 _28719_ (.A(net364),
    .B(_22206_),
    .C(_22207_),
    .Y(_22208_));
 sky130_as_sc_hs__nand3_2 _28720_ (.A(net236),
    .B(_22205_),
    .C(_22208_),
    .Y(_22209_));
 sky130_as_sc_hs__or2_2 _28721_ (.A(net396),
    .B(\tholin_riscv.regs[12][4] ),
    .Y(_22210_));
 sky130_as_sc_hs__nand3_2 _28723_ (.A(net226),
    .B(_22210_),
    .C(_22211_),
    .Y(_22212_));
 sky130_as_sc_hs__or2_2 _28724_ (.A(net396),
    .B(\tholin_riscv.regs[14][4] ),
    .Y(_22213_));
 sky130_as_sc_hs__nand3_2 _28726_ (.A(net364),
    .B(_22213_),
    .C(_22214_),
    .Y(_22215_));
 sky130_as_sc_hs__nand3_2 _28727_ (.A(net348),
    .B(_22212_),
    .C(_22215_),
    .Y(_22216_));
 sky130_as_sc_hs__or2_2 _28728_ (.A(net396),
    .B(\tholin_riscv.regs[0][4] ),
    .Y(_22217_));
 sky130_as_sc_hs__nand3_2 _28730_ (.A(net225),
    .B(_22217_),
    .C(_22218_),
    .Y(_22219_));
 sky130_as_sc_hs__or2_2 _28731_ (.A(net396),
    .B(\tholin_riscv.regs[2][4] ),
    .Y(_22220_));
 sky130_as_sc_hs__nand3_2 _28733_ (.A(net364),
    .B(_22220_),
    .C(_22221_),
    .Y(_22222_));
 sky130_as_sc_hs__nand3_2 _28734_ (.A(net237),
    .B(_22219_),
    .C(_22222_),
    .Y(_22223_));
 sky130_as_sc_hs__or2_2 _28735_ (.A(net396),
    .B(\tholin_riscv.regs[6][4] ),
    .Y(_22224_));
 sky130_as_sc_hs__nand3_2 _28737_ (.A(net364),
    .B(_22224_),
    .C(_22225_),
    .Y(_22226_));
 sky130_as_sc_hs__or2_2 _28738_ (.A(net396),
    .B(\tholin_riscv.regs[4][4] ),
    .Y(_22227_));
 sky130_as_sc_hs__nand3_2 _28740_ (.A(net220),
    .B(_22227_),
    .C(_22228_),
    .Y(_22229_));
 sky130_as_sc_hs__nand3_2 _28741_ (.A(net348),
    .B(_22226_),
    .C(_22229_),
    .Y(_22230_));
 sky130_as_sc_hs__nand3_2 _28742_ (.A(net243),
    .B(_22223_),
    .C(_22230_),
    .Y(_22231_));
 sky130_as_sc_hs__nand3_2 _28743_ (.A(net339),
    .B(_22209_),
    .C(_22216_),
    .Y(_22232_));
 sky130_as_sc_hs__nand3_2 _28744_ (.A(net246),
    .B(_22231_),
    .C(_22232_),
    .Y(_22233_));
 sky130_as_sc_hs__and2_2 _28745_ (.A(_22202_),
    .B(_22233_),
    .Y(_22234_));
 sky130_as_sc_hs__inv_2 _28746_ (.Y(_22235_),
    .A(_22234_));
 sky130_as_sc_hs__nor2_2 _28748_ (.A(_21914_),
    .B(_22234_),
    .Y(_22237_));
 sky130_as_sc_hs__or2_2 _28750_ (.A(net385),
    .B(\tholin_riscv.regs[24][7] ),
    .Y(_22239_));
 sky130_as_sc_hs__or2_2 _28751_ (.A(net203),
    .B(\tholin_riscv.regs[25][7] ),
    .Y(_22240_));
 sky130_as_sc_hs__nand3_2 _28752_ (.A(net217),
    .B(_22239_),
    .C(_22240_),
    .Y(_22241_));
 sky130_as_sc_hs__or2_2 _28753_ (.A(net385),
    .B(\tholin_riscv.regs[26][7] ),
    .Y(_22242_));
 sky130_as_sc_hs__or2_2 _28754_ (.A(net203),
    .B(\tholin_riscv.regs[27][7] ),
    .Y(_22243_));
 sky130_as_sc_hs__nand3_2 _28755_ (.A(net358),
    .B(_22242_),
    .C(_22243_),
    .Y(_22244_));
 sky130_as_sc_hs__nand3_2 _28756_ (.A(net233),
    .B(_22241_),
    .C(_22244_),
    .Y(_22245_));
 sky130_as_sc_hs__or2_2 _28757_ (.A(net384),
    .B(\tholin_riscv.regs[28][7] ),
    .Y(_22246_));
 sky130_as_sc_hs__or2_2 _28758_ (.A(net208),
    .B(\tholin_riscv.regs[29][7] ),
    .Y(_22247_));
 sky130_as_sc_hs__nand3_2 _28759_ (.A(net215),
    .B(_22246_),
    .C(_22247_),
    .Y(_22248_));
 sky130_as_sc_hs__or2_2 _28760_ (.A(net390),
    .B(\tholin_riscv.regs[30][7] ),
    .Y(_22249_));
 sky130_as_sc_hs__or2_2 _28761_ (.A(net208),
    .B(\tholin_riscv.regs[31][7] ),
    .Y(_22250_));
 sky130_as_sc_hs__nand3_2 _28762_ (.A(net355),
    .B(_22249_),
    .C(_22250_),
    .Y(_22251_));
 sky130_as_sc_hs__nand3_2 _28763_ (.A(net344),
    .B(_22248_),
    .C(_22251_),
    .Y(_22252_));
 sky130_as_sc_hs__or2_2 _28764_ (.A(net384),
    .B(\tholin_riscv.regs[16][7] ),
    .Y(_22253_));
 sky130_as_sc_hs__or2_2 _28765_ (.A(net203),
    .B(\tholin_riscv.regs[17][7] ),
    .Y(_22254_));
 sky130_as_sc_hs__nand3_2 _28766_ (.A(net215),
    .B(_22253_),
    .C(_22254_),
    .Y(_22255_));
 sky130_as_sc_hs__or2_2 _28767_ (.A(net385),
    .B(\tholin_riscv.regs[18][7] ),
    .Y(_22256_));
 sky130_as_sc_hs__or2_2 _28768_ (.A(net210),
    .B(\tholin_riscv.regs[19][7] ),
    .Y(_22257_));
 sky130_as_sc_hs__nand3_2 _28769_ (.A(net355),
    .B(_22256_),
    .C(_22257_),
    .Y(_22258_));
 sky130_as_sc_hs__nand3_2 _28770_ (.A(net233),
    .B(_22255_),
    .C(_22258_),
    .Y(_22259_));
 sky130_as_sc_hs__or2_2 _28771_ (.A(net384),
    .B(\tholin_riscv.regs[22][7] ),
    .Y(_22260_));
 sky130_as_sc_hs__or2_2 _28772_ (.A(net203),
    .B(\tholin_riscv.regs[23][7] ),
    .Y(_22261_));
 sky130_as_sc_hs__nand3_2 _28773_ (.A(net355),
    .B(_22260_),
    .C(_22261_),
    .Y(_22262_));
 sky130_as_sc_hs__or2_2 _28774_ (.A(net384),
    .B(\tholin_riscv.regs[20][7] ),
    .Y(_22263_));
 sky130_as_sc_hs__or2_2 _28775_ (.A(net203),
    .B(\tholin_riscv.regs[21][7] ),
    .Y(_22264_));
 sky130_as_sc_hs__nand3_2 _28776_ (.A(net215),
    .B(_22263_),
    .C(_22264_),
    .Y(_22265_));
 sky130_as_sc_hs__nand3_2 _28777_ (.A(net344),
    .B(_22262_),
    .C(_22265_),
    .Y(_22266_));
 sky130_as_sc_hs__nand3_2 _28778_ (.A(net241),
    .B(_22259_),
    .C(_22266_),
    .Y(_22267_));
 sky130_as_sc_hs__nand3_2 _28779_ (.A(net338),
    .B(_22245_),
    .C(_22252_),
    .Y(_22268_));
 sky130_as_sc_hs__nand3_2 _28780_ (.A(net336),
    .B(_22267_),
    .C(_22268_),
    .Y(_22269_));
 sky130_as_sc_hs__or2_2 _28781_ (.A(net385),
    .B(\tholin_riscv.regs[8][7] ),
    .Y(_22270_));
 sky130_as_sc_hs__or2_2 _28782_ (.A(net209),
    .B(\tholin_riscv.regs[9][7] ),
    .Y(_22271_));
 sky130_as_sc_hs__nand3_2 _28783_ (.A(net217),
    .B(_22270_),
    .C(_22271_),
    .Y(_22272_));
 sky130_as_sc_hs__or2_2 _28784_ (.A(net385),
    .B(\tholin_riscv.regs[10][7] ),
    .Y(_22273_));
 sky130_as_sc_hs__or2_2 _28785_ (.A(net205),
    .B(\tholin_riscv.regs[11][7] ),
    .Y(_22274_));
 sky130_as_sc_hs__nand3_2 _28786_ (.A(net358),
    .B(_22273_),
    .C(_22274_),
    .Y(_22275_));
 sky130_as_sc_hs__nand3_2 _28787_ (.A(net234),
    .B(_22272_),
    .C(_22275_),
    .Y(_22276_));
 sky130_as_sc_hs__or2_2 _28788_ (.A(net390),
    .B(\tholin_riscv.regs[12][7] ),
    .Y(_22277_));
 sky130_as_sc_hs__or2_2 _28789_ (.A(net209),
    .B(\tholin_riscv.regs[13][7] ),
    .Y(_22278_));
 sky130_as_sc_hs__nand3_2 _28790_ (.A(net217),
    .B(_22277_),
    .C(_22278_),
    .Y(_22279_));
 sky130_as_sc_hs__or2_2 _28791_ (.A(net385),
    .B(\tholin_riscv.regs[14][7] ),
    .Y(_22280_));
 sky130_as_sc_hs__or2_2 _28792_ (.A(net209),
    .B(\tholin_riscv.regs[15][7] ),
    .Y(_22281_));
 sky130_as_sc_hs__nand3_2 _28793_ (.A(net358),
    .B(_22280_),
    .C(_22281_),
    .Y(_22282_));
 sky130_as_sc_hs__nand3_2 _28794_ (.A(net345),
    .B(_22279_),
    .C(_22282_),
    .Y(_22283_));
 sky130_as_sc_hs__or2_2 _28795_ (.A(net390),
    .B(\tholin_riscv.regs[0][7] ),
    .Y(_22284_));
 sky130_as_sc_hs__or2_2 _28796_ (.A(net209),
    .B(\tholin_riscv.regs[1][7] ),
    .Y(_22285_));
 sky130_as_sc_hs__nand3_2 _28797_ (.A(net217),
    .B(_22284_),
    .C(_22285_),
    .Y(_22286_));
 sky130_as_sc_hs__or2_2 _28798_ (.A(net385),
    .B(\tholin_riscv.regs[2][7] ),
    .Y(_22287_));
 sky130_as_sc_hs__or2_2 _28799_ (.A(net209),
    .B(\tholin_riscv.regs[3][7] ),
    .Y(_22288_));
 sky130_as_sc_hs__nand3_2 _28800_ (.A(net358),
    .B(_22287_),
    .C(_22288_),
    .Y(_22289_));
 sky130_as_sc_hs__nand3_2 _28801_ (.A(net234),
    .B(_22286_),
    .C(_22289_),
    .Y(_22290_));
 sky130_as_sc_hs__or2_2 _28802_ (.A(net390),
    .B(\tholin_riscv.regs[6][7] ),
    .Y(_22291_));
 sky130_as_sc_hs__or2_2 _28803_ (.A(net209),
    .B(\tholin_riscv.regs[7][7] ),
    .Y(_22292_));
 sky130_as_sc_hs__nand3_2 _28804_ (.A(net357),
    .B(_22291_),
    .C(_22292_),
    .Y(_22293_));
 sky130_as_sc_hs__or2_2 _28805_ (.A(net390),
    .B(\tholin_riscv.regs[4][7] ),
    .Y(_22294_));
 sky130_as_sc_hs__or2_2 _28806_ (.A(net209),
    .B(\tholin_riscv.regs[5][7] ),
    .Y(_22295_));
 sky130_as_sc_hs__nand3_2 _28807_ (.A(net217),
    .B(_22294_),
    .C(_22295_),
    .Y(_22296_));
 sky130_as_sc_hs__nand3_2 _28808_ (.A(net345),
    .B(_22293_),
    .C(_22296_),
    .Y(_22297_));
 sky130_as_sc_hs__nand3_2 _28809_ (.A(net241),
    .B(_22290_),
    .C(_22297_),
    .Y(_22298_));
 sky130_as_sc_hs__nand3_2 _28810_ (.A(net338),
    .B(_22276_),
    .C(_22283_),
    .Y(_22299_));
 sky130_as_sc_hs__nand3_2 _28811_ (.A(net245),
    .B(_22298_),
    .C(_22299_),
    .Y(_22300_));
 sky130_as_sc_hs__and2_2 _28812_ (.A(_22269_),
    .B(_22300_),
    .Y(_22301_));
 sky130_as_sc_hs__or2_2 _28813_ (.A(net386),
    .B(\tholin_riscv.regs[24][6] ),
    .Y(_22302_));
 sky130_as_sc_hs__or2_2 _28814_ (.A(net204),
    .B(\tholin_riscv.regs[25][6] ),
    .Y(_22303_));
 sky130_as_sc_hs__nand3_2 _28815_ (.A(net214),
    .B(_22302_),
    .C(_22303_),
    .Y(_22304_));
 sky130_as_sc_hs__or2_2 _28816_ (.A(net375),
    .B(\tholin_riscv.regs[26][6] ),
    .Y(_22305_));
 sky130_as_sc_hs__or2_2 _28817_ (.A(net206),
    .B(\tholin_riscv.regs[27][6] ),
    .Y(_22306_));
 sky130_as_sc_hs__nand3_2 _28818_ (.A(net354),
    .B(_22305_),
    .C(_22306_),
    .Y(_22307_));
 sky130_as_sc_hs__nand3_2 _28819_ (.A(_19483_),
    .B(_22304_),
    .C(_22307_),
    .Y(_22308_));
 sky130_as_sc_hs__or2_2 _28820_ (.A(net395),
    .B(\tholin_riscv.regs[28][6] ),
    .Y(_22309_));
 sky130_as_sc_hs__or2_2 _28821_ (.A(net204),
    .B(\tholin_riscv.regs[29][6] ),
    .Y(_22310_));
 sky130_as_sc_hs__nand3_2 _28822_ (.A(net220),
    .B(_22309_),
    .C(_22310_),
    .Y(_22311_));
 sky130_as_sc_hs__or2_2 _28823_ (.A(net395),
    .B(\tholin_riscv.regs[30][6] ),
    .Y(_22312_));
 sky130_as_sc_hs__or2_2 _28824_ (.A(net204),
    .B(\tholin_riscv.regs[31][6] ),
    .Y(_22313_));
 sky130_as_sc_hs__nand3_2 _28825_ (.A(net361),
    .B(_22312_),
    .C(_22313_),
    .Y(_22314_));
 sky130_as_sc_hs__nand3_2 _28826_ (.A(net347),
    .B(_22311_),
    .C(_22314_),
    .Y(_22315_));
 sky130_as_sc_hs__or2_2 _28827_ (.A(net386),
    .B(\tholin_riscv.regs[16][6] ),
    .Y(_22316_));
 sky130_as_sc_hs__or2_2 _28828_ (.A(net204),
    .B(\tholin_riscv.regs[17][6] ),
    .Y(_22317_));
 sky130_as_sc_hs__nand3_2 _28829_ (.A(net214),
    .B(_22316_),
    .C(_22317_),
    .Y(_22318_));
 sky130_as_sc_hs__or2_2 _28830_ (.A(net386),
    .B(\tholin_riscv.regs[18][6] ),
    .Y(_22319_));
 sky130_as_sc_hs__or2_2 _28831_ (.A(net204),
    .B(\tholin_riscv.regs[19][6] ),
    .Y(_22320_));
 sky130_as_sc_hs__nand3_2 _28832_ (.A(net354),
    .B(_22319_),
    .C(_22320_),
    .Y(_22321_));
 sky130_as_sc_hs__nand3_2 _28833_ (.A(net232),
    .B(_22318_),
    .C(_22321_),
    .Y(_22322_));
 sky130_as_sc_hs__or2_2 _28834_ (.A(net386),
    .B(\tholin_riscv.regs[22][6] ),
    .Y(_22323_));
 sky130_as_sc_hs__or2_2 _28835_ (.A(net206),
    .B(\tholin_riscv.regs[23][6] ),
    .Y(_22324_));
 sky130_as_sc_hs__nand3_2 _28836_ (.A(net354),
    .B(_22323_),
    .C(_22324_),
    .Y(_22325_));
 sky130_as_sc_hs__or2_2 _28837_ (.A(net395),
    .B(\tholin_riscv.regs[20][6] ),
    .Y(_22326_));
 sky130_as_sc_hs__or2_2 _28838_ (.A(net206),
    .B(\tholin_riscv.regs[21][6] ),
    .Y(_22327_));
 sky130_as_sc_hs__nand3_2 _28839_ (.A(net220),
    .B(_22326_),
    .C(_22327_),
    .Y(_22328_));
 sky130_as_sc_hs__nand3_2 _28840_ (.A(net342),
    .B(_22325_),
    .C(_22328_),
    .Y(_22329_));
 sky130_as_sc_hs__nand3_2 _28841_ (.A(net242),
    .B(_22322_),
    .C(_22329_),
    .Y(_22330_));
 sky130_as_sc_hs__nand3_2 _28842_ (.A(net337),
    .B(_22308_),
    .C(_22315_),
    .Y(_22331_));
 sky130_as_sc_hs__nand3_2 _28843_ (.A(net335),
    .B(_22330_),
    .C(_22331_),
    .Y(_22332_));
 sky130_as_sc_hs__or2_2 _28844_ (.A(net395),
    .B(\tholin_riscv.regs[8][6] ),
    .Y(_22333_));
 sky130_as_sc_hs__or2_2 _28845_ (.A(net204),
    .B(\tholin_riscv.regs[9][6] ),
    .Y(_22334_));
 sky130_as_sc_hs__nand3_2 _28846_ (.A(net220),
    .B(_22333_),
    .C(_22334_),
    .Y(_22335_));
 sky130_as_sc_hs__or2_2 _28847_ (.A(net395),
    .B(\tholin_riscv.regs[10][6] ),
    .Y(_22336_));
 sky130_as_sc_hs__or2_2 _28848_ (.A(net204),
    .B(\tholin_riscv.regs[11][6] ),
    .Y(_22337_));
 sky130_as_sc_hs__nand3_2 _28849_ (.A(net361),
    .B(_22336_),
    .C(_22337_),
    .Y(_22338_));
 sky130_as_sc_hs__nand3_2 _28850_ (.A(net236),
    .B(_22335_),
    .C(_22338_),
    .Y(_22339_));
 sky130_as_sc_hs__or2_2 _28851_ (.A(net395),
    .B(\tholin_riscv.regs[12][6] ),
    .Y(_22340_));
 sky130_as_sc_hs__or2_2 _28852_ (.A(net206),
    .B(\tholin_riscv.regs[13][6] ),
    .Y(_22341_));
 sky130_as_sc_hs__nand3_2 _28853_ (.A(net220),
    .B(_22340_),
    .C(_22341_),
    .Y(_22342_));
 sky130_as_sc_hs__or2_2 _28854_ (.A(net395),
    .B(\tholin_riscv.regs[14][6] ),
    .Y(_22343_));
 sky130_as_sc_hs__or2_2 _28855_ (.A(net206),
    .B(\tholin_riscv.regs[15][6] ),
    .Y(_22344_));
 sky130_as_sc_hs__nand3_2 _28856_ (.A(net360),
    .B(_22343_),
    .C(_22344_),
    .Y(_22345_));
 sky130_as_sc_hs__nand3_2 _28857_ (.A(net347),
    .B(_22342_),
    .C(_22345_),
    .Y(_22346_));
 sky130_as_sc_hs__or2_2 _28858_ (.A(net395),
    .B(\tholin_riscv.regs[0][6] ),
    .Y(_22347_));
 sky130_as_sc_hs__or2_2 _28859_ (.A(net206),
    .B(\tholin_riscv.regs[1][6] ),
    .Y(_22348_));
 sky130_as_sc_hs__nand3_2 _28860_ (.A(net220),
    .B(_22347_),
    .C(_22348_),
    .Y(_22349_));
 sky130_as_sc_hs__or2_2 _28861_ (.A(net395),
    .B(\tholin_riscv.regs[2][6] ),
    .Y(_22350_));
 sky130_as_sc_hs__or2_2 _28862_ (.A(net206),
    .B(\tholin_riscv.regs[3][6] ),
    .Y(_22351_));
 sky130_as_sc_hs__nand3_2 _28863_ (.A(net365),
    .B(_22350_),
    .C(_22351_),
    .Y(_22352_));
 sky130_as_sc_hs__nand3_2 _28864_ (.A(net236),
    .B(_22349_),
    .C(_22352_),
    .Y(_22353_));
 sky130_as_sc_hs__or2_2 _28865_ (.A(net396),
    .B(\tholin_riscv.regs[6][6] ),
    .Y(_22354_));
 sky130_as_sc_hs__or2_2 _28866_ (.A(net206),
    .B(\tholin_riscv.regs[7][6] ),
    .Y(_22355_));
 sky130_as_sc_hs__nand3_2 _28867_ (.A(net365),
    .B(_22354_),
    .C(_22355_),
    .Y(_22356_));
 sky130_as_sc_hs__or2_2 _28868_ (.A(net396),
    .B(\tholin_riscv.regs[4][6] ),
    .Y(_22357_));
 sky130_as_sc_hs__or2_2 _28869_ (.A(net206),
    .B(\tholin_riscv.regs[5][6] ),
    .Y(_22358_));
 sky130_as_sc_hs__nand3_2 _28870_ (.A(net225),
    .B(_22357_),
    .C(_22358_),
    .Y(_22359_));
 sky130_as_sc_hs__nand3_2 _28871_ (.A(net348),
    .B(_22356_),
    .C(_22359_),
    .Y(_22360_));
 sky130_as_sc_hs__nand3_2 _28872_ (.A(net242),
    .B(_22353_),
    .C(_22360_),
    .Y(_22361_));
 sky130_as_sc_hs__nand3_2 _28873_ (.A(net340),
    .B(_22339_),
    .C(_22346_),
    .Y(_22362_));
 sky130_as_sc_hs__nand3_2 _28874_ (.A(net246),
    .B(_22361_),
    .C(_22362_),
    .Y(_22363_));
 sky130_as_sc_hs__and2_2 _28875_ (.A(_22332_),
    .B(_22363_),
    .Y(_22364_));
 sky130_as_sc_hs__inv_2 _28876_ (.Y(_22365_),
    .A(_22364_));
 sky130_as_sc_hs__nor2_2 _28877_ (.A(_22301_),
    .B(_22364_),
    .Y(_22366_));
 sky130_as_sc_hs__nand3_2 _28878_ (.A(_22171_),
    .B(_22237_),
    .C(_22366_),
    .Y(_22367_));
 sky130_as_sc_hs__or2_2 _28879_ (.A(net387),
    .B(\tholin_riscv.regs[24][11] ),
    .Y(_22368_));
 sky130_as_sc_hs__nand2b_2 _28880_ (.B(net387),
    .Y(_22369_),
    .A(\tholin_riscv.regs[25][11] ));
 sky130_as_sc_hs__nand3_2 _28881_ (.A(net216),
    .B(_22368_),
    .C(_22369_),
    .Y(_22370_));
 sky130_as_sc_hs__or2_2 _28882_ (.A(net388),
    .B(\tholin_riscv.regs[26][11] ),
    .Y(_22371_));
 sky130_as_sc_hs__nand2b_2 _28883_ (.B(net387),
    .Y(_22372_),
    .A(\tholin_riscv.regs[27][11] ));
 sky130_as_sc_hs__nand3_2 _28884_ (.A(net356),
    .B(_22371_),
    .C(_22372_),
    .Y(_22373_));
 sky130_as_sc_hs__nand3_2 _28885_ (.A(net233),
    .B(_22370_),
    .C(_22373_),
    .Y(_22374_));
 sky130_as_sc_hs__or2_2 _28886_ (.A(net387),
    .B(\tholin_riscv.regs[28][11] ),
    .Y(_22375_));
 sky130_as_sc_hs__nand2b_2 _28887_ (.B(net387),
    .Y(_22376_),
    .A(\tholin_riscv.regs[29][11] ));
 sky130_as_sc_hs__nand3_2 _28888_ (.A(net216),
    .B(_22375_),
    .C(_22376_),
    .Y(_22377_));
 sky130_as_sc_hs__or2_2 _28889_ (.A(net394),
    .B(\tholin_riscv.regs[30][11] ),
    .Y(_22378_));
 sky130_as_sc_hs__nand2b_2 _28890_ (.B(net394),
    .Y(_22379_),
    .A(\tholin_riscv.regs[31][11] ));
 sky130_as_sc_hs__nand3_2 _28891_ (.A(net356),
    .B(_22378_),
    .C(_22379_),
    .Y(_22380_));
 sky130_as_sc_hs__nand3_2 _28892_ (.A(net344),
    .B(_22377_),
    .C(_22380_),
    .Y(_22381_));
 sky130_as_sc_hs__or2_2 _28893_ (.A(net384),
    .B(\tholin_riscv.regs[16][11] ),
    .Y(_22382_));
 sky130_as_sc_hs__nand2b_2 _28894_ (.B(net387),
    .Y(_22383_),
    .A(\tholin_riscv.regs[17][11] ));
 sky130_as_sc_hs__nand3_2 _28895_ (.A(net215),
    .B(_22382_),
    .C(_22383_),
    .Y(_22384_));
 sky130_as_sc_hs__or2_2 _28896_ (.A(net387),
    .B(\tholin_riscv.regs[18][11] ),
    .Y(_22385_));
 sky130_as_sc_hs__nand2b_2 _28897_ (.B(net387),
    .Y(_22386_),
    .A(\tholin_riscv.regs[19][11] ));
 sky130_as_sc_hs__nand3_2 _28898_ (.A(net355),
    .B(_22385_),
    .C(_22386_),
    .Y(_22387_));
 sky130_as_sc_hs__nand3_2 _28899_ (.A(net233),
    .B(_22384_),
    .C(_22387_),
    .Y(_22388_));
 sky130_as_sc_hs__or2_2 _28900_ (.A(net387),
    .B(\tholin_riscv.regs[22][11] ),
    .Y(_22389_));
 sky130_as_sc_hs__nand2b_2 _28901_ (.B(net387),
    .Y(_22390_),
    .A(\tholin_riscv.regs[23][11] ));
 sky130_as_sc_hs__nand3_2 _28902_ (.A(net355),
    .B(_22389_),
    .C(_22390_),
    .Y(_22391_));
 sky130_as_sc_hs__or2_2 _28903_ (.A(net387),
    .B(\tholin_riscv.regs[20][11] ),
    .Y(_22392_));
 sky130_as_sc_hs__nand2b_2 _28904_ (.B(net387),
    .Y(_22393_),
    .A(\tholin_riscv.regs[21][11] ));
 sky130_as_sc_hs__nand3_2 _28905_ (.A(net215),
    .B(_22392_),
    .C(_22393_),
    .Y(_22394_));
 sky130_as_sc_hs__nand3_2 _28906_ (.A(net344),
    .B(_22391_),
    .C(_22394_),
    .Y(_22395_));
 sky130_as_sc_hs__nand3_2 _28907_ (.A(net240),
    .B(_22388_),
    .C(_22395_),
    .Y(_22396_));
 sky130_as_sc_hs__nand3_2 _28908_ (.A(net338),
    .B(_22374_),
    .C(_22381_),
    .Y(_22397_));
 sky130_as_sc_hs__nand3_2 _28909_ (.A(net336),
    .B(_22396_),
    .C(_22397_),
    .Y(_22398_));
 sky130_as_sc_hs__or2_2 _28910_ (.A(net390),
    .B(\tholin_riscv.regs[8][11] ),
    .Y(_22399_));
 sky130_as_sc_hs__nand2b_2 _28911_ (.B(net390),
    .Y(_22400_),
    .A(\tholin_riscv.regs[9][11] ));
 sky130_as_sc_hs__nand3_2 _28912_ (.A(net218),
    .B(_22399_),
    .C(_22400_),
    .Y(_22401_));
 sky130_as_sc_hs__or2_2 _28913_ (.A(net393),
    .B(\tholin_riscv.regs[10][11] ),
    .Y(_22402_));
 sky130_as_sc_hs__nand2b_2 _28914_ (.B(net393),
    .Y(_22403_),
    .A(\tholin_riscv.regs[11][11] ));
 sky130_as_sc_hs__nand3_2 _28915_ (.A(net357),
    .B(_22402_),
    .C(_22403_),
    .Y(_22404_));
 sky130_as_sc_hs__nand3_2 _28916_ (.A(net234),
    .B(_22401_),
    .C(_22404_),
    .Y(_22405_));
 sky130_as_sc_hs__or2_2 _28917_ (.A(net390),
    .B(\tholin_riscv.regs[12][11] ),
    .Y(_22406_));
 sky130_as_sc_hs__nand2b_2 _28918_ (.B(net390),
    .Y(_22407_),
    .A(\tholin_riscv.regs[13][11] ));
 sky130_as_sc_hs__nand3_2 _28919_ (.A(net218),
    .B(_22406_),
    .C(_22407_),
    .Y(_22408_));
 sky130_as_sc_hs__or2_2 _28920_ (.A(net390),
    .B(\tholin_riscv.regs[14][11] ),
    .Y(_22409_));
 sky130_as_sc_hs__nand2b_2 _28921_ (.B(net390),
    .Y(_22410_),
    .A(\tholin_riscv.regs[15][11] ));
 sky130_as_sc_hs__nand3_2 _28922_ (.A(net357),
    .B(_22409_),
    .C(_22410_),
    .Y(_22411_));
 sky130_as_sc_hs__nand3_2 _28923_ (.A(net345),
    .B(_22408_),
    .C(_22411_),
    .Y(_22412_));
 sky130_as_sc_hs__or2_2 _28924_ (.A(net387),
    .B(\tholin_riscv.regs[0][11] ),
    .Y(_22413_));
 sky130_as_sc_hs__nand2b_2 _28925_ (.B(net387),
    .Y(_22414_),
    .A(\tholin_riscv.regs[1][11] ));
 sky130_as_sc_hs__nand3_2 _28926_ (.A(net215),
    .B(_22413_),
    .C(_22414_),
    .Y(_22415_));
 sky130_as_sc_hs__or2_2 _28927_ (.A(net387),
    .B(\tholin_riscv.regs[2][11] ),
    .Y(_22416_));
 sky130_as_sc_hs__nand2b_2 _28928_ (.B(net388),
    .Y(_22417_),
    .A(\tholin_riscv.regs[3][11] ));
 sky130_as_sc_hs__nand3_2 _28929_ (.A(net355),
    .B(_22416_),
    .C(_22417_),
    .Y(_22418_));
 sky130_as_sc_hs__nand3_2 _28930_ (.A(net233),
    .B(_22415_),
    .C(_22418_),
    .Y(_22419_));
 sky130_as_sc_hs__or2_2 _28931_ (.A(net388),
    .B(\tholin_riscv.regs[6][11] ),
    .Y(_22420_));
 sky130_as_sc_hs__nand2b_2 _28932_ (.B(net388),
    .Y(_22421_),
    .A(\tholin_riscv.regs[7][11] ));
 sky130_as_sc_hs__nand3_2 _28933_ (.A(net356),
    .B(_22420_),
    .C(_22421_),
    .Y(_22422_));
 sky130_as_sc_hs__or2_2 _28934_ (.A(net388),
    .B(\tholin_riscv.regs[4][11] ),
    .Y(_22423_));
 sky130_as_sc_hs__nand2b_2 _28935_ (.B(net387),
    .Y(_22424_),
    .A(\tholin_riscv.regs[5][11] ));
 sky130_as_sc_hs__nand3_2 _28936_ (.A(net216),
    .B(_22423_),
    .C(_22424_),
    .Y(_22425_));
 sky130_as_sc_hs__nand3_2 _28937_ (.A(net344),
    .B(_22422_),
    .C(_22425_),
    .Y(_22426_));
 sky130_as_sc_hs__nand3_2 _28938_ (.A(net241),
    .B(_22419_),
    .C(_22426_),
    .Y(_22427_));
 sky130_as_sc_hs__nand3_2 _28939_ (.A(net338),
    .B(_22405_),
    .C(_22412_),
    .Y(_22428_));
 sky130_as_sc_hs__nand3_2 _28940_ (.A(net245),
    .B(_22427_),
    .C(_22428_),
    .Y(_22429_));
 sky130_as_sc_hs__and2_2 _28941_ (.A(_22398_),
    .B(_22429_),
    .Y(_22430_));
 sky130_as_sc_hs__or2_2 _28942_ (.A(net392),
    .B(\tholin_riscv.regs[24][10] ),
    .Y(_22431_));
 sky130_as_sc_hs__nand2b_2 _28943_ (.B(net392),
    .Y(_22432_),
    .A(\tholin_riscv.regs[25][10] ));
 sky130_as_sc_hs__nand3_2 _28944_ (.A(net217),
    .B(_22431_),
    .C(_22432_),
    .Y(_22433_));
 sky130_as_sc_hs__or2_2 _28945_ (.A(net394),
    .B(\tholin_riscv.regs[26][10] ),
    .Y(_22434_));
 sky130_as_sc_hs__nand2b_2 _28946_ (.B(net392),
    .Y(_22435_),
    .A(\tholin_riscv.regs[27][10] ));
 sky130_as_sc_hs__nand3_2 _28947_ (.A(net357),
    .B(_22434_),
    .C(_22435_),
    .Y(_22436_));
 sky130_as_sc_hs__nand3_2 _28948_ (.A(net234),
    .B(_22433_),
    .C(_22436_),
    .Y(_22437_));
 sky130_as_sc_hs__or2_2 _28949_ (.A(net392),
    .B(\tholin_riscv.regs[28][10] ),
    .Y(_22438_));
 sky130_as_sc_hs__nand2b_2 _28950_ (.B(net392),
    .Y(_22439_),
    .A(\tholin_riscv.regs[29][10] ));
 sky130_as_sc_hs__nand3_2 _28951_ (.A(net218),
    .B(_22438_),
    .C(_22439_),
    .Y(_22440_));
 sky130_as_sc_hs__or2_2 _28952_ (.A(net392),
    .B(\tholin_riscv.regs[30][10] ),
    .Y(_22441_));
 sky130_as_sc_hs__nand2b_2 _28953_ (.B(net392),
    .Y(_22442_),
    .A(\tholin_riscv.regs[31][10] ));
 sky130_as_sc_hs__nand3_2 _28954_ (.A(net357),
    .B(_22441_),
    .C(_22442_),
    .Y(_22443_));
 sky130_as_sc_hs__nand3_2 _28955_ (.A(net345),
    .B(_22440_),
    .C(_22443_),
    .Y(_22444_));
 sky130_as_sc_hs__or2_2 _28956_ (.A(net393),
    .B(\tholin_riscv.regs[16][10] ),
    .Y(_22445_));
 sky130_as_sc_hs__nand2b_2 _28957_ (.B(net393),
    .Y(_22446_),
    .A(\tholin_riscv.regs[17][10] ));
 sky130_as_sc_hs__nand3_2 _28958_ (.A(net218),
    .B(_22445_),
    .C(_22446_),
    .Y(_22447_));
 sky130_as_sc_hs__or2_2 _28959_ (.A(net393),
    .B(\tholin_riscv.regs[18][10] ),
    .Y(_22448_));
 sky130_as_sc_hs__nand2b_2 _28960_ (.B(net393),
    .Y(_22449_),
    .A(\tholin_riscv.regs[19][10] ));
 sky130_as_sc_hs__nand3_2 _28961_ (.A(net357),
    .B(_22448_),
    .C(_22449_),
    .Y(_22450_));
 sky130_as_sc_hs__nand3_2 _28962_ (.A(net234),
    .B(_22447_),
    .C(_22450_),
    .Y(_22451_));
 sky130_as_sc_hs__or2_2 _28963_ (.A(net393),
    .B(\tholin_riscv.regs[22][10] ),
    .Y(_22452_));
 sky130_as_sc_hs__nand2b_2 _28964_ (.B(net393),
    .Y(_22453_),
    .A(\tholin_riscv.regs[23][10] ));
 sky130_as_sc_hs__nand3_2 _28965_ (.A(net357),
    .B(_22452_),
    .C(_22453_),
    .Y(_22454_));
 sky130_as_sc_hs__or2_2 _28966_ (.A(net390),
    .B(\tholin_riscv.regs[20][10] ),
    .Y(_22455_));
 sky130_as_sc_hs__nand2b_2 _28967_ (.B(net390),
    .Y(_22456_),
    .A(\tholin_riscv.regs[21][10] ));
 sky130_as_sc_hs__nand3_2 _28968_ (.A(net218),
    .B(_22455_),
    .C(_22456_),
    .Y(_22457_));
 sky130_as_sc_hs__nand3_2 _28969_ (.A(net345),
    .B(_22454_),
    .C(_22457_),
    .Y(_22458_));
 sky130_as_sc_hs__nand3_2 _28970_ (.A(net240),
    .B(_22451_),
    .C(_22458_),
    .Y(_22459_));
 sky130_as_sc_hs__nand3_2 _28971_ (.A(net338),
    .B(_22437_),
    .C(_22444_),
    .Y(_22460_));
 sky130_as_sc_hs__nand3_2 _28972_ (.A(net336),
    .B(_22459_),
    .C(_22460_),
    .Y(_22461_));
 sky130_as_sc_hs__or2_2 _28973_ (.A(net391),
    .B(\tholin_riscv.regs[8][10] ),
    .Y(_22462_));
 sky130_as_sc_hs__nand2b_2 _28974_ (.B(net391),
    .Y(_22463_),
    .A(\tholin_riscv.regs[9][10] ));
 sky130_as_sc_hs__nand3_2 _28975_ (.A(net217),
    .B(_22462_),
    .C(_22463_),
    .Y(_22464_));
 sky130_as_sc_hs__or2_2 _28976_ (.A(net390),
    .B(\tholin_riscv.regs[10][10] ),
    .Y(_22465_));
 sky130_as_sc_hs__nand2b_2 _28977_ (.B(net391),
    .Y(_22466_),
    .A(\tholin_riscv.regs[11][10] ));
 sky130_as_sc_hs__nand3_2 _28978_ (.A(net357),
    .B(_22465_),
    .C(_22466_),
    .Y(_22467_));
 sky130_as_sc_hs__nand3_2 _28979_ (.A(net234),
    .B(_22464_),
    .C(_22467_),
    .Y(_22468_));
 sky130_as_sc_hs__or2_2 _28980_ (.A(net391),
    .B(\tholin_riscv.regs[12][10] ),
    .Y(_22469_));
 sky130_as_sc_hs__nand2b_2 _28981_ (.B(net391),
    .Y(_22470_),
    .A(\tholin_riscv.regs[13][10] ));
 sky130_as_sc_hs__nand3_2 _28982_ (.A(net217),
    .B(_22469_),
    .C(_22470_),
    .Y(_22471_));
 sky130_as_sc_hs__or2_2 _28983_ (.A(net392),
    .B(\tholin_riscv.regs[14][10] ),
    .Y(_22472_));
 sky130_as_sc_hs__nand2b_2 _28984_ (.B(net392),
    .Y(_22473_),
    .A(\tholin_riscv.regs[15][10] ));
 sky130_as_sc_hs__nand3_2 _28985_ (.A(net357),
    .B(_22472_),
    .C(_22473_),
    .Y(_22474_));
 sky130_as_sc_hs__nand3_2 _28986_ (.A(net345),
    .B(_22471_),
    .C(_22474_),
    .Y(_22475_));
 sky130_as_sc_hs__or2_2 _28987_ (.A(net391),
    .B(\tholin_riscv.regs[0][10] ),
    .Y(_22476_));
 sky130_as_sc_hs__nand2b_2 _28988_ (.B(net390),
    .Y(_22477_),
    .A(\tholin_riscv.regs[1][10] ));
 sky130_as_sc_hs__nand3_2 _28989_ (.A(net217),
    .B(_22476_),
    .C(_22477_),
    .Y(_22478_));
 sky130_as_sc_hs__or2_2 _28990_ (.A(net391),
    .B(\tholin_riscv.regs[2][10] ),
    .Y(_22479_));
 sky130_as_sc_hs__nand2b_2 _28991_ (.B(net391),
    .Y(_22480_),
    .A(\tholin_riscv.regs[3][10] ));
 sky130_as_sc_hs__nand3_2 _28992_ (.A(net357),
    .B(_22479_),
    .C(_22480_),
    .Y(_22481_));
 sky130_as_sc_hs__nand3_2 _28993_ (.A(net234),
    .B(_22478_),
    .C(_22481_),
    .Y(_22482_));
 sky130_as_sc_hs__or2_2 _28994_ (.A(net391),
    .B(\tholin_riscv.regs[6][10] ),
    .Y(_22483_));
 sky130_as_sc_hs__nand2b_2 _28995_ (.B(net391),
    .Y(_22484_),
    .A(\tholin_riscv.regs[7][10] ));
 sky130_as_sc_hs__nand3_2 _28996_ (.A(net357),
    .B(_22483_),
    .C(_22484_),
    .Y(_22485_));
 sky130_as_sc_hs__or2_2 _28997_ (.A(net391),
    .B(\tholin_riscv.regs[4][10] ),
    .Y(_22486_));
 sky130_as_sc_hs__nand2b_2 _28998_ (.B(net401),
    .Y(_22487_),
    .A(\tholin_riscv.regs[5][10] ));
 sky130_as_sc_hs__nand3_2 _28999_ (.A(net217),
    .B(_22486_),
    .C(_22487_),
    .Y(_22488_));
 sky130_as_sc_hs__nand3_2 _29000_ (.A(net345),
    .B(_22485_),
    .C(_22488_),
    .Y(_22489_));
 sky130_as_sc_hs__nand3_2 _29001_ (.A(net241),
    .B(_22482_),
    .C(_22489_),
    .Y(_22490_));
 sky130_as_sc_hs__nand3_2 _29002_ (.A(net338),
    .B(_22468_),
    .C(_22475_),
    .Y(_22491_));
 sky130_as_sc_hs__nand3_2 _29003_ (.A(net245),
    .B(_22490_),
    .C(_22491_),
    .Y(_22492_));
 sky130_as_sc_hs__and2_2 _29004_ (.A(_22461_),
    .B(_22492_),
    .Y(_22493_));
 sky130_as_sc_hs__nor2_2 _29006_ (.A(_22430_),
    .B(_22493_),
    .Y(_22495_));
 sky130_as_sc_hs__or2_2 _29007_ (.A(net392),
    .B(\tholin_riscv.regs[24][9] ),
    .Y(_22496_));
 sky130_as_sc_hs__nand2b_2 _29008_ (.B(net392),
    .Y(_22497_),
    .A(\tholin_riscv.regs[25][9] ));
 sky130_as_sc_hs__nand3_2 _29009_ (.A(net217),
    .B(_22496_),
    .C(_22497_),
    .Y(_22498_));
 sky130_as_sc_hs__or2_2 _29010_ (.A(net392),
    .B(\tholin_riscv.regs[26][9] ),
    .Y(_22499_));
 sky130_as_sc_hs__nand2b_2 _29011_ (.B(net392),
    .Y(_22500_),
    .A(\tholin_riscv.regs[27][9] ));
 sky130_as_sc_hs__nand3_2 _29012_ (.A(net357),
    .B(_22499_),
    .C(_22500_),
    .Y(_22501_));
 sky130_as_sc_hs__nand3_2 _29013_ (.A(net233),
    .B(_22498_),
    .C(_22501_),
    .Y(_22502_));
 sky130_as_sc_hs__or2_2 _29014_ (.A(net403),
    .B(\tholin_riscv.regs[28][9] ),
    .Y(_22503_));
 sky130_as_sc_hs__nand2b_2 _29015_ (.B(net403),
    .Y(_22504_),
    .A(\tholin_riscv.regs[29][9] ));
 sky130_as_sc_hs__nand3_2 _29016_ (.A(net227),
    .B(_22503_),
    .C(_22504_),
    .Y(_22505_));
 sky130_as_sc_hs__or2_2 _29017_ (.A(net403),
    .B(\tholin_riscv.regs[30][9] ),
    .Y(_22506_));
 sky130_as_sc_hs__nand2b_2 _29018_ (.B(net403),
    .Y(_22507_),
    .A(\tholin_riscv.regs[31][9] ));
 sky130_as_sc_hs__nand3_2 _29019_ (.A(net366),
    .B(_22506_),
    .C(_22507_),
    .Y(_22508_));
 sky130_as_sc_hs__nand3_2 _29020_ (.A(net350),
    .B(_22505_),
    .C(_22508_),
    .Y(_22509_));
 sky130_as_sc_hs__or2_2 _29021_ (.A(net392),
    .B(\tholin_riscv.regs[16][9] ),
    .Y(_22510_));
 sky130_as_sc_hs__nand2b_2 _29022_ (.B(net394),
    .Y(_22511_),
    .A(\tholin_riscv.regs[17][9] ));
 sky130_as_sc_hs__nand3_2 _29023_ (.A(net218),
    .B(_22510_),
    .C(_22511_),
    .Y(_22512_));
 sky130_as_sc_hs__or2_2 _29024_ (.A(net392),
    .B(\tholin_riscv.regs[18][9] ),
    .Y(_22513_));
 sky130_as_sc_hs__nand2b_2 _29025_ (.B(net392),
    .Y(_22514_),
    .A(\tholin_riscv.regs[19][9] ));
 sky130_as_sc_hs__nand3_2 _29026_ (.A(net357),
    .B(_22513_),
    .C(_22514_),
    .Y(_22515_));
 sky130_as_sc_hs__nand3_2 _29027_ (.A(net234),
    .B(_22512_),
    .C(_22515_),
    .Y(_22516_));
 sky130_as_sc_hs__or2_2 _29028_ (.A(net393),
    .B(\tholin_riscv.regs[22][9] ),
    .Y(_22517_));
 sky130_as_sc_hs__nand2b_2 _29029_ (.B(net393),
    .Y(_22518_),
    .A(\tholin_riscv.regs[23][9] ));
 sky130_as_sc_hs__nand3_2 _29030_ (.A(net358),
    .B(_22517_),
    .C(_22518_),
    .Y(_22519_));
 sky130_as_sc_hs__or2_2 _29031_ (.A(net403),
    .B(\tholin_riscv.regs[20][9] ),
    .Y(_22520_));
 sky130_as_sc_hs__nand2b_2 _29032_ (.B(net403),
    .Y(_22521_),
    .A(\tholin_riscv.regs[21][9] ));
 sky130_as_sc_hs__nand3_2 _29033_ (.A(net227),
    .B(_22520_),
    .C(_22521_),
    .Y(_22522_));
 sky130_as_sc_hs__nand3_2 _29034_ (.A(net345),
    .B(_22519_),
    .C(_22522_),
    .Y(_22523_));
 sky130_as_sc_hs__nand3_2 _29035_ (.A(net241),
    .B(_22516_),
    .C(_22523_),
    .Y(_22524_));
 sky130_as_sc_hs__nand3_2 _29036_ (.A(net338),
    .B(_22502_),
    .C(_22509_),
    .Y(_22525_));
 sky130_as_sc_hs__nand3_2 _29037_ (.A(net336),
    .B(_22524_),
    .C(_22525_),
    .Y(_22526_));
 sky130_as_sc_hs__or2_2 _29038_ (.A(net403),
    .B(\tholin_riscv.regs[8][9] ),
    .Y(_22527_));
 sky130_as_sc_hs__nand2b_2 _29039_ (.B(net403),
    .Y(_22528_),
    .A(\tholin_riscv.regs[9][9] ));
 sky130_as_sc_hs__nand3_2 _29040_ (.A(net227),
    .B(_22527_),
    .C(_22528_),
    .Y(_22529_));
 sky130_as_sc_hs__or2_2 _29041_ (.A(net403),
    .B(\tholin_riscv.regs[10][9] ),
    .Y(_22530_));
 sky130_as_sc_hs__nand2b_2 _29042_ (.B(net403),
    .Y(_22531_),
    .A(\tholin_riscv.regs[11][9] ));
 sky130_as_sc_hs__nand3_2 _29043_ (.A(net366),
    .B(_22530_),
    .C(_22531_),
    .Y(_22532_));
 sky130_as_sc_hs__nand3_2 _29044_ (.A(net237),
    .B(_22529_),
    .C(_22532_),
    .Y(_22533_));
 sky130_as_sc_hs__or2_2 _29045_ (.A(net402),
    .B(\tholin_riscv.regs[12][9] ),
    .Y(_22534_));
 sky130_as_sc_hs__nand2b_2 _29046_ (.B(net402),
    .Y(_22535_),
    .A(\tholin_riscv.regs[13][9] ));
 sky130_as_sc_hs__nand3_2 _29047_ (.A(net230),
    .B(_22534_),
    .C(_22535_),
    .Y(_22536_));
 sky130_as_sc_hs__or2_2 _29048_ (.A(net404),
    .B(\tholin_riscv.regs[14][9] ),
    .Y(_22537_));
 sky130_as_sc_hs__nand2b_2 _29049_ (.B(net404),
    .Y(_22538_),
    .A(\tholin_riscv.regs[15][9] ));
 sky130_as_sc_hs__nand3_2 _29050_ (.A(net366),
    .B(_22537_),
    .C(_22538_),
    .Y(_22539_));
 sky130_as_sc_hs__nand3_2 _29051_ (.A(net350),
    .B(_22536_),
    .C(_22539_),
    .Y(_22540_));
 sky130_as_sc_hs__or2_2 _29052_ (.A(net401),
    .B(\tholin_riscv.regs[0][9] ),
    .Y(_22541_));
 sky130_as_sc_hs__nand2b_2 _29053_ (.B(net401),
    .Y(_22542_),
    .A(\tholin_riscv.regs[1][9] ));
 sky130_as_sc_hs__nand3_2 _29054_ (.A(net227),
    .B(_22541_),
    .C(_22542_),
    .Y(_22543_));
 sky130_as_sc_hs__or2_2 _29055_ (.A(net401),
    .B(\tholin_riscv.regs[2][9] ),
    .Y(_22544_));
 sky130_as_sc_hs__nand2b_2 _29056_ (.B(net401),
    .Y(_22545_),
    .A(\tholin_riscv.regs[3][9] ));
 sky130_as_sc_hs__nand3_2 _29057_ (.A(net366),
    .B(_22544_),
    .C(_22545_),
    .Y(_22546_));
 sky130_as_sc_hs__nand3_2 _29058_ (.A(net237),
    .B(_22543_),
    .C(_22546_),
    .Y(_22547_));
 sky130_as_sc_hs__or2_2 _29059_ (.A(net401),
    .B(\tholin_riscv.regs[6][9] ),
    .Y(_22548_));
 sky130_as_sc_hs__nand2b_2 _29060_ (.B(net401),
    .Y(_22549_),
    .A(\tholin_riscv.regs[7][9] ));
 sky130_as_sc_hs__nand3_2 _29061_ (.A(net366),
    .B(_22548_),
    .C(_22549_),
    .Y(_22550_));
 sky130_as_sc_hs__or2_2 _29062_ (.A(net401),
    .B(\tholin_riscv.regs[4][9] ),
    .Y(_22551_));
 sky130_as_sc_hs__nand2b_2 _29063_ (.B(net401),
    .Y(_22552_),
    .A(\tholin_riscv.regs[5][9] ));
 sky130_as_sc_hs__nand3_2 _29064_ (.A(net227),
    .B(_22551_),
    .C(_22552_),
    .Y(_22553_));
 sky130_as_sc_hs__nand3_2 _29065_ (.A(net348),
    .B(_22550_),
    .C(_22553_),
    .Y(_22554_));
 sky130_as_sc_hs__nand3_2 _29066_ (.A(net243),
    .B(_22547_),
    .C(_22554_),
    .Y(_22555_));
 sky130_as_sc_hs__nand3_2 _29067_ (.A(net339),
    .B(_22533_),
    .C(_22540_),
    .Y(_22556_));
 sky130_as_sc_hs__nand3_2 _29068_ (.A(net245),
    .B(_22555_),
    .C(_22556_),
    .Y(_22557_));
 sky130_as_sc_hs__and2_2 _29069_ (.A(_22526_),
    .B(_22557_),
    .Y(_22558_));
 sky130_as_sc_hs__or2_2 _29071_ (.A(net405),
    .B(\tholin_riscv.regs[24][8] ),
    .Y(_22560_));
 sky130_as_sc_hs__nand2b_2 _29072_ (.B(net405),
    .Y(_22561_),
    .A(\tholin_riscv.regs[25][8] ));
 sky130_as_sc_hs__nand3_2 _29073_ (.A(net229),
    .B(_22560_),
    .C(_22561_),
    .Y(_22562_));
 sky130_as_sc_hs__or2_2 _29074_ (.A(net405),
    .B(\tholin_riscv.regs[26][8] ),
    .Y(_22563_));
 sky130_as_sc_hs__nand2b_2 _29075_ (.B(net405),
    .Y(_22564_),
    .A(\tholin_riscv.regs[27][8] ));
 sky130_as_sc_hs__nand3_2 _29076_ (.A(net369),
    .B(_22563_),
    .C(_22564_),
    .Y(_22565_));
 sky130_as_sc_hs__nand3_2 _29077_ (.A(net238),
    .B(_22562_),
    .C(_22565_),
    .Y(_22566_));
 sky130_as_sc_hs__or2_2 _29078_ (.A(net405),
    .B(\tholin_riscv.regs[28][8] ),
    .Y(_22567_));
 sky130_as_sc_hs__nand2b_2 _29079_ (.B(net406),
    .Y(_22568_),
    .A(\tholin_riscv.regs[29][8] ));
 sky130_as_sc_hs__nand3_2 _29080_ (.A(net229),
    .B(_22567_),
    .C(_22568_),
    .Y(_22569_));
 sky130_as_sc_hs__or2_2 _29081_ (.A(net406),
    .B(\tholin_riscv.regs[30][8] ),
    .Y(_22570_));
 sky130_as_sc_hs__nand2b_2 _29082_ (.B(net406),
    .Y(_22571_),
    .A(\tholin_riscv.regs[31][8] ));
 sky130_as_sc_hs__nand3_2 _29083_ (.A(net369),
    .B(_22570_),
    .C(_22571_),
    .Y(_22572_));
 sky130_as_sc_hs__nand3_2 _29084_ (.A(net349),
    .B(_22569_),
    .C(_22572_),
    .Y(_22573_));
 sky130_as_sc_hs__or2_2 _29085_ (.A(net407),
    .B(\tholin_riscv.regs[16][8] ),
    .Y(_22574_));
 sky130_as_sc_hs__nand2b_2 _29086_ (.B(net407),
    .Y(_22575_),
    .A(\tholin_riscv.regs[17][8] ));
 sky130_as_sc_hs__nand3_2 _29087_ (.A(net229),
    .B(_22574_),
    .C(_22575_),
    .Y(_22576_));
 sky130_as_sc_hs__or2_2 _29088_ (.A(net407),
    .B(\tholin_riscv.regs[18][8] ),
    .Y(_22577_));
 sky130_as_sc_hs__nand2b_2 _29089_ (.B(net407),
    .Y(_22578_),
    .A(\tholin_riscv.regs[19][8] ));
 sky130_as_sc_hs__nand3_2 _29090_ (.A(net369),
    .B(_22577_),
    .C(_22578_),
    .Y(_22579_));
 sky130_as_sc_hs__nand3_2 _29091_ (.A(net238),
    .B(_22576_),
    .C(_22579_),
    .Y(_22580_));
 sky130_as_sc_hs__or2_2 _29092_ (.A(net407),
    .B(\tholin_riscv.regs[22][8] ),
    .Y(_22581_));
 sky130_as_sc_hs__nand2b_2 _29093_ (.B(net407),
    .Y(_22582_),
    .A(\tholin_riscv.regs[23][8] ));
 sky130_as_sc_hs__nand3_2 _29094_ (.A(net369),
    .B(_22581_),
    .C(_22582_),
    .Y(_22583_));
 sky130_as_sc_hs__or2_2 _29095_ (.A(net407),
    .B(\tholin_riscv.regs[20][8] ),
    .Y(_22584_));
 sky130_as_sc_hs__nand2b_2 _29096_ (.B(net408),
    .Y(_22585_),
    .A(\tholin_riscv.regs[21][8] ));
 sky130_as_sc_hs__nand3_2 _29097_ (.A(net229),
    .B(_22584_),
    .C(_22585_),
    .Y(_22586_));
 sky130_as_sc_hs__nand3_2 _29098_ (.A(net350),
    .B(_22583_),
    .C(_22586_),
    .Y(_22587_));
 sky130_as_sc_hs__nand3_2 _29099_ (.A(net243),
    .B(_22580_),
    .C(_22587_),
    .Y(_22588_));
 sky130_as_sc_hs__nand3_2 _29100_ (.A(net341),
    .B(_22566_),
    .C(_22573_),
    .Y(_22589_));
 sky130_as_sc_hs__nand3_2 _29101_ (.A(\tholin_riscv.Jimm[19] ),
    .B(_22588_),
    .C(_22589_),
    .Y(_22590_));
 sky130_as_sc_hs__or2_2 _29102_ (.A(net402),
    .B(\tholin_riscv.regs[8][8] ),
    .Y(_22591_));
 sky130_as_sc_hs__nand2b_2 _29103_ (.B(net402),
    .Y(_22592_),
    .A(\tholin_riscv.regs[9][8] ));
 sky130_as_sc_hs__nand3_2 _29104_ (.A(net230),
    .B(_22591_),
    .C(_22592_),
    .Y(_22593_));
 sky130_as_sc_hs__or2_2 _29105_ (.A(net402),
    .B(\tholin_riscv.regs[10][8] ),
    .Y(_22594_));
 sky130_as_sc_hs__nand2b_2 _29106_ (.B(net402),
    .Y(_22595_),
    .A(\tholin_riscv.regs[11][8] ));
 sky130_as_sc_hs__nand3_2 _29107_ (.A(net370),
    .B(_22594_),
    .C(_22595_),
    .Y(_22596_));
 sky130_as_sc_hs__nand3_2 _29108_ (.A(net238),
    .B(_22593_),
    .C(_22596_),
    .Y(_22597_));
 sky130_as_sc_hs__or2_2 _29109_ (.A(net405),
    .B(\tholin_riscv.regs[12][8] ),
    .Y(_22598_));
 sky130_as_sc_hs__nand2b_2 _29110_ (.B(net405),
    .Y(_22599_),
    .A(\tholin_riscv.regs[13][8] ));
 sky130_as_sc_hs__nand3_2 _29111_ (.A(net229),
    .B(_22598_),
    .C(_22599_),
    .Y(_22600_));
 sky130_as_sc_hs__or2_2 _29112_ (.A(net405),
    .B(\tholin_riscv.regs[14][8] ),
    .Y(_22601_));
 sky130_as_sc_hs__nand2b_2 _29113_ (.B(net405),
    .Y(_22602_),
    .A(\tholin_riscv.regs[15][8] ));
 sky130_as_sc_hs__nand3_2 _29114_ (.A(net369),
    .B(_22601_),
    .C(_22602_),
    .Y(_22603_));
 sky130_as_sc_hs__nand3_2 _29115_ (.A(net350),
    .B(_22600_),
    .C(_22603_),
    .Y(_22604_));
 sky130_as_sc_hs__or2_2 _29116_ (.A(net408),
    .B(\tholin_riscv.regs[0][8] ),
    .Y(_22605_));
 sky130_as_sc_hs__nand2b_2 _29117_ (.B(net404),
    .Y(_22606_),
    .A(\tholin_riscv.regs[1][8] ));
 sky130_as_sc_hs__nand3_2 _29118_ (.A(net227),
    .B(_22605_),
    .C(_22606_),
    .Y(_22607_));
 sky130_as_sc_hs__or2_2 _29119_ (.A(net401),
    .B(\tholin_riscv.regs[2][8] ),
    .Y(_22608_));
 sky130_as_sc_hs__nand2b_2 _29120_ (.B(net401),
    .Y(_22609_),
    .A(\tholin_riscv.regs[3][8] ));
 sky130_as_sc_hs__nand3_2 _29121_ (.A(net366),
    .B(_22608_),
    .C(_22609_),
    .Y(_22610_));
 sky130_as_sc_hs__nand3_2 _29122_ (.A(net238),
    .B(_22607_),
    .C(_22610_),
    .Y(_22611_));
 sky130_as_sc_hs__or2_2 _29123_ (.A(net404),
    .B(\tholin_riscv.regs[6][8] ),
    .Y(_22612_));
 sky130_as_sc_hs__nand2b_2 _29124_ (.B(net404),
    .Y(_22613_),
    .A(\tholin_riscv.regs[7][8] ));
 sky130_as_sc_hs__nand3_2 _29125_ (.A(net366),
    .B(_22612_),
    .C(_22613_),
    .Y(_22614_));
 sky130_as_sc_hs__or2_2 _29126_ (.A(net407),
    .B(\tholin_riscv.regs[4][8] ),
    .Y(_22615_));
 sky130_as_sc_hs__nand2b_2 _29127_ (.B(net407),
    .Y(_22616_),
    .A(\tholin_riscv.regs[5][8] ));
 sky130_as_sc_hs__nand3_2 _29128_ (.A(net229),
    .B(_22615_),
    .C(_22616_),
    .Y(_22617_));
 sky130_as_sc_hs__nand3_2 _29129_ (.A(net350),
    .B(_22614_),
    .C(_22617_),
    .Y(_22618_));
 sky130_as_sc_hs__nand3_2 _29130_ (.A(net243),
    .B(_22611_),
    .C(_22618_),
    .Y(_22619_));
 sky130_as_sc_hs__nand3_2 _29131_ (.A(net339),
    .B(_22597_),
    .C(_22604_),
    .Y(_22620_));
 sky130_as_sc_hs__nand3_2 _29132_ (.A(net245),
    .B(_22619_),
    .C(_22620_),
    .Y(_22621_));
 sky130_as_sc_hs__and2_2 _29133_ (.A(_22590_),
    .B(_22621_),
    .Y(_22622_));
 sky130_as_sc_hs__nor2_2 _29134_ (.A(_22558_),
    .B(_22622_),
    .Y(_22623_));
 sky130_as_sc_hs__and2_2 _29135_ (.A(_22495_),
    .B(_22623_),
    .Y(_22624_));
 sky130_as_sc_hs__or2_2 _29136_ (.A(net383),
    .B(\tholin_riscv.regs[24][14] ),
    .Y(_22625_));
 sky130_as_sc_hs__or2_2 _29137_ (.A(net201),
    .B(\tholin_riscv.regs[25][14] ),
    .Y(_22626_));
 sky130_as_sc_hs__nand3_2 _29138_ (.A(net211),
    .B(_22625_),
    .C(_22626_),
    .Y(_22627_));
 sky130_as_sc_hs__or2_2 _29139_ (.A(net383),
    .B(\tholin_riscv.regs[26][14] ),
    .Y(_22628_));
 sky130_as_sc_hs__or2_2 _29140_ (.A(net201),
    .B(\tholin_riscv.regs[27][14] ),
    .Y(_22629_));
 sky130_as_sc_hs__nand3_2 _29141_ (.A(net351),
    .B(_22628_),
    .C(_22629_),
    .Y(_22630_));
 sky130_as_sc_hs__nand3_2 _29142_ (.A(net232),
    .B(_22627_),
    .C(_22630_),
    .Y(_22631_));
 sky130_as_sc_hs__or2_2 _29143_ (.A(net372),
    .B(\tholin_riscv.regs[28][14] ),
    .Y(_22632_));
 sky130_as_sc_hs__or2_2 _29144_ (.A(net201),
    .B(\tholin_riscv.regs[29][14] ),
    .Y(_22633_));
 sky130_as_sc_hs__nand3_2 _29145_ (.A(net211),
    .B(_22632_),
    .C(_22633_),
    .Y(_22634_));
 sky130_as_sc_hs__or2_2 _29146_ (.A(net372),
    .B(\tholin_riscv.regs[30][14] ),
    .Y(_22635_));
 sky130_as_sc_hs__or2_2 _29147_ (.A(net201),
    .B(\tholin_riscv.regs[31][14] ),
    .Y(_22636_));
 sky130_as_sc_hs__nand3_2 _29148_ (.A(net351),
    .B(_22635_),
    .C(_22636_),
    .Y(_22637_));
 sky130_as_sc_hs__nand3_2 _29149_ (.A(net343),
    .B(_22634_),
    .C(_22637_),
    .Y(_22638_));
 sky130_as_sc_hs__or2_2 _29150_ (.A(net372),
    .B(\tholin_riscv.regs[16][14] ),
    .Y(_22639_));
 sky130_as_sc_hs__or2_2 _29151_ (.A(net201),
    .B(\tholin_riscv.regs[17][14] ),
    .Y(_22640_));
 sky130_as_sc_hs__nand3_2 _29152_ (.A(net211),
    .B(_22639_),
    .C(_22640_),
    .Y(_22641_));
 sky130_as_sc_hs__or2_2 _29153_ (.A(net372),
    .B(\tholin_riscv.regs[18][14] ),
    .Y(_22642_));
 sky130_as_sc_hs__or2_2 _29154_ (.A(net201),
    .B(\tholin_riscv.regs[19][14] ),
    .Y(_22643_));
 sky130_as_sc_hs__nand3_2 _29155_ (.A(net351),
    .B(_22642_),
    .C(_22643_),
    .Y(_22644_));
 sky130_as_sc_hs__nand3_2 _29156_ (.A(net232),
    .B(_22641_),
    .C(_22644_),
    .Y(_22645_));
 sky130_as_sc_hs__or2_2 _29157_ (.A(net383),
    .B(\tholin_riscv.regs[22][14] ),
    .Y(_22646_));
 sky130_as_sc_hs__or2_2 _29158_ (.A(net201),
    .B(\tholin_riscv.regs[23][14] ),
    .Y(_22647_));
 sky130_as_sc_hs__nand3_2 _29159_ (.A(net351),
    .B(_22646_),
    .C(_22647_),
    .Y(_22648_));
 sky130_as_sc_hs__or2_2 _29160_ (.A(net383),
    .B(\tholin_riscv.regs[20][14] ),
    .Y(_22649_));
 sky130_as_sc_hs__or2_2 _29161_ (.A(net201),
    .B(\tholin_riscv.regs[21][14] ),
    .Y(_22650_));
 sky130_as_sc_hs__nand3_2 _29162_ (.A(net211),
    .B(_22649_),
    .C(_22650_),
    .Y(_22651_));
 sky130_as_sc_hs__nand3_2 _29163_ (.A(net343),
    .B(_22648_),
    .C(_22651_),
    .Y(_22652_));
 sky130_as_sc_hs__nand3_2 _29164_ (.A(net240),
    .B(_22645_),
    .C(_22652_),
    .Y(_22653_));
 sky130_as_sc_hs__nand3_2 _29165_ (.A(net337),
    .B(_22631_),
    .C(_22638_),
    .Y(_22654_));
 sky130_as_sc_hs__nand3_2 _29166_ (.A(net336),
    .B(_22653_),
    .C(_22654_),
    .Y(_22655_));
 sky130_as_sc_hs__or2_2 _29167_ (.A(net384),
    .B(\tholin_riscv.regs[8][14] ),
    .Y(_22656_));
 sky130_as_sc_hs__or2_2 _29168_ (.A(net202),
    .B(\tholin_riscv.regs[9][14] ),
    .Y(_22657_));
 sky130_as_sc_hs__nand3_2 _29169_ (.A(net211),
    .B(_22656_),
    .C(_22657_),
    .Y(_22658_));
 sky130_as_sc_hs__or2_2 _29170_ (.A(net383),
    .B(\tholin_riscv.regs[10][14] ),
    .Y(_22659_));
 sky130_as_sc_hs__or2_2 _29171_ (.A(net202),
    .B(\tholin_riscv.regs[11][14] ),
    .Y(_22660_));
 sky130_as_sc_hs__nand3_2 _29172_ (.A(net351),
    .B(_22659_),
    .C(_22660_),
    .Y(_22661_));
 sky130_as_sc_hs__nand3_2 _29173_ (.A(net232),
    .B(_22658_),
    .C(_22661_),
    .Y(_22662_));
 sky130_as_sc_hs__or2_2 _29174_ (.A(net383),
    .B(\tholin_riscv.regs[12][14] ),
    .Y(_22663_));
 sky130_as_sc_hs__or2_2 _29175_ (.A(net202),
    .B(\tholin_riscv.regs[13][14] ),
    .Y(_22664_));
 sky130_as_sc_hs__nand3_2 _29176_ (.A(net211),
    .B(_22663_),
    .C(_22664_),
    .Y(_22665_));
 sky130_as_sc_hs__or2_2 _29177_ (.A(net383),
    .B(\tholin_riscv.regs[14][14] ),
    .Y(_22666_));
 sky130_as_sc_hs__or2_2 _29178_ (.A(net202),
    .B(\tholin_riscv.regs[15][14] ),
    .Y(_22667_));
 sky130_as_sc_hs__nand3_2 _29179_ (.A(net351),
    .B(_22666_),
    .C(_22667_),
    .Y(_22668_));
 sky130_as_sc_hs__nand3_2 _29180_ (.A(net343),
    .B(_22665_),
    .C(_22668_),
    .Y(_22669_));
 sky130_as_sc_hs__or2_2 _29181_ (.A(net372),
    .B(\tholin_riscv.regs[0][14] ),
    .Y(_22670_));
 sky130_as_sc_hs__or2_2 _29182_ (.A(net202),
    .B(\tholin_riscv.regs[1][14] ),
    .Y(_22671_));
 sky130_as_sc_hs__nand3_2 _29183_ (.A(net211),
    .B(_22670_),
    .C(_22671_),
    .Y(_22672_));
 sky130_as_sc_hs__or2_2 _29184_ (.A(net372),
    .B(\tholin_riscv.regs[2][14] ),
    .Y(_22673_));
 sky130_as_sc_hs__or2_2 _29185_ (.A(net202),
    .B(\tholin_riscv.regs[3][14] ),
    .Y(_22674_));
 sky130_as_sc_hs__nand3_2 _29186_ (.A(net351),
    .B(_22673_),
    .C(_22674_),
    .Y(_22675_));
 sky130_as_sc_hs__nand3_2 _29187_ (.A(net232),
    .B(_22672_),
    .C(_22675_),
    .Y(_22676_));
 sky130_as_sc_hs__or2_2 _29188_ (.A(net372),
    .B(\tholin_riscv.regs[6][14] ),
    .Y(_22677_));
 sky130_as_sc_hs__or2_2 _29189_ (.A(net202),
    .B(\tholin_riscv.regs[7][14] ),
    .Y(_22678_));
 sky130_as_sc_hs__nand3_2 _29190_ (.A(net351),
    .B(_22677_),
    .C(_22678_),
    .Y(_22679_));
 sky130_as_sc_hs__or2_2 _29191_ (.A(net372),
    .B(\tholin_riscv.regs[4][14] ),
    .Y(_22680_));
 sky130_as_sc_hs__or2_2 _29192_ (.A(net202),
    .B(\tholin_riscv.regs[5][14] ),
    .Y(_22681_));
 sky130_as_sc_hs__nand3_2 _29193_ (.A(net211),
    .B(_22680_),
    .C(_22681_),
    .Y(_22682_));
 sky130_as_sc_hs__nand3_2 _29194_ (.A(net343),
    .B(_22679_),
    .C(_22682_),
    .Y(_22683_));
 sky130_as_sc_hs__nand3_2 _29195_ (.A(net240),
    .B(_22676_),
    .C(_22683_),
    .Y(_22684_));
 sky130_as_sc_hs__nand3_2 _29196_ (.A(net337),
    .B(_22662_),
    .C(_22669_),
    .Y(_22685_));
 sky130_as_sc_hs__nand3_2 _29197_ (.A(net246),
    .B(_22684_),
    .C(_22685_),
    .Y(_22686_));
 sky130_as_sc_hs__and2_2 _29198_ (.A(_22655_),
    .B(_22686_),
    .Y(_22687_));
 sky130_as_sc_hs__or2_2 _29199_ (.A(net383),
    .B(\tholin_riscv.regs[24][15] ),
    .Y(_22688_));
 sky130_as_sc_hs__or2_2 _29200_ (.A(net201),
    .B(\tholin_riscv.regs[25][15] ),
    .Y(_22689_));
 sky130_as_sc_hs__nand3_2 _29201_ (.A(net211),
    .B(_22688_),
    .C(_22689_),
    .Y(_22690_));
 sky130_as_sc_hs__or2_2 _29202_ (.A(net383),
    .B(\tholin_riscv.regs[26][15] ),
    .Y(_22691_));
 sky130_as_sc_hs__or2_2 _29203_ (.A(net201),
    .B(\tholin_riscv.regs[27][15] ),
    .Y(_22692_));
 sky130_as_sc_hs__nand3_2 _29204_ (.A(net351),
    .B(_22691_),
    .C(_22692_),
    .Y(_22693_));
 sky130_as_sc_hs__nand3_2 _29205_ (.A(net232),
    .B(_22690_),
    .C(_22693_),
    .Y(_22694_));
 sky130_as_sc_hs__or2_2 _29206_ (.A(net383),
    .B(\tholin_riscv.regs[28][15] ),
    .Y(_22695_));
 sky130_as_sc_hs__or2_2 _29207_ (.A(net201),
    .B(\tholin_riscv.regs[29][15] ),
    .Y(_22696_));
 sky130_as_sc_hs__nand3_2 _29208_ (.A(net211),
    .B(_22695_),
    .C(_22696_),
    .Y(_22697_));
 sky130_as_sc_hs__or2_2 _29209_ (.A(net383),
    .B(\tholin_riscv.regs[30][15] ),
    .Y(_22698_));
 sky130_as_sc_hs__or2_2 _29210_ (.A(net203),
    .B(\tholin_riscv.regs[31][15] ),
    .Y(_22699_));
 sky130_as_sc_hs__nand3_2 _29211_ (.A(net355),
    .B(_22698_),
    .C(_22699_),
    .Y(_22700_));
 sky130_as_sc_hs__nand3_2 _29212_ (.A(net344),
    .B(_22697_),
    .C(_22700_),
    .Y(_22701_));
 sky130_as_sc_hs__or2_2 _29213_ (.A(net384),
    .B(\tholin_riscv.regs[16][15] ),
    .Y(_22702_));
 sky130_as_sc_hs__or2_2 _29214_ (.A(net203),
    .B(\tholin_riscv.regs[17][15] ),
    .Y(_22703_));
 sky130_as_sc_hs__nand3_2 _29215_ (.A(net219),
    .B(_22702_),
    .C(_22703_),
    .Y(_22704_));
 sky130_as_sc_hs__or2_2 _29216_ (.A(net383),
    .B(\tholin_riscv.regs[18][15] ),
    .Y(_22705_));
 sky130_as_sc_hs__or2_2 _29217_ (.A(net203),
    .B(\tholin_riscv.regs[19][15] ),
    .Y(_22706_));
 sky130_as_sc_hs__nand3_2 _29218_ (.A(net355),
    .B(_22705_),
    .C(_22706_),
    .Y(_22707_));
 sky130_as_sc_hs__nand3_2 _29219_ (.A(net232),
    .B(_22704_),
    .C(_22707_),
    .Y(_22708_));
 sky130_as_sc_hs__or2_2 _29220_ (.A(net384),
    .B(\tholin_riscv.regs[22][15] ),
    .Y(_22709_));
 sky130_as_sc_hs__or2_2 _29221_ (.A(net203),
    .B(\tholin_riscv.regs[23][15] ),
    .Y(_22710_));
 sky130_as_sc_hs__nand3_2 _29222_ (.A(net355),
    .B(_22709_),
    .C(_22710_),
    .Y(_22711_));
 sky130_as_sc_hs__or2_2 _29223_ (.A(net383),
    .B(\tholin_riscv.regs[20][15] ),
    .Y(_22712_));
 sky130_as_sc_hs__or2_2 _29224_ (.A(net203),
    .B(\tholin_riscv.regs[21][15] ),
    .Y(_22713_));
 sky130_as_sc_hs__nand3_2 _29225_ (.A(net211),
    .B(_22712_),
    .C(_22713_),
    .Y(_22714_));
 sky130_as_sc_hs__nand3_2 _29226_ (.A(net344),
    .B(_22711_),
    .C(_22714_),
    .Y(_22715_));
 sky130_as_sc_hs__nand3_2 _29227_ (.A(net240),
    .B(_22708_),
    .C(_22715_),
    .Y(_22716_));
 sky130_as_sc_hs__nand3_2 _29228_ (.A(net338),
    .B(_22694_),
    .C(_22701_),
    .Y(_22717_));
 sky130_as_sc_hs__nand3_2 _29229_ (.A(net336),
    .B(_22716_),
    .C(_22717_),
    .Y(_22718_));
 sky130_as_sc_hs__or2_2 _29230_ (.A(net384),
    .B(\tholin_riscv.regs[8][15] ),
    .Y(_22719_));
 sky130_as_sc_hs__or2_2 _29231_ (.A(net203),
    .B(\tholin_riscv.regs[9][15] ),
    .Y(_22720_));
 sky130_as_sc_hs__nand3_2 _29232_ (.A(net215),
    .B(_22719_),
    .C(_22720_),
    .Y(_22721_));
 sky130_as_sc_hs__or2_2 _29233_ (.A(net384),
    .B(\tholin_riscv.regs[10][15] ),
    .Y(_22722_));
 sky130_as_sc_hs__or2_2 _29234_ (.A(net210),
    .B(\tholin_riscv.regs[11][15] ),
    .Y(_22723_));
 sky130_as_sc_hs__nand3_2 _29235_ (.A(net355),
    .B(_22722_),
    .C(_22723_),
    .Y(_22724_));
 sky130_as_sc_hs__nand3_2 _29236_ (.A(net233),
    .B(_22721_),
    .C(_22724_),
    .Y(_22725_));
 sky130_as_sc_hs__or2_2 _29237_ (.A(net384),
    .B(\tholin_riscv.regs[12][15] ),
    .Y(_22726_));
 sky130_as_sc_hs__or2_2 _29238_ (.A(net203),
    .B(\tholin_riscv.regs[13][15] ),
    .Y(_22727_));
 sky130_as_sc_hs__nand3_2 _29239_ (.A(net215),
    .B(_22726_),
    .C(_22727_),
    .Y(_22728_));
 sky130_as_sc_hs__or2_2 _29240_ (.A(net384),
    .B(\tholin_riscv.regs[14][15] ),
    .Y(_22729_));
 sky130_as_sc_hs__or2_2 _29241_ (.A(net203),
    .B(\tholin_riscv.regs[15][15] ),
    .Y(_22730_));
 sky130_as_sc_hs__nand3_2 _29242_ (.A(net355),
    .B(_22729_),
    .C(_22730_),
    .Y(_22731_));
 sky130_as_sc_hs__nand3_2 _29243_ (.A(net344),
    .B(_22728_),
    .C(_22731_),
    .Y(_22732_));
 sky130_as_sc_hs__or2_2 _29244_ (.A(net384),
    .B(\tholin_riscv.regs[0][15] ),
    .Y(_22733_));
 sky130_as_sc_hs__or2_2 _29245_ (.A(net201),
    .B(\tholin_riscv.regs[1][15] ),
    .Y(_22734_));
 sky130_as_sc_hs__nand3_2 _29246_ (.A(net211),
    .B(_22733_),
    .C(_22734_),
    .Y(_22735_));
 sky130_as_sc_hs__or2_2 _29247_ (.A(net383),
    .B(\tholin_riscv.regs[2][15] ),
    .Y(_22736_));
 sky130_as_sc_hs__or2_2 _29248_ (.A(net210),
    .B(\tholin_riscv.regs[3][15] ),
    .Y(_22737_));
 sky130_as_sc_hs__nand3_2 _29249_ (.A(net355),
    .B(_22736_),
    .C(_22737_),
    .Y(_22738_));
 sky130_as_sc_hs__nand3_2 _29250_ (.A(net232),
    .B(_22735_),
    .C(_22738_),
    .Y(_22739_));
 sky130_as_sc_hs__or2_2 _29251_ (.A(net383),
    .B(\tholin_riscv.regs[6][15] ),
    .Y(_22740_));
 sky130_as_sc_hs__or2_2 _29252_ (.A(net203),
    .B(\tholin_riscv.regs[7][15] ),
    .Y(_22741_));
 sky130_as_sc_hs__nand3_2 _29253_ (.A(net355),
    .B(_22740_),
    .C(_22741_),
    .Y(_22742_));
 sky130_as_sc_hs__or2_2 _29254_ (.A(net383),
    .B(\tholin_riscv.regs[4][15] ),
    .Y(_22743_));
 sky130_as_sc_hs__or2_2 _29255_ (.A(net203),
    .B(\tholin_riscv.regs[5][15] ),
    .Y(_22744_));
 sky130_as_sc_hs__nand3_2 _29256_ (.A(net219),
    .B(_22743_),
    .C(_22744_),
    .Y(_22745_));
 sky130_as_sc_hs__nand3_2 _29257_ (.A(net344),
    .B(_22742_),
    .C(_22745_),
    .Y(_22746_));
 sky130_as_sc_hs__nand3_2 _29258_ (.A(net240),
    .B(_22739_),
    .C(_22746_),
    .Y(_22747_));
 sky130_as_sc_hs__nand3_2 _29259_ (.A(net338),
    .B(_22725_),
    .C(_22732_),
    .Y(_22748_));
 sky130_as_sc_hs__nand3_2 _29260_ (.A(net246),
    .B(_22747_),
    .C(_22748_),
    .Y(_22749_));
 sky130_as_sc_hs__inv_2 _29262_ (.Y(_22751_),
    .A(_22750_));
 sky130_as_sc_hs__nor2b_2 _29263_ (.A(_22687_),
    .Y(_22752_),
    .B(_22750_));
 sky130_as_sc_hs__or2_2 _29264_ (.A(net388),
    .B(\tholin_riscv.regs[24][13] ),
    .Y(_22753_));
 sky130_as_sc_hs__or2_2 _29265_ (.A(net208),
    .B(\tholin_riscv.regs[25][13] ),
    .Y(_22754_));
 sky130_as_sc_hs__nand3_2 _29266_ (.A(net215),
    .B(_22753_),
    .C(_22754_),
    .Y(_22755_));
 sky130_as_sc_hs__or2_2 _29267_ (.A(net388),
    .B(\tholin_riscv.regs[26][13] ),
    .Y(_22756_));
 sky130_as_sc_hs__or2_2 _29268_ (.A(net208),
    .B(\tholin_riscv.regs[27][13] ),
    .Y(_22757_));
 sky130_as_sc_hs__nand3_2 _29269_ (.A(net355),
    .B(_22756_),
    .C(_22757_),
    .Y(_22758_));
 sky130_as_sc_hs__nand3_2 _29270_ (.A(net233),
    .B(_22755_),
    .C(_22758_),
    .Y(_22759_));
 sky130_as_sc_hs__or2_2 _29271_ (.A(net388),
    .B(\tholin_riscv.regs[28][13] ),
    .Y(_22760_));
 sky130_as_sc_hs__or2_2 _29272_ (.A(net208),
    .B(\tholin_riscv.regs[29][13] ),
    .Y(_22761_));
 sky130_as_sc_hs__nand3_2 _29273_ (.A(net216),
    .B(_22760_),
    .C(_22761_),
    .Y(_22762_));
 sky130_as_sc_hs__or2_2 _29274_ (.A(net388),
    .B(\tholin_riscv.regs[30][13] ),
    .Y(_22763_));
 sky130_as_sc_hs__or2_2 _29275_ (.A(net208),
    .B(\tholin_riscv.regs[31][13] ),
    .Y(_22764_));
 sky130_as_sc_hs__nand3_2 _29276_ (.A(net356),
    .B(_22763_),
    .C(_22764_),
    .Y(_22765_));
 sky130_as_sc_hs__nand3_2 _29277_ (.A(net344),
    .B(_22762_),
    .C(_22765_),
    .Y(_22766_));
 sky130_as_sc_hs__or2_2 _29278_ (.A(net388),
    .B(\tholin_riscv.regs[16][13] ),
    .Y(_22767_));
 sky130_as_sc_hs__or2_2 _29279_ (.A(net208),
    .B(\tholin_riscv.regs[17][13] ),
    .Y(_22768_));
 sky130_as_sc_hs__nand3_2 _29280_ (.A(net215),
    .B(_22767_),
    .C(_22768_),
    .Y(_22769_));
 sky130_as_sc_hs__or2_2 _29281_ (.A(net388),
    .B(\tholin_riscv.regs[18][13] ),
    .Y(_22770_));
 sky130_as_sc_hs__or2_2 _29282_ (.A(net208),
    .B(\tholin_riscv.regs[19][13] ),
    .Y(_22771_));
 sky130_as_sc_hs__nand3_2 _29283_ (.A(net355),
    .B(_22770_),
    .C(_22771_),
    .Y(_22772_));
 sky130_as_sc_hs__nand3_2 _29284_ (.A(net233),
    .B(_22769_),
    .C(_22772_),
    .Y(_22773_));
 sky130_as_sc_hs__or2_2 _29285_ (.A(net384),
    .B(\tholin_riscv.regs[22][13] ),
    .Y(_22774_));
 sky130_as_sc_hs__or2_2 _29286_ (.A(net208),
    .B(\tholin_riscv.regs[23][13] ),
    .Y(_22775_));
 sky130_as_sc_hs__nand3_2 _29287_ (.A(net355),
    .B(_22774_),
    .C(_22775_),
    .Y(_22776_));
 sky130_as_sc_hs__or2_2 _29288_ (.A(net388),
    .B(\tholin_riscv.regs[20][13] ),
    .Y(_22777_));
 sky130_as_sc_hs__or2_2 _29289_ (.A(net208),
    .B(\tholin_riscv.regs[21][13] ),
    .Y(_22778_));
 sky130_as_sc_hs__nand3_2 _29290_ (.A(net215),
    .B(_22777_),
    .C(_22778_),
    .Y(_22779_));
 sky130_as_sc_hs__nand3_2 _29291_ (.A(net344),
    .B(_22776_),
    .C(_22779_),
    .Y(_22780_));
 sky130_as_sc_hs__nand3_2 _29292_ (.A(net241),
    .B(_22773_),
    .C(_22780_),
    .Y(_22781_));
 sky130_as_sc_hs__nand3_2 _29293_ (.A(net338),
    .B(_22759_),
    .C(_22766_),
    .Y(_22782_));
 sky130_as_sc_hs__nand3_2 _29294_ (.A(net336),
    .B(_22781_),
    .C(_22782_),
    .Y(_22783_));
 sky130_as_sc_hs__or2_2 _29295_ (.A(net389),
    .B(\tholin_riscv.regs[8][13] ),
    .Y(_22784_));
 sky130_as_sc_hs__or2_2 _29296_ (.A(net207),
    .B(\tholin_riscv.regs[9][13] ),
    .Y(_22785_));
 sky130_as_sc_hs__nand3_2 _29297_ (.A(net215),
    .B(_22784_),
    .C(_22785_),
    .Y(_22786_));
 sky130_as_sc_hs__or2_2 _29298_ (.A(net389),
    .B(\tholin_riscv.regs[10][13] ),
    .Y(_22787_));
 sky130_as_sc_hs__or2_2 _29299_ (.A(net207),
    .B(\tholin_riscv.regs[11][13] ),
    .Y(_22788_));
 sky130_as_sc_hs__nand3_2 _29300_ (.A(net356),
    .B(_22787_),
    .C(_22788_),
    .Y(_22789_));
 sky130_as_sc_hs__nand3_2 _29301_ (.A(net233),
    .B(_22786_),
    .C(_22789_),
    .Y(_22790_));
 sky130_as_sc_hs__or2_2 _29302_ (.A(net389),
    .B(\tholin_riscv.regs[12][13] ),
    .Y(_22791_));
 sky130_as_sc_hs__or2_2 _29303_ (.A(net207),
    .B(\tholin_riscv.regs[13][13] ),
    .Y(_22792_));
 sky130_as_sc_hs__nand3_2 _29304_ (.A(net215),
    .B(_22791_),
    .C(_22792_),
    .Y(_22793_));
 sky130_as_sc_hs__or2_2 _29305_ (.A(net394),
    .B(\tholin_riscv.regs[14][13] ),
    .Y(_22794_));
 sky130_as_sc_hs__or2_2 _29306_ (.A(net207),
    .B(\tholin_riscv.regs[15][13] ),
    .Y(_22795_));
 sky130_as_sc_hs__nand3_2 _29307_ (.A(net356),
    .B(_22794_),
    .C(_22795_),
    .Y(_22796_));
 sky130_as_sc_hs__nand3_2 _29308_ (.A(net344),
    .B(_22793_),
    .C(_22796_),
    .Y(_22797_));
 sky130_as_sc_hs__or2_2 _29309_ (.A(net389),
    .B(\tholin_riscv.regs[0][13] ),
    .Y(_22798_));
 sky130_as_sc_hs__or2_2 _29310_ (.A(net207),
    .B(\tholin_riscv.regs[1][13] ),
    .Y(_22799_));
 sky130_as_sc_hs__nand3_2 _29311_ (.A(net215),
    .B(_22798_),
    .C(_22799_),
    .Y(_22800_));
 sky130_as_sc_hs__or2_2 _29312_ (.A(net389),
    .B(\tholin_riscv.regs[2][13] ),
    .Y(_22801_));
 sky130_as_sc_hs__or2_2 _29313_ (.A(net207),
    .B(\tholin_riscv.regs[3][13] ),
    .Y(_22802_));
 sky130_as_sc_hs__nand3_2 _29314_ (.A(net356),
    .B(_22801_),
    .C(_22802_),
    .Y(_22803_));
 sky130_as_sc_hs__nand3_2 _29315_ (.A(net233),
    .B(_22800_),
    .C(_22803_),
    .Y(_22804_));
 sky130_as_sc_hs__or2_2 _29316_ (.A(net389),
    .B(\tholin_riscv.regs[6][13] ),
    .Y(_22805_));
 sky130_as_sc_hs__or2_2 _29317_ (.A(net208),
    .B(\tholin_riscv.regs[7][13] ),
    .Y(_22806_));
 sky130_as_sc_hs__nand3_2 _29318_ (.A(net356),
    .B(_22805_),
    .C(_22806_),
    .Y(_22807_));
 sky130_as_sc_hs__or2_2 _29319_ (.A(net389),
    .B(\tholin_riscv.regs[4][13] ),
    .Y(_22808_));
 sky130_as_sc_hs__or2_2 _29320_ (.A(net207),
    .B(\tholin_riscv.regs[5][13] ),
    .Y(_22809_));
 sky130_as_sc_hs__nand3_2 _29321_ (.A(net215),
    .B(_22808_),
    .C(_22809_),
    .Y(_22810_));
 sky130_as_sc_hs__nand3_2 _29322_ (.A(net344),
    .B(_22807_),
    .C(_22810_),
    .Y(_22811_));
 sky130_as_sc_hs__nand3_2 _29323_ (.A(net241),
    .B(_22804_),
    .C(_22811_),
    .Y(_22812_));
 sky130_as_sc_hs__nand3_2 _29324_ (.A(net338),
    .B(_22790_),
    .C(_22797_),
    .Y(_22813_));
 sky130_as_sc_hs__nand3_2 _29325_ (.A(net245),
    .B(_22812_),
    .C(_22813_),
    .Y(_22814_));
 sky130_as_sc_hs__inv_2 _29327_ (.Y(_22816_),
    .A(_22815_));
 sky130_as_sc_hs__or2_2 _29328_ (.A(net389),
    .B(\tholin_riscv.regs[24][12] ),
    .Y(_22817_));
 sky130_as_sc_hs__or2_2 _29329_ (.A(net207),
    .B(\tholin_riscv.regs[25][12] ),
    .Y(_22818_));
 sky130_as_sc_hs__nand3_2 _29330_ (.A(net215),
    .B(_22817_),
    .C(_22818_),
    .Y(_22819_));
 sky130_as_sc_hs__or2_2 _29331_ (.A(net389),
    .B(\tholin_riscv.regs[26][12] ),
    .Y(_22820_));
 sky130_as_sc_hs__or2_2 _29332_ (.A(net207),
    .B(\tholin_riscv.regs[27][12] ),
    .Y(_22821_));
 sky130_as_sc_hs__nand3_2 _29333_ (.A(net356),
    .B(_22820_),
    .C(_22821_),
    .Y(_22822_));
 sky130_as_sc_hs__nand3_2 _29334_ (.A(net233),
    .B(_22819_),
    .C(_22822_),
    .Y(_22823_));
 sky130_as_sc_hs__or2_2 _29335_ (.A(net389),
    .B(\tholin_riscv.regs[28][12] ),
    .Y(_22824_));
 sky130_as_sc_hs__or2_2 _29336_ (.A(net207),
    .B(\tholin_riscv.regs[29][12] ),
    .Y(_22825_));
 sky130_as_sc_hs__nand3_2 _29337_ (.A(net216),
    .B(_22824_),
    .C(_22825_),
    .Y(_22826_));
 sky130_as_sc_hs__or2_2 _29338_ (.A(net389),
    .B(\tholin_riscv.regs[30][12] ),
    .Y(_22827_));
 sky130_as_sc_hs__or2_2 _29339_ (.A(net207),
    .B(\tholin_riscv.regs[31][12] ),
    .Y(_22828_));
 sky130_as_sc_hs__nand3_2 _29340_ (.A(net356),
    .B(_22827_),
    .C(_22828_),
    .Y(_22829_));
 sky130_as_sc_hs__nand3_2 _29341_ (.A(net344),
    .B(_22826_),
    .C(_22829_),
    .Y(_22830_));
 sky130_as_sc_hs__or2_2 _29342_ (.A(net389),
    .B(\tholin_riscv.regs[16][12] ),
    .Y(_22831_));
 sky130_as_sc_hs__or2_2 _29343_ (.A(net207),
    .B(\tholin_riscv.regs[17][12] ),
    .Y(_22832_));
 sky130_as_sc_hs__nand3_2 _29344_ (.A(net216),
    .B(_22831_),
    .C(_22832_),
    .Y(_22833_));
 sky130_as_sc_hs__or2_2 _29345_ (.A(net388),
    .B(\tholin_riscv.regs[18][12] ),
    .Y(_22834_));
 sky130_as_sc_hs__or2_2 _29346_ (.A(net208),
    .B(\tholin_riscv.regs[19][12] ),
    .Y(_22835_));
 sky130_as_sc_hs__nand3_2 _29347_ (.A(net356),
    .B(_22834_),
    .C(_22835_),
    .Y(_22836_));
 sky130_as_sc_hs__nand3_2 _29348_ (.A(net233),
    .B(_22833_),
    .C(_22836_),
    .Y(_22837_));
 sky130_as_sc_hs__or2_2 _29349_ (.A(net388),
    .B(\tholin_riscv.regs[22][12] ),
    .Y(_22838_));
 sky130_as_sc_hs__or2_2 _29350_ (.A(net208),
    .B(\tholin_riscv.regs[23][12] ),
    .Y(_22839_));
 sky130_as_sc_hs__nand3_2 _29351_ (.A(net356),
    .B(_22838_),
    .C(_22839_),
    .Y(_22840_));
 sky130_as_sc_hs__or2_2 _29352_ (.A(net389),
    .B(\tholin_riscv.regs[20][12] ),
    .Y(_22841_));
 sky130_as_sc_hs__or2_2 _29353_ (.A(net207),
    .B(\tholin_riscv.regs[21][12] ),
    .Y(_22842_));
 sky130_as_sc_hs__nand3_2 _29354_ (.A(net216),
    .B(_22841_),
    .C(_22842_),
    .Y(_22843_));
 sky130_as_sc_hs__nand3_2 _29355_ (.A(net344),
    .B(_22840_),
    .C(_22843_),
    .Y(_22844_));
 sky130_as_sc_hs__nand3_2 _29356_ (.A(net241),
    .B(_22837_),
    .C(_22844_),
    .Y(_22845_));
 sky130_as_sc_hs__nand3_2 _29357_ (.A(net338),
    .B(_22823_),
    .C(_22830_),
    .Y(_22846_));
 sky130_as_sc_hs__nand3_2 _29358_ (.A(net336),
    .B(_22845_),
    .C(_22846_),
    .Y(_22847_));
 sky130_as_sc_hs__or2_2 _29359_ (.A(net389),
    .B(\tholin_riscv.regs[8][12] ),
    .Y(_22848_));
 sky130_as_sc_hs__or2_2 _29360_ (.A(net207),
    .B(\tholin_riscv.regs[9][12] ),
    .Y(_22849_));
 sky130_as_sc_hs__nand3_2 _29361_ (.A(net218),
    .B(_22848_),
    .C(_22849_),
    .Y(_22850_));
 sky130_as_sc_hs__or2_2 _29362_ (.A(net393),
    .B(\tholin_riscv.regs[10][12] ),
    .Y(_22851_));
 sky130_as_sc_hs__or2_2 _29363_ (.A(net208),
    .B(\tholin_riscv.regs[11][12] ),
    .Y(_22852_));
 sky130_as_sc_hs__nand3_2 _29364_ (.A(net357),
    .B(_22851_),
    .C(_22852_),
    .Y(_22853_));
 sky130_as_sc_hs__nand3_2 _29365_ (.A(net234),
    .B(_22850_),
    .C(_22853_),
    .Y(_22854_));
 sky130_as_sc_hs__or2_2 _29366_ (.A(net389),
    .B(\tholin_riscv.regs[12][12] ),
    .Y(_22855_));
 sky130_as_sc_hs__or2_2 _29367_ (.A(net209),
    .B(\tholin_riscv.regs[13][12] ),
    .Y(_22856_));
 sky130_as_sc_hs__nand3_2 _29368_ (.A(net216),
    .B(_22855_),
    .C(_22856_),
    .Y(_22857_));
 sky130_as_sc_hs__or2_2 _29369_ (.A(net389),
    .B(\tholin_riscv.regs[14][12] ),
    .Y(_22858_));
 sky130_as_sc_hs__or2_2 _29370_ (.A(net207),
    .B(\tholin_riscv.regs[15][12] ),
    .Y(_22859_));
 sky130_as_sc_hs__nand3_2 _29371_ (.A(net356),
    .B(_22858_),
    .C(_22859_),
    .Y(_22860_));
 sky130_as_sc_hs__nand3_2 _29372_ (.A(net344),
    .B(_22857_),
    .C(_22860_),
    .Y(_22861_));
 sky130_as_sc_hs__or2_2 _29373_ (.A(net393),
    .B(\tholin_riscv.regs[0][12] ),
    .Y(_22862_));
 sky130_as_sc_hs__or2_2 _29374_ (.A(net207),
    .B(\tholin_riscv.regs[1][12] ),
    .Y(_22863_));
 sky130_as_sc_hs__nand3_2 _29375_ (.A(net218),
    .B(_22862_),
    .C(_22863_),
    .Y(_22864_));
 sky130_as_sc_hs__or2_2 _29376_ (.A(net393),
    .B(\tholin_riscv.regs[2][12] ),
    .Y(_22865_));
 sky130_as_sc_hs__or2_2 _29377_ (.A(net208),
    .B(\tholin_riscv.regs[3][12] ),
    .Y(_22866_));
 sky130_as_sc_hs__nand3_2 _29378_ (.A(net357),
    .B(_22865_),
    .C(_22866_),
    .Y(_22867_));
 sky130_as_sc_hs__nand3_2 _29379_ (.A(net233),
    .B(_22864_),
    .C(_22867_),
    .Y(_22868_));
 sky130_as_sc_hs__or2_2 _29380_ (.A(net393),
    .B(\tholin_riscv.regs[6][12] ),
    .Y(_22869_));
 sky130_as_sc_hs__or2_2 _29381_ (.A(net209),
    .B(\tholin_riscv.regs[7][12] ),
    .Y(_22870_));
 sky130_as_sc_hs__nand3_2 _29382_ (.A(net357),
    .B(_22869_),
    .C(_22870_),
    .Y(_22871_));
 sky130_as_sc_hs__or2_2 _29383_ (.A(net393),
    .B(\tholin_riscv.regs[4][12] ),
    .Y(_22872_));
 sky130_as_sc_hs__or2_2 _29384_ (.A(net209),
    .B(\tholin_riscv.regs[5][12] ),
    .Y(_22873_));
 sky130_as_sc_hs__nand3_2 _29385_ (.A(net218),
    .B(_22872_),
    .C(_22873_),
    .Y(_22874_));
 sky130_as_sc_hs__nand3_2 _29386_ (.A(net345),
    .B(_22871_),
    .C(_22874_),
    .Y(_22875_));
 sky130_as_sc_hs__nand3_2 _29387_ (.A(net241),
    .B(_22868_),
    .C(_22875_),
    .Y(_22876_));
 sky130_as_sc_hs__nand3_2 _29388_ (.A(net338),
    .B(_22854_),
    .C(_22861_),
    .Y(_22877_));
 sky130_as_sc_hs__nand3_2 _29389_ (.A(net245),
    .B(_22876_),
    .C(_22877_),
    .Y(_22878_));
 sky130_as_sc_hs__and2_2 _29391_ (.A(_22815_),
    .B(_22879_),
    .Y(_22880_));
 sky130_as_sc_hs__nand3_2 _29392_ (.A(_22624_),
    .B(_22752_),
    .C(_22880_),
    .Y(_22881_));
 sky130_as_sc_hs__nor2_2 _29393_ (.A(_22367_),
    .B(_22881_),
    .Y(_22882_));
 sky130_as_sc_hs__or2_2 _29394_ (.A(net399),
    .B(\tholin_riscv.regs[24][16] ),
    .Y(_22883_));
 sky130_as_sc_hs__nand3_2 _29396_ (.A(net228),
    .B(_22883_),
    .C(_22884_),
    .Y(_22885_));
 sky130_as_sc_hs__or2_2 _29397_ (.A(net399),
    .B(\tholin_riscv.regs[26][16] ),
    .Y(_22886_));
 sky130_as_sc_hs__nand3_2 _29399_ (.A(net368),
    .B(_22886_),
    .C(_22887_),
    .Y(_22888_));
 sky130_as_sc_hs__nand3_2 _29400_ (.A(net239),
    .B(_22885_),
    .C(_22888_),
    .Y(_22889_));
 sky130_as_sc_hs__or2_2 _29401_ (.A(net399),
    .B(\tholin_riscv.regs[28][16] ),
    .Y(_22890_));
 sky130_as_sc_hs__nand3_2 _29403_ (.A(net228),
    .B(_22890_),
    .C(_22891_),
    .Y(_22892_));
 sky130_as_sc_hs__or2_2 _29404_ (.A(net399),
    .B(\tholin_riscv.regs[30][16] ),
    .Y(_22893_));
 sky130_as_sc_hs__nand3_2 _29406_ (.A(net368),
    .B(_22893_),
    .C(_22894_),
    .Y(_22895_));
 sky130_as_sc_hs__nand3_2 _29407_ (.A(net349),
    .B(_22892_),
    .C(_22895_),
    .Y(_22896_));
 sky130_as_sc_hs__or2_2 _29408_ (.A(net398),
    .B(\tholin_riscv.regs[16][16] ),
    .Y(_22897_));
 sky130_as_sc_hs__nand3_2 _29410_ (.A(net229),
    .B(_22897_),
    .C(_22898_),
    .Y(_22899_));
 sky130_as_sc_hs__or2_2 _29411_ (.A(net399),
    .B(\tholin_riscv.regs[18][16] ),
    .Y(_22900_));
 sky130_as_sc_hs__nand3_2 _29413_ (.A(net368),
    .B(_22900_),
    .C(_22901_),
    .Y(_22902_));
 sky130_as_sc_hs__nand3_2 _29414_ (.A(net239),
    .B(_22899_),
    .C(_22902_),
    .Y(_22903_));
 sky130_as_sc_hs__or2_2 _29415_ (.A(net399),
    .B(\tholin_riscv.regs[22][16] ),
    .Y(_22904_));
 sky130_as_sc_hs__nand3_2 _29417_ (.A(net368),
    .B(_22904_),
    .C(_22905_),
    .Y(_22906_));
 sky130_as_sc_hs__or2_2 _29418_ (.A(net399),
    .B(\tholin_riscv.regs[20][16] ),
    .Y(_22907_));
 sky130_as_sc_hs__nand3_2 _29420_ (.A(net229),
    .B(_22907_),
    .C(_22908_),
    .Y(_22909_));
 sky130_as_sc_hs__nand3_2 _29421_ (.A(net349),
    .B(_22906_),
    .C(_22909_),
    .Y(_22910_));
 sky130_as_sc_hs__nand3_2 _29422_ (.A(net244),
    .B(_22903_),
    .C(_22910_),
    .Y(_22911_));
 sky130_as_sc_hs__nand3_2 _29423_ (.A(net339),
    .B(_22889_),
    .C(_22896_),
    .Y(_22912_));
 sky130_as_sc_hs__nand3_2 _29424_ (.A(\tholin_riscv.Jimm[19] ),
    .B(_22911_),
    .C(_22912_),
    .Y(_22913_));
 sky130_as_sc_hs__or2_2 _29425_ (.A(net407),
    .B(\tholin_riscv.regs[8][16] ),
    .Y(_22914_));
 sky130_as_sc_hs__nand3_2 _29427_ (.A(net229),
    .B(_22914_),
    .C(_22915_),
    .Y(_22916_));
 sky130_as_sc_hs__or2_2 _29428_ (.A(net407),
    .B(\tholin_riscv.regs[10][16] ),
    .Y(_22917_));
 sky130_as_sc_hs__nand3_2 _29430_ (.A(net369),
    .B(_22917_),
    .C(_22918_),
    .Y(_22919_));
 sky130_as_sc_hs__nand3_2 _29431_ (.A(net238),
    .B(_22916_),
    .C(_22919_),
    .Y(_22920_));
 sky130_as_sc_hs__or2_2 _29432_ (.A(net407),
    .B(\tholin_riscv.regs[12][16] ),
    .Y(_22921_));
 sky130_as_sc_hs__nand3_2 _29434_ (.A(net229),
    .B(_22921_),
    .C(_22922_),
    .Y(_22923_));
 sky130_as_sc_hs__or2_2 _29435_ (.A(net407),
    .B(\tholin_riscv.regs[14][16] ),
    .Y(_22924_));
 sky130_as_sc_hs__nand3_2 _29437_ (.A(net369),
    .B(_22924_),
    .C(_22925_),
    .Y(_22926_));
 sky130_as_sc_hs__nand3_2 _29438_ (.A(net350),
    .B(_22923_),
    .C(_22926_),
    .Y(_22927_));
 sky130_as_sc_hs__or2_2 _29439_ (.A(net407),
    .B(\tholin_riscv.regs[0][16] ),
    .Y(_22928_));
 sky130_as_sc_hs__nand3_2 _29441_ (.A(net229),
    .B(_22928_),
    .C(_22929_),
    .Y(_22930_));
 sky130_as_sc_hs__or2_2 _29442_ (.A(net407),
    .B(\tholin_riscv.regs[2][16] ),
    .Y(_22931_));
 sky130_as_sc_hs__nand3_2 _29444_ (.A(net369),
    .B(_22931_),
    .C(_22932_),
    .Y(_22933_));
 sky130_as_sc_hs__nand3_2 _29445_ (.A(net238),
    .B(_22930_),
    .C(_22933_),
    .Y(_22934_));
 sky130_as_sc_hs__or2_2 _29446_ (.A(net407),
    .B(\tholin_riscv.regs[6][16] ),
    .Y(_22935_));
 sky130_as_sc_hs__nand3_2 _29448_ (.A(net369),
    .B(_22935_),
    .C(_22936_),
    .Y(_22937_));
 sky130_as_sc_hs__or2_2 _29449_ (.A(net408),
    .B(\tholin_riscv.regs[4][16] ),
    .Y(_22938_));
 sky130_as_sc_hs__nand3_2 _29451_ (.A(net229),
    .B(_22938_),
    .C(_22939_),
    .Y(_22940_));
 sky130_as_sc_hs__nand3_2 _29452_ (.A(net349),
    .B(_22937_),
    .C(_22940_),
    .Y(_22941_));
 sky130_as_sc_hs__nand3_2 _29453_ (.A(net243),
    .B(_22934_),
    .C(_22941_),
    .Y(_22942_));
 sky130_as_sc_hs__nand3_2 _29454_ (.A(net341),
    .B(_22920_),
    .C(_22927_),
    .Y(_22943_));
 sky130_as_sc_hs__nand3_2 _29455_ (.A(net245),
    .B(_22942_),
    .C(_22943_),
    .Y(_22944_));
 sky130_as_sc_hs__nor2_2 _29458_ (.A(_21851_),
    .B(_22946_),
    .Y(_22947_));
 sky130_as_sc_hs__nand3_2 _29459_ (.A(_21850_),
    .B(_22882_),
    .C(_22945_),
    .Y(_22948_));
 sky130_as_sc_hs__or2_2 _29460_ (.A(net397),
    .B(\tholin_riscv.regs[24][18] ),
    .Y(_22949_));
 sky130_as_sc_hs__nand3_2 _29462_ (.A(net224),
    .B(_22949_),
    .C(_22950_),
    .Y(_22951_));
 sky130_as_sc_hs__or2_2 _29463_ (.A(net400),
    .B(\tholin_riscv.regs[26][18] ),
    .Y(_22952_));
 sky130_as_sc_hs__nand3_2 _29465_ (.A(net363),
    .B(_22952_),
    .C(_22953_),
    .Y(_22954_));
 sky130_as_sc_hs__nand3_2 _29466_ (.A(net235),
    .B(_22951_),
    .C(_22954_),
    .Y(_22955_));
 sky130_as_sc_hs__or2_2 _29467_ (.A(net397),
    .B(\tholin_riscv.regs[28][18] ),
    .Y(_22956_));
 sky130_as_sc_hs__nand3_2 _29469_ (.A(net224),
    .B(_22956_),
    .C(_22957_),
    .Y(_22958_));
 sky130_as_sc_hs__or2_2 _29470_ (.A(net400),
    .B(\tholin_riscv.regs[30][18] ),
    .Y(_22959_));
 sky130_as_sc_hs__nand3_2 _29472_ (.A(net362),
    .B(_22959_),
    .C(_22960_),
    .Y(_22961_));
 sky130_as_sc_hs__nand3_2 _29473_ (.A(net346),
    .B(_22958_),
    .C(_22961_),
    .Y(_22962_));
 sky130_as_sc_hs__or2_2 _29474_ (.A(net397),
    .B(\tholin_riscv.regs[16][18] ),
    .Y(_22963_));
 sky130_as_sc_hs__nand3_2 _29476_ (.A(net222),
    .B(_22963_),
    .C(_22964_),
    .Y(_22965_));
 sky130_as_sc_hs__or2_2 _29477_ (.A(net397),
    .B(\tholin_riscv.regs[18][18] ),
    .Y(_22966_));
 sky130_as_sc_hs__nand3_2 _29479_ (.A(net362),
    .B(_22966_),
    .C(_22967_),
    .Y(_22968_));
 sky130_as_sc_hs__nand3_2 _29480_ (.A(net235),
    .B(_22965_),
    .C(_22968_),
    .Y(_22969_));
 sky130_as_sc_hs__or2_2 _29481_ (.A(net397),
    .B(\tholin_riscv.regs[22][18] ),
    .Y(_22970_));
 sky130_as_sc_hs__nand3_2 _29483_ (.A(net363),
    .B(_22970_),
    .C(_22971_),
    .Y(_22972_));
 sky130_as_sc_hs__or2_2 _29484_ (.A(net397),
    .B(\tholin_riscv.regs[20][18] ),
    .Y(_22973_));
 sky130_as_sc_hs__nand3_2 _29486_ (.A(net222),
    .B(_22973_),
    .C(_22974_),
    .Y(_22975_));
 sky130_as_sc_hs__nand3_2 _29487_ (.A(net346),
    .B(_22972_),
    .C(_22975_),
    .Y(_22976_));
 sky130_as_sc_hs__nand3_2 _29488_ (.A(net242),
    .B(_22969_),
    .C(_22976_),
    .Y(_22977_));
 sky130_as_sc_hs__nand3_2 _29489_ (.A(net340),
    .B(_22955_),
    .C(_22962_),
    .Y(_22978_));
 sky130_as_sc_hs__nand3_2 _29490_ (.A(net335),
    .B(_22977_),
    .C(_22978_),
    .Y(_22979_));
 sky130_as_sc_hs__or2_2 _29491_ (.A(net402),
    .B(\tholin_riscv.regs[8][18] ),
    .Y(_22980_));
 sky130_as_sc_hs__nand3_2 _29493_ (.A(net226),
    .B(_22980_),
    .C(_22981_),
    .Y(_22982_));
 sky130_as_sc_hs__or2_2 _29494_ (.A(net396),
    .B(\tholin_riscv.regs[10][18] ),
    .Y(_22983_));
 sky130_as_sc_hs__nand3_2 _29496_ (.A(net364),
    .B(_22983_),
    .C(_22984_),
    .Y(_22985_));
 sky130_as_sc_hs__nand3_2 _29497_ (.A(net237),
    .B(_22982_),
    .C(_22985_),
    .Y(_22986_));
 sky130_as_sc_hs__or2_2 _29498_ (.A(net402),
    .B(\tholin_riscv.regs[12][18] ),
    .Y(_22987_));
 sky130_as_sc_hs__nand3_2 _29500_ (.A(net228),
    .B(_22987_),
    .C(_22988_),
    .Y(_22989_));
 sky130_as_sc_hs__or2_2 _29501_ (.A(net402),
    .B(\tholin_riscv.regs[14][18] ),
    .Y(_22990_));
 sky130_as_sc_hs__nand3_2 _29503_ (.A(net364),
    .B(_22990_),
    .C(_22991_),
    .Y(_22992_));
 sky130_as_sc_hs__nand3_2 _29504_ (.A(net348),
    .B(_22989_),
    .C(_22992_),
    .Y(_22993_));
 sky130_as_sc_hs__or2_2 _29505_ (.A(net402),
    .B(\tholin_riscv.regs[0][18] ),
    .Y(_22994_));
 sky130_as_sc_hs__nand3_2 _29507_ (.A(net226),
    .B(_22994_),
    .C(_22995_),
    .Y(_22996_));
 sky130_as_sc_hs__or2_2 _29508_ (.A(net402),
    .B(\tholin_riscv.regs[2][18] ),
    .Y(_22997_));
 sky130_as_sc_hs__nand3_2 _29510_ (.A(net370),
    .B(_22997_),
    .C(_22998_),
    .Y(_22999_));
 sky130_as_sc_hs__nand3_2 _29511_ (.A(net237),
    .B(_22996_),
    .C(_22999_),
    .Y(_23000_));
 sky130_as_sc_hs__or2_2 _29512_ (.A(net402),
    .B(\tholin_riscv.regs[6][18] ),
    .Y(_23001_));
 sky130_as_sc_hs__nand3_2 _29514_ (.A(net364),
    .B(_23001_),
    .C(_23002_),
    .Y(_23003_));
 sky130_as_sc_hs__or2_2 _29515_ (.A(net402),
    .B(\tholin_riscv.regs[4][18] ),
    .Y(_23004_));
 sky130_as_sc_hs__nand3_2 _29517_ (.A(net226),
    .B(_23004_),
    .C(_23005_),
    .Y(_23006_));
 sky130_as_sc_hs__nand3_2 _29518_ (.A(net348),
    .B(_23003_),
    .C(_23006_),
    .Y(_23007_));
 sky130_as_sc_hs__nand3_2 _29519_ (.A(net243),
    .B(_23000_),
    .C(_23007_),
    .Y(_23008_));
 sky130_as_sc_hs__nand3_2 _29520_ (.A(net339),
    .B(_22986_),
    .C(_22993_),
    .Y(_23009_));
 sky130_as_sc_hs__nand3_2 _29521_ (.A(_19481_),
    .B(_23008_),
    .C(_23009_),
    .Y(_23010_));
 sky130_as_sc_hs__nor2_2 _29525_ (.A(_22948_),
    .B(_23013_),
    .Y(_23014_));
 sky130_as_sc_hs__or2_2 _29526_ (.A(net382),
    .B(\tholin_riscv.regs[24][22] ),
    .Y(_23015_));
 sky130_as_sc_hs__nand3_2 _29528_ (.A(net223),
    .B(_23015_),
    .C(_23016_),
    .Y(_23017_));
 sky130_as_sc_hs__or2_2 _29529_ (.A(net382),
    .B(\tholin_riscv.regs[26][22] ),
    .Y(_23018_));
 sky130_as_sc_hs__nand3_2 _29531_ (.A(net363),
    .B(_23018_),
    .C(_23019_),
    .Y(_23020_));
 sky130_as_sc_hs__nand3_2 _29532_ (.A(net235),
    .B(_23017_),
    .C(_23020_),
    .Y(_23021_));
 sky130_as_sc_hs__or2_2 _29533_ (.A(net380),
    .B(\tholin_riscv.regs[28][22] ),
    .Y(_23022_));
 sky130_as_sc_hs__nand3_2 _29535_ (.A(net222),
    .B(_23022_),
    .C(_23023_),
    .Y(_23024_));
 sky130_as_sc_hs__or2_2 _29536_ (.A(net380),
    .B(\tholin_riscv.regs[30][22] ),
    .Y(_23025_));
 sky130_as_sc_hs__nand3_2 _29538_ (.A(net363),
    .B(_23025_),
    .C(_23026_),
    .Y(_23027_));
 sky130_as_sc_hs__nand3_2 _29539_ (.A(net346),
    .B(_23024_),
    .C(_23027_),
    .Y(_23028_));
 sky130_as_sc_hs__or2_2 _29540_ (.A(net380),
    .B(\tholin_riscv.regs[16][22] ),
    .Y(_23029_));
 sky130_as_sc_hs__nand3_2 _29542_ (.A(net224),
    .B(_23029_),
    .C(_23030_),
    .Y(_23031_));
 sky130_as_sc_hs__or2_2 _29543_ (.A(net380),
    .B(\tholin_riscv.regs[18][22] ),
    .Y(_23032_));
 sky130_as_sc_hs__nand3_2 _29545_ (.A(net363),
    .B(_23032_),
    .C(_23033_),
    .Y(_23034_));
 sky130_as_sc_hs__nand3_2 _29546_ (.A(net235),
    .B(_23031_),
    .C(_23034_),
    .Y(_23035_));
 sky130_as_sc_hs__or2_2 _29547_ (.A(net380),
    .B(\tholin_riscv.regs[22][22] ),
    .Y(_23036_));
 sky130_as_sc_hs__nand3_2 _29549_ (.A(net362),
    .B(_23036_),
    .C(_23037_),
    .Y(_23038_));
 sky130_as_sc_hs__or2_2 _29550_ (.A(net380),
    .B(\tholin_riscv.regs[20][22] ),
    .Y(_23039_));
 sky130_as_sc_hs__nand3_2 _29552_ (.A(net223),
    .B(_23039_),
    .C(_23040_),
    .Y(_23041_));
 sky130_as_sc_hs__nand3_2 _29553_ (.A(net346),
    .B(_23038_),
    .C(_23041_),
    .Y(_23042_));
 sky130_as_sc_hs__nand3_2 _29554_ (.A(net242),
    .B(_23035_),
    .C(_23042_),
    .Y(_23043_));
 sky130_as_sc_hs__nand3_2 _29555_ (.A(net340),
    .B(_23021_),
    .C(_23028_),
    .Y(_23044_));
 sky130_as_sc_hs__nand3_2 _29556_ (.A(net335),
    .B(_23043_),
    .C(_23044_),
    .Y(_23045_));
 sky130_as_sc_hs__or2_2 _29557_ (.A(net396),
    .B(\tholin_riscv.regs[8][22] ),
    .Y(_23046_));
 sky130_as_sc_hs__nand3_2 _29559_ (.A(net225),
    .B(_23046_),
    .C(_23047_),
    .Y(_23048_));
 sky130_as_sc_hs__or2_2 _29560_ (.A(net396),
    .B(\tholin_riscv.regs[10][22] ),
    .Y(_23049_));
 sky130_as_sc_hs__nand3_2 _29562_ (.A(net365),
    .B(_23049_),
    .C(_23050_),
    .Y(_23051_));
 sky130_as_sc_hs__nand3_2 _29563_ (.A(net237),
    .B(_23048_),
    .C(_23051_),
    .Y(_23052_));
 sky130_as_sc_hs__or2_2 _29564_ (.A(net398),
    .B(\tholin_riscv.regs[12][22] ),
    .Y(_23053_));
 sky130_as_sc_hs__nand3_2 _29566_ (.A(net228),
    .B(_23053_),
    .C(_23054_),
    .Y(_23055_));
 sky130_as_sc_hs__or2_2 _29567_ (.A(net398),
    .B(\tholin_riscv.regs[14][22] ),
    .Y(_23056_));
 sky130_as_sc_hs__nand3_2 _29569_ (.A(net367),
    .B(_23056_),
    .C(_23057_),
    .Y(_23058_));
 sky130_as_sc_hs__nand3_2 _29570_ (.A(net349),
    .B(_23055_),
    .C(_23058_),
    .Y(_23059_));
 sky130_as_sc_hs__or2_2 _29571_ (.A(net396),
    .B(\tholin_riscv.regs[0][22] ),
    .Y(_23060_));
 sky130_as_sc_hs__nand3_2 _29573_ (.A(net228),
    .B(_23060_),
    .C(_23061_),
    .Y(_23062_));
 sky130_as_sc_hs__or2_2 _29574_ (.A(net398),
    .B(\tholin_riscv.regs[2][22] ),
    .Y(_23063_));
 sky130_as_sc_hs__nand3_2 _29576_ (.A(net367),
    .B(_23063_),
    .C(_23064_),
    .Y(_23065_));
 sky130_as_sc_hs__nand3_2 _29577_ (.A(net239),
    .B(_23062_),
    .C(_23065_),
    .Y(_23066_));
 sky130_as_sc_hs__or2_2 _29578_ (.A(net398),
    .B(\tholin_riscv.regs[6][22] ),
    .Y(_23067_));
 sky130_as_sc_hs__nand3_2 _29580_ (.A(net367),
    .B(_23067_),
    .C(_23068_),
    .Y(_23069_));
 sky130_as_sc_hs__or2_2 _29581_ (.A(net398),
    .B(\tholin_riscv.regs[4][22] ),
    .Y(_23070_));
 sky130_as_sc_hs__nand3_2 _29583_ (.A(net228),
    .B(_23070_),
    .C(_23071_),
    .Y(_23072_));
 sky130_as_sc_hs__nand3_2 _29584_ (.A(net349),
    .B(_23069_),
    .C(_23072_),
    .Y(_23073_));
 sky130_as_sc_hs__nand3_2 _29585_ (.A(net243),
    .B(_23066_),
    .C(_23073_),
    .Y(_23074_));
 sky130_as_sc_hs__nand3_2 _29586_ (.A(net339),
    .B(_23052_),
    .C(_23059_),
    .Y(_23075_));
 sky130_as_sc_hs__nand3_2 _29587_ (.A(net245),
    .B(_23074_),
    .C(_23075_),
    .Y(_23076_));
 sky130_as_sc_hs__inv_2 _29589_ (.Y(_23078_),
    .A(_23077_));
 sky130_as_sc_hs__or2_2 _29590_ (.A(net381),
    .B(\tholin_riscv.regs[24][23] ),
    .Y(_23079_));
 sky130_as_sc_hs__nand3_2 _29592_ (.A(net223),
    .B(_23079_),
    .C(_23080_),
    .Y(_23081_));
 sky130_as_sc_hs__or2_2 _29593_ (.A(net381),
    .B(\tholin_riscv.regs[26][23] ),
    .Y(_23082_));
 sky130_as_sc_hs__nand3_2 _29595_ (.A(net362),
    .B(_23082_),
    .C(_23083_),
    .Y(_23084_));
 sky130_as_sc_hs__nand3_2 _29596_ (.A(net235),
    .B(_23081_),
    .C(_23084_),
    .Y(_23085_));
 sky130_as_sc_hs__or2_2 _29597_ (.A(net378),
    .B(\tholin_riscv.regs[28][23] ),
    .Y(_23086_));
 sky130_as_sc_hs__nand3_2 _29599_ (.A(net223),
    .B(_23086_),
    .C(_23087_),
    .Y(_23088_));
 sky130_as_sc_hs__or2_2 _29600_ (.A(net378),
    .B(\tholin_riscv.regs[30][23] ),
    .Y(_23089_));
 sky130_as_sc_hs__nand3_2 _29602_ (.A(net363),
    .B(_23089_),
    .C(_23090_),
    .Y(_23091_));
 sky130_as_sc_hs__nand3_2 _29603_ (.A(net346),
    .B(_23088_),
    .C(_23091_),
    .Y(_23092_));
 sky130_as_sc_hs__or2_2 _29604_ (.A(net376),
    .B(\tholin_riscv.regs[16][23] ),
    .Y(_23093_));
 sky130_as_sc_hs__nand3_2 _29606_ (.A(net221),
    .B(_23093_),
    .C(_23094_),
    .Y(_23095_));
 sky130_as_sc_hs__or2_2 _29607_ (.A(net376),
    .B(\tholin_riscv.regs[18][23] ),
    .Y(_23096_));
 sky130_as_sc_hs__nand3_2 _29609_ (.A(net361),
    .B(_23096_),
    .C(_23097_),
    .Y(_23098_));
 sky130_as_sc_hs__nand3_2 _29610_ (.A(net236),
    .B(_23095_),
    .C(_23098_),
    .Y(_23099_));
 sky130_as_sc_hs__or2_2 _29611_ (.A(net377),
    .B(\tholin_riscv.regs[22][23] ),
    .Y(_23100_));
 sky130_as_sc_hs__nand3_2 _29613_ (.A(net360),
    .B(_23100_),
    .C(_23101_),
    .Y(_23102_));
 sky130_as_sc_hs__or2_2 _29614_ (.A(net376),
    .B(\tholin_riscv.regs[20][23] ),
    .Y(_23103_));
 sky130_as_sc_hs__nand3_2 _29616_ (.A(net221),
    .B(_23103_),
    .C(_23104_),
    .Y(_23105_));
 sky130_as_sc_hs__nand3_2 _29617_ (.A(net347),
    .B(_23102_),
    .C(_23105_),
    .Y(_23106_));
 sky130_as_sc_hs__nand3_2 _29618_ (.A(net242),
    .B(_23099_),
    .C(_23106_),
    .Y(_23107_));
 sky130_as_sc_hs__nand3_2 _29619_ (.A(net340),
    .B(_23085_),
    .C(_23092_),
    .Y(_23108_));
 sky130_as_sc_hs__nand3_2 _29620_ (.A(net335),
    .B(_23107_),
    .C(_23108_),
    .Y(_23109_));
 sky130_as_sc_hs__or2_2 _29621_ (.A(net375),
    .B(\tholin_riscv.regs[8][23] ),
    .Y(_23110_));
 sky130_as_sc_hs__nand3_2 _29623_ (.A(net220),
    .B(_23110_),
    .C(_23111_),
    .Y(_23112_));
 sky130_as_sc_hs__or2_2 _29624_ (.A(net395),
    .B(\tholin_riscv.regs[10][23] ),
    .Y(_23113_));
 sky130_as_sc_hs__nand3_2 _29626_ (.A(net361),
    .B(_23113_),
    .C(_23114_),
    .Y(_23115_));
 sky130_as_sc_hs__nand3_2 _29627_ (.A(net236),
    .B(_23112_),
    .C(_23115_),
    .Y(_23116_));
 sky130_as_sc_hs__or2_2 _29628_ (.A(net397),
    .B(\tholin_riscv.regs[12][23] ),
    .Y(_23117_));
 sky130_as_sc_hs__nand3_2 _29630_ (.A(net222),
    .B(_23117_),
    .C(_23118_),
    .Y(_23119_));
 sky130_as_sc_hs__or2_2 _29631_ (.A(net381),
    .B(\tholin_riscv.regs[14][23] ),
    .Y(_23120_));
 sky130_as_sc_hs__nand3_2 _29633_ (.A(net362),
    .B(_23120_),
    .C(_23121_),
    .Y(_23122_));
 sky130_as_sc_hs__nand3_2 _29634_ (.A(net346),
    .B(_23119_),
    .C(_23122_),
    .Y(_23123_));
 sky130_as_sc_hs__or2_2 _29635_ (.A(net376),
    .B(\tholin_riscv.regs[0][23] ),
    .Y(_23124_));
 sky130_as_sc_hs__nand3_2 _29637_ (.A(net220),
    .B(_23124_),
    .C(_23125_),
    .Y(_23126_));
 sky130_as_sc_hs__or2_2 _29638_ (.A(net376),
    .B(\tholin_riscv.regs[2][23] ),
    .Y(_23127_));
 sky130_as_sc_hs__nand3_2 _29640_ (.A(net360),
    .B(_23127_),
    .C(_23128_),
    .Y(_23129_));
 sky130_as_sc_hs__nand3_2 _29641_ (.A(net236),
    .B(_23126_),
    .C(_23129_),
    .Y(_23130_));
 sky130_as_sc_hs__or2_2 _29642_ (.A(net376),
    .B(\tholin_riscv.regs[6][23] ),
    .Y(_23131_));
 sky130_as_sc_hs__nand3_2 _29644_ (.A(net361),
    .B(_23131_),
    .C(_23132_),
    .Y(_23133_));
 sky130_as_sc_hs__or2_2 _29645_ (.A(net381),
    .B(\tholin_riscv.regs[4][23] ),
    .Y(_23134_));
 sky130_as_sc_hs__nand3_2 _29647_ (.A(net223),
    .B(_23134_),
    .C(_23135_),
    .Y(_23136_));
 sky130_as_sc_hs__nand3_2 _29648_ (.A(net347),
    .B(_23133_),
    .C(_23136_),
    .Y(_23137_));
 sky130_as_sc_hs__nand3_2 _29649_ (.A(net242),
    .B(_23130_),
    .C(_23137_),
    .Y(_23138_));
 sky130_as_sc_hs__nand3_2 _29650_ (.A(net340),
    .B(_23116_),
    .C(_23123_),
    .Y(_23139_));
 sky130_as_sc_hs__nand3_2 _29651_ (.A(net246),
    .B(_23138_),
    .C(_23139_),
    .Y(_23140_));
 sky130_as_sc_hs__and2_2 _29652_ (.A(_23109_),
    .B(_23140_),
    .Y(_23141_));
 sky130_as_sc_hs__or2_2 _29653_ (.A(net398),
    .B(\tholin_riscv.regs[24][21] ),
    .Y(_23142_));
 sky130_as_sc_hs__nand3_2 _29655_ (.A(net228),
    .B(_23142_),
    .C(_23143_),
    .Y(_23144_));
 sky130_as_sc_hs__or2_2 _29656_ (.A(net398),
    .B(\tholin_riscv.regs[26][21] ),
    .Y(_23145_));
 sky130_as_sc_hs__nand3_2 _29658_ (.A(net367),
    .B(_23145_),
    .C(_23146_),
    .Y(_23147_));
 sky130_as_sc_hs__nand3_2 _29659_ (.A(net239),
    .B(_23144_),
    .C(_23147_),
    .Y(_23148_));
 sky130_as_sc_hs__or2_2 _29660_ (.A(net399),
    .B(\tholin_riscv.regs[28][21] ),
    .Y(_23149_));
 sky130_as_sc_hs__nand3_2 _29662_ (.A(net228),
    .B(_23149_),
    .C(_23150_),
    .Y(_23151_));
 sky130_as_sc_hs__or2_2 _29663_ (.A(net406),
    .B(\tholin_riscv.regs[30][21] ),
    .Y(_23152_));
 sky130_as_sc_hs__nand3_2 _29665_ (.A(net367),
    .B(_23152_),
    .C(_23153_),
    .Y(_23154_));
 sky130_as_sc_hs__nand3_2 _29666_ (.A(net349),
    .B(_23151_),
    .C(_23154_),
    .Y(_23155_));
 sky130_as_sc_hs__or2_2 _29667_ (.A(net405),
    .B(\tholin_riscv.regs[16][21] ),
    .Y(_23156_));
 sky130_as_sc_hs__nand3_2 _29669_ (.A(net228),
    .B(_23156_),
    .C(_23157_),
    .Y(_23158_));
 sky130_as_sc_hs__or2_2 _29670_ (.A(net405),
    .B(\tholin_riscv.regs[18][21] ),
    .Y(_23159_));
 sky130_as_sc_hs__nand3_2 _29672_ (.A(net367),
    .B(_23159_),
    .C(_23160_),
    .Y(_23161_));
 sky130_as_sc_hs__nand3_2 _29673_ (.A(net238),
    .B(_23158_),
    .C(_23161_),
    .Y(_23162_));
 sky130_as_sc_hs__or2_2 _29674_ (.A(net405),
    .B(\tholin_riscv.regs[22][21] ),
    .Y(_23163_));
 sky130_as_sc_hs__nand3_2 _29676_ (.A(net369),
    .B(_23163_),
    .C(_23164_),
    .Y(_23165_));
 sky130_as_sc_hs__or2_2 _29677_ (.A(net405),
    .B(\tholin_riscv.regs[20][21] ),
    .Y(_23166_));
 sky130_as_sc_hs__nand3_2 _29679_ (.A(net229),
    .B(_23166_),
    .C(_23167_),
    .Y(_23168_));
 sky130_as_sc_hs__nand3_2 _29680_ (.A(net349),
    .B(_23165_),
    .C(_23168_),
    .Y(_23169_));
 sky130_as_sc_hs__nand3_2 _29681_ (.A(net243),
    .B(_23162_),
    .C(_23169_),
    .Y(_23170_));
 sky130_as_sc_hs__nand3_2 _29682_ (.A(net341),
    .B(_23148_),
    .C(_23155_),
    .Y(_23171_));
 sky130_as_sc_hs__nand3_2 _29683_ (.A(net335),
    .B(_23170_),
    .C(_23171_),
    .Y(_23172_));
 sky130_as_sc_hs__or2_2 _29684_ (.A(net404),
    .B(\tholin_riscv.regs[8][21] ),
    .Y(_23173_));
 sky130_as_sc_hs__nand3_2 _29686_ (.A(net227),
    .B(_23173_),
    .C(_23174_),
    .Y(_23175_));
 sky130_as_sc_hs__or2_2 _29687_ (.A(net404),
    .B(\tholin_riscv.regs[10][21] ),
    .Y(_23176_));
 sky130_as_sc_hs__nand3_2 _29689_ (.A(net366),
    .B(_23176_),
    .C(_23177_),
    .Y(_23178_));
 sky130_as_sc_hs__nand3_2 _29690_ (.A(net238),
    .B(_23175_),
    .C(_23178_),
    .Y(_23179_));
 sky130_as_sc_hs__or2_2 _29691_ (.A(net404),
    .B(\tholin_riscv.regs[12][21] ),
    .Y(_23180_));
 sky130_as_sc_hs__nand3_2 _29693_ (.A(net227),
    .B(_23180_),
    .C(_23181_),
    .Y(_23182_));
 sky130_as_sc_hs__or2_2 _29694_ (.A(net404),
    .B(\tholin_riscv.regs[14][21] ),
    .Y(_23183_));
 sky130_as_sc_hs__nand3_2 _29696_ (.A(net366),
    .B(_23183_),
    .C(_23184_),
    .Y(_23185_));
 sky130_as_sc_hs__nand3_2 _29697_ (.A(net348),
    .B(_23182_),
    .C(_23185_),
    .Y(_23186_));
 sky130_as_sc_hs__or2_2 _29698_ (.A(net404),
    .B(\tholin_riscv.regs[0][21] ),
    .Y(_23187_));
 sky130_as_sc_hs__nand3_2 _29700_ (.A(net227),
    .B(_23187_),
    .C(_23188_),
    .Y(_23189_));
 sky130_as_sc_hs__or2_2 _29701_ (.A(net404),
    .B(\tholin_riscv.regs[2][21] ),
    .Y(_23190_));
 sky130_as_sc_hs__nand3_2 _29703_ (.A(net366),
    .B(_23190_),
    .C(_23191_),
    .Y(_23192_));
 sky130_as_sc_hs__nand3_2 _29704_ (.A(net238),
    .B(_23189_),
    .C(_23192_),
    .Y(_23193_));
 sky130_as_sc_hs__or2_2 _29705_ (.A(net404),
    .B(\tholin_riscv.regs[6][21] ),
    .Y(_23194_));
 sky130_as_sc_hs__nand3_2 _29707_ (.A(net366),
    .B(_23194_),
    .C(_23195_),
    .Y(_23196_));
 sky130_as_sc_hs__or2_2 _29708_ (.A(net404),
    .B(\tholin_riscv.regs[4][21] ),
    .Y(_23197_));
 sky130_as_sc_hs__nand3_2 _29710_ (.A(net227),
    .B(_23197_),
    .C(_23198_),
    .Y(_23199_));
 sky130_as_sc_hs__nand3_2 _29711_ (.A(net348),
    .B(_23196_),
    .C(_23199_),
    .Y(_23200_));
 sky130_as_sc_hs__nand3_2 _29712_ (.A(net243),
    .B(_23193_),
    .C(_23200_),
    .Y(_23201_));
 sky130_as_sc_hs__nand3_2 _29713_ (.A(net339),
    .B(_23179_),
    .C(_23186_),
    .Y(_23202_));
 sky130_as_sc_hs__nand3_2 _29714_ (.A(net245),
    .B(_23201_),
    .C(_23202_),
    .Y(_23203_));
 sky130_as_sc_hs__inv_2 _29716_ (.Y(_23205_),
    .A(_23204_));
 sky130_as_sc_hs__or2_2 _29717_ (.A(net398),
    .B(\tholin_riscv.regs[24][20] ),
    .Y(_23206_));
 sky130_as_sc_hs__nand3_2 _29719_ (.A(net228),
    .B(_23206_),
    .C(_23207_),
    .Y(_23208_));
 sky130_as_sc_hs__or2_2 _29720_ (.A(net398),
    .B(\tholin_riscv.regs[26][20] ),
    .Y(_23209_));
 sky130_as_sc_hs__nand3_2 _29722_ (.A(net367),
    .B(_23209_),
    .C(_23210_),
    .Y(_23211_));
 sky130_as_sc_hs__nand3_2 _29723_ (.A(net238),
    .B(_23208_),
    .C(_23211_),
    .Y(_23212_));
 sky130_as_sc_hs__or2_2 _29724_ (.A(net398),
    .B(\tholin_riscv.regs[28][20] ),
    .Y(_23213_));
 sky130_as_sc_hs__nand3_2 _29726_ (.A(net228),
    .B(_23213_),
    .C(_23214_),
    .Y(_23215_));
 sky130_as_sc_hs__or2_2 _29727_ (.A(net398),
    .B(\tholin_riscv.regs[30][20] ),
    .Y(_23216_));
 sky130_as_sc_hs__nand3_2 _29729_ (.A(net367),
    .B(_23216_),
    .C(_23217_),
    .Y(_23218_));
 sky130_as_sc_hs__nand3_2 _29730_ (.A(net349),
    .B(_23215_),
    .C(_23218_),
    .Y(_23219_));
 sky130_as_sc_hs__or2_2 _29731_ (.A(net397),
    .B(\tholin_riscv.regs[16][20] ),
    .Y(_23220_));
 sky130_as_sc_hs__nand3_2 _29733_ (.A(net224),
    .B(_23220_),
    .C(_23221_),
    .Y(_23222_));
 sky130_as_sc_hs__or2_2 _29734_ (.A(net400),
    .B(\tholin_riscv.regs[18][20] ),
    .Y(_23223_));
 sky130_as_sc_hs__nand3_2 _29736_ (.A(net367),
    .B(_23223_),
    .C(_23224_),
    .Y(_23225_));
 sky130_as_sc_hs__nand3_2 _29737_ (.A(net239),
    .B(_23222_),
    .C(_23225_),
    .Y(_23226_));
 sky130_as_sc_hs__or2_2 _29738_ (.A(net398),
    .B(\tholin_riscv.regs[22][20] ),
    .Y(_23227_));
 sky130_as_sc_hs__nand3_2 _29740_ (.A(net367),
    .B(_23227_),
    .C(_23228_),
    .Y(_23229_));
 sky130_as_sc_hs__or2_2 _29741_ (.A(net398),
    .B(\tholin_riscv.regs[20][20] ),
    .Y(_23230_));
 sky130_as_sc_hs__nand3_2 _29743_ (.A(net222),
    .B(_23230_),
    .C(_23231_),
    .Y(_23232_));
 sky130_as_sc_hs__nand3_2 _29744_ (.A(net349),
    .B(_23229_),
    .C(_23232_),
    .Y(_23233_));
 sky130_as_sc_hs__nand3_2 _29745_ (.A(net243),
    .B(_23226_),
    .C(_23233_),
    .Y(_23234_));
 sky130_as_sc_hs__nand3_2 _29746_ (.A(net341),
    .B(_23212_),
    .C(_23219_),
    .Y(_23235_));
 sky130_as_sc_hs__nand3_2 _29747_ (.A(net335),
    .B(_23234_),
    .C(_23235_),
    .Y(_23236_));
 sky130_as_sc_hs__or2_2 _29748_ (.A(net397),
    .B(\tholin_riscv.regs[8][20] ),
    .Y(_23237_));
 sky130_as_sc_hs__nand3_2 _29750_ (.A(net222),
    .B(_23237_),
    .C(_23238_),
    .Y(_23239_));
 sky130_as_sc_hs__or2_2 _29751_ (.A(net397),
    .B(\tholin_riscv.regs[10][20] ),
    .Y(_23240_));
 sky130_as_sc_hs__nand3_2 _29753_ (.A(net362),
    .B(_23240_),
    .C(_23241_),
    .Y(_23242_));
 sky130_as_sc_hs__nand3_2 _29754_ (.A(net235),
    .B(_23239_),
    .C(_23242_),
    .Y(_23243_));
 sky130_as_sc_hs__or2_2 _29755_ (.A(net397),
    .B(\tholin_riscv.regs[12][20] ),
    .Y(_23244_));
 sky130_as_sc_hs__nand3_2 _29757_ (.A(net222),
    .B(_23244_),
    .C(_23245_),
    .Y(_23246_));
 sky130_as_sc_hs__or2_2 _29758_ (.A(net397),
    .B(\tholin_riscv.regs[14][20] ),
    .Y(_23247_));
 sky130_as_sc_hs__nand3_2 _29760_ (.A(net362),
    .B(_23247_),
    .C(_23248_),
    .Y(_23249_));
 sky130_as_sc_hs__nand3_2 _29761_ (.A(\tholin_riscv.Jimm[17] ),
    .B(_23246_),
    .C(_23249_),
    .Y(_23250_));
 sky130_as_sc_hs__or2_2 _29762_ (.A(net397),
    .B(\tholin_riscv.regs[0][20] ),
    .Y(_23251_));
 sky130_as_sc_hs__nand3_2 _29764_ (.A(net222),
    .B(_23251_),
    .C(_23252_),
    .Y(_23253_));
 sky130_as_sc_hs__or2_2 _29765_ (.A(net397),
    .B(\tholin_riscv.regs[2][20] ),
    .Y(_23254_));
 sky130_as_sc_hs__nand3_2 _29767_ (.A(net362),
    .B(_23254_),
    .C(_23255_),
    .Y(_23256_));
 sky130_as_sc_hs__nand3_2 _29768_ (.A(net235),
    .B(_23253_),
    .C(_23256_),
    .Y(_23257_));
 sky130_as_sc_hs__or2_2 _29769_ (.A(net397),
    .B(\tholin_riscv.regs[6][20] ),
    .Y(_23258_));
 sky130_as_sc_hs__nand3_2 _29771_ (.A(net367),
    .B(_23258_),
    .C(_23259_),
    .Y(_23260_));
 sky130_as_sc_hs__or2_2 _29772_ (.A(net397),
    .B(\tholin_riscv.regs[4][20] ),
    .Y(_23261_));
 sky130_as_sc_hs__nand3_2 _29774_ (.A(net222),
    .B(_23261_),
    .C(_23262_),
    .Y(_23263_));
 sky130_as_sc_hs__nand3_2 _29775_ (.A(net346),
    .B(_23260_),
    .C(_23263_),
    .Y(_23264_));
 sky130_as_sc_hs__nand3_2 _29776_ (.A(net242),
    .B(_23257_),
    .C(_23264_),
    .Y(_23265_));
 sky130_as_sc_hs__nand3_2 _29777_ (.A(net340),
    .B(_23243_),
    .C(_23250_),
    .Y(_23266_));
 sky130_as_sc_hs__nand3_2 _29778_ (.A(net246),
    .B(_23265_),
    .C(_23266_),
    .Y(_23267_));
 sky130_as_sc_hs__nand3_2 _29780_ (.A(_23077_),
    .B(_23204_),
    .C(_23268_),
    .Y(_23269_));
 sky130_as_sc_hs__nor2_2 _29781_ (.A(_23141_),
    .B(_23269_),
    .Y(_23270_));
 sky130_as_sc_hs__and2_2 _29782_ (.A(_23014_),
    .B(_23270_),
    .Y(_23271_));
 sky130_as_sc_hs__nand3_2 _29785_ (.A(net220),
    .B(_23272_),
    .C(_23273_),
    .Y(_23274_));
 sky130_as_sc_hs__nand3_2 _29788_ (.A(net364),
    .B(_23275_),
    .C(_23276_),
    .Y(_23277_));
 sky130_as_sc_hs__nand3_2 _29789_ (.A(net236),
    .B(_23274_),
    .C(_23277_),
    .Y(_23278_));
 sky130_as_sc_hs__nand3_2 _29792_ (.A(net222),
    .B(_23279_),
    .C(_23280_),
    .Y(_23281_));
 sky130_as_sc_hs__nand3_2 _29795_ (.A(net367),
    .B(_23282_),
    .C(_23283_),
    .Y(_23284_));
 sky130_as_sc_hs__nand3_2 _29796_ (.A(net349),
    .B(_23281_),
    .C(_23284_),
    .Y(_23285_));
 sky130_as_sc_hs__nand3_2 _29799_ (.A(net220),
    .B(_23286_),
    .C(_23287_),
    .Y(_23288_));
 sky130_as_sc_hs__nand3_2 _29802_ (.A(net364),
    .B(_23289_),
    .C(_23290_),
    .Y(_23291_));
 sky130_as_sc_hs__nand3_2 _29803_ (.A(net236),
    .B(_23288_),
    .C(_23291_),
    .Y(_23292_));
 sky130_as_sc_hs__nand3_2 _29806_ (.A(net364),
    .B(_23293_),
    .C(_23294_),
    .Y(_23295_));
 sky130_as_sc_hs__nand3_2 _29809_ (.A(net222),
    .B(_23296_),
    .C(_23297_),
    .Y(_23298_));
 sky130_as_sc_hs__nand3_2 _29810_ (.A(net348),
    .B(_23295_),
    .C(_23298_),
    .Y(_23299_));
 sky130_as_sc_hs__nand3_2 _29811_ (.A(net242),
    .B(_23292_),
    .C(_23299_),
    .Y(_23300_));
 sky130_as_sc_hs__nand3_2 _29812_ (.A(net339),
    .B(_23278_),
    .C(_23285_),
    .Y(_23301_));
 sky130_as_sc_hs__nand3_2 _29813_ (.A(net335),
    .B(_23300_),
    .C(_23301_),
    .Y(_23302_));
 sky130_as_sc_hs__nand3_2 _29816_ (.A(net228),
    .B(_23303_),
    .C(_23304_),
    .Y(_23305_));
 sky130_as_sc_hs__nand3_2 _29819_ (.A(net367),
    .B(_23306_),
    .C(_23307_),
    .Y(_23308_));
 sky130_as_sc_hs__nand3_2 _29820_ (.A(net238),
    .B(_23305_),
    .C(_23308_),
    .Y(_23309_));
 sky130_as_sc_hs__nand3_2 _29823_ (.A(net228),
    .B(_23310_),
    .C(_23311_),
    .Y(_23312_));
 sky130_as_sc_hs__nand3_2 _29826_ (.A(net367),
    .B(_23313_),
    .C(_23314_),
    .Y(_23315_));
 sky130_as_sc_hs__nand3_2 _29827_ (.A(net349),
    .B(_23312_),
    .C(_23315_),
    .Y(_23316_));
 sky130_as_sc_hs__nand3_2 _29830_ (.A(net226),
    .B(_23317_),
    .C(_23318_),
    .Y(_23319_));
 sky130_as_sc_hs__nand3_2 _29833_ (.A(net364),
    .B(_23320_),
    .C(_23321_),
    .Y(_23322_));
 sky130_as_sc_hs__nand3_2 _29834_ (.A(net237),
    .B(_23319_),
    .C(_23322_),
    .Y(_23323_));
 sky130_as_sc_hs__nand3_2 _29837_ (.A(net364),
    .B(_23324_),
    .C(_23325_),
    .Y(_23326_));
 sky130_as_sc_hs__nand3_2 _29840_ (.A(net228),
    .B(_23327_),
    .C(_23328_),
    .Y(_23329_));
 sky130_as_sc_hs__nand3_2 _29841_ (.A(net349),
    .B(_23326_),
    .C(_23329_),
    .Y(_23330_));
 sky130_as_sc_hs__nand3_2 _29842_ (.A(net244),
    .B(_23323_),
    .C(_23330_),
    .Y(_23331_));
 sky130_as_sc_hs__nand3_2 _29843_ (.A(net339),
    .B(_23309_),
    .C(_23316_),
    .Y(_23332_));
 sky130_as_sc_hs__nand3_2 _29844_ (.A(net245),
    .B(_23331_),
    .C(_23332_),
    .Y(_23333_));
 sky130_as_sc_hs__nand3_2 _29848_ (.A(net213),
    .B(_23335_),
    .C(_23336_),
    .Y(_23337_));
 sky130_as_sc_hs__nand3_2 _29851_ (.A(net353),
    .B(_23338_),
    .C(_23339_),
    .Y(_23340_));
 sky130_as_sc_hs__nand3_2 _29852_ (.A(net231),
    .B(_23337_),
    .C(_23340_),
    .Y(_23341_));
 sky130_as_sc_hs__nand3_2 _29855_ (.A(net213),
    .B(_23342_),
    .C(_23343_),
    .Y(_23344_));
 sky130_as_sc_hs__nand3_2 _29858_ (.A(net352),
    .B(_23345_),
    .C(_23346_),
    .Y(_23347_));
 sky130_as_sc_hs__nand3_2 _29859_ (.A(net342),
    .B(_23344_),
    .C(_23347_),
    .Y(_23348_));
 sky130_as_sc_hs__nand3_2 _29862_ (.A(net221),
    .B(_23349_),
    .C(_23350_),
    .Y(_23351_));
 sky130_as_sc_hs__nand3_2 _29865_ (.A(net360),
    .B(_23352_),
    .C(_23353_),
    .Y(_23354_));
 sky130_as_sc_hs__nand3_2 _29866_ (.A(net236),
    .B(_23351_),
    .C(_23354_),
    .Y(_23355_));
 sky130_as_sc_hs__nand3_2 _29869_ (.A(net360),
    .B(_23356_),
    .C(_23357_),
    .Y(_23358_));
 sky130_as_sc_hs__nand3_2 _29872_ (.A(net221),
    .B(_23359_),
    .C(_23360_),
    .Y(_23361_));
 sky130_as_sc_hs__nand3_2 _29873_ (.A(net347),
    .B(_23358_),
    .C(_23361_),
    .Y(_23362_));
 sky130_as_sc_hs__nand3_2 _29874_ (.A(net242),
    .B(_23355_),
    .C(_23362_),
    .Y(_23363_));
 sky130_as_sc_hs__nand3_2 _29875_ (.A(net337),
    .B(_23341_),
    .C(_23348_),
    .Y(_23364_));
 sky130_as_sc_hs__nand3_2 _29876_ (.A(net335),
    .B(_23363_),
    .C(_23364_),
    .Y(_23365_));
 sky130_as_sc_hs__nand3_2 _29879_ (.A(net213),
    .B(_23366_),
    .C(_23367_),
    .Y(_23368_));
 sky130_as_sc_hs__nand3_2 _29882_ (.A(net352),
    .B(_23369_),
    .C(_23370_),
    .Y(_23371_));
 sky130_as_sc_hs__nand3_2 _29883_ (.A(net231),
    .B(_23368_),
    .C(_23371_),
    .Y(_23372_));
 sky130_as_sc_hs__nand3_2 _29886_ (.A(net221),
    .B(_23373_),
    .C(_23374_),
    .Y(_23375_));
 sky130_as_sc_hs__nand3_2 _29889_ (.A(net360),
    .B(_23376_),
    .C(_23377_),
    .Y(_23378_));
 sky130_as_sc_hs__nand3_2 _29890_ (.A(net347),
    .B(_23375_),
    .C(_23378_),
    .Y(_23379_));
 sky130_as_sc_hs__nand3_2 _29893_ (.A(net221),
    .B(_23380_),
    .C(_23381_),
    .Y(_23382_));
 sky130_as_sc_hs__nand3_2 _29896_ (.A(net360),
    .B(_23383_),
    .C(_23384_),
    .Y(_23385_));
 sky130_as_sc_hs__nand3_2 _29897_ (.A(net236),
    .B(_23382_),
    .C(_23385_),
    .Y(_23386_));
 sky130_as_sc_hs__nand3_2 _29900_ (.A(net360),
    .B(_23387_),
    .C(_23388_),
    .Y(_23389_));
 sky130_as_sc_hs__nand3_2 _29903_ (.A(net221),
    .B(_23390_),
    .C(_23391_),
    .Y(_23392_));
 sky130_as_sc_hs__nand3_2 _29904_ (.A(net347),
    .B(_23389_),
    .C(_23392_),
    .Y(_23393_));
 sky130_as_sc_hs__nand3_2 _29905_ (.A(net242),
    .B(_23386_),
    .C(_23393_),
    .Y(_23394_));
 sky130_as_sc_hs__nand3_2 _29906_ (.A(net337),
    .B(_23372_),
    .C(_23379_),
    .Y(_23395_));
 sky130_as_sc_hs__nand3_2 _29907_ (.A(net246),
    .B(_23394_),
    .C(_23395_),
    .Y(_23396_));
 sky130_as_sc_hs__and2_2 _29908_ (.A(_23365_),
    .B(_23396_),
    .Y(_23397_));
 sky130_as_sc_hs__inv_2 _29909_ (.Y(_23398_),
    .A(_23397_));
 sky130_as_sc_hs__nand3_2 _29912_ (.A(net212),
    .B(_23399_),
    .C(_23400_),
    .Y(_23401_));
 sky130_as_sc_hs__nand3_2 _29915_ (.A(net352),
    .B(_23402_),
    .C(_23403_),
    .Y(_23404_));
 sky130_as_sc_hs__nand3_2 _29916_ (.A(net231),
    .B(_23401_),
    .C(_23404_),
    .Y(_23405_));
 sky130_as_sc_hs__nand3_2 _29919_ (.A(net212),
    .B(_23406_),
    .C(_23407_),
    .Y(_23408_));
 sky130_as_sc_hs__nand3_2 _29922_ (.A(net352),
    .B(_23409_),
    .C(_23410_),
    .Y(_23411_));
 sky130_as_sc_hs__nand3_2 _29923_ (.A(net342),
    .B(_23408_),
    .C(_23411_),
    .Y(_23412_));
 sky130_as_sc_hs__nand3_2 _29926_ (.A(net212),
    .B(_23413_),
    .C(_23414_),
    .Y(_23415_));
 sky130_as_sc_hs__nand3_2 _29929_ (.A(net352),
    .B(_23416_),
    .C(_23417_),
    .Y(_23418_));
 sky130_as_sc_hs__nand3_2 _29930_ (.A(net231),
    .B(_23415_),
    .C(_23418_),
    .Y(_23419_));
 sky130_as_sc_hs__nand3_2 _29933_ (.A(net352),
    .B(_23420_),
    .C(_23421_),
    .Y(_23422_));
 sky130_as_sc_hs__nand3_2 _29936_ (.A(net213),
    .B(_23423_),
    .C(_23424_),
    .Y(_23425_));
 sky130_as_sc_hs__nand3_2 _29937_ (.A(net342),
    .B(_23422_),
    .C(_23425_),
    .Y(_23426_));
 sky130_as_sc_hs__nand3_2 _29938_ (.A(net240),
    .B(_23419_),
    .C(_23426_),
    .Y(_23427_));
 sky130_as_sc_hs__nand3_2 _29939_ (.A(net337),
    .B(_23405_),
    .C(_23412_),
    .Y(_23428_));
 sky130_as_sc_hs__nand3_2 _29940_ (.A(net336),
    .B(_23427_),
    .C(_23428_),
    .Y(_23429_));
 sky130_as_sc_hs__nand3_2 _29943_ (.A(net212),
    .B(_23430_),
    .C(_23431_),
    .Y(_23432_));
 sky130_as_sc_hs__nand3_2 _29946_ (.A(net352),
    .B(_23433_),
    .C(_23434_),
    .Y(_23435_));
 sky130_as_sc_hs__nand3_2 _29947_ (.A(net231),
    .B(_23432_),
    .C(_23435_),
    .Y(_23436_));
 sky130_as_sc_hs__nand3_2 _29950_ (.A(net212),
    .B(_23437_),
    .C(_23438_),
    .Y(_23439_));
 sky130_as_sc_hs__nand3_2 _29953_ (.A(net352),
    .B(_23440_),
    .C(_23441_),
    .Y(_23442_));
 sky130_as_sc_hs__nand3_2 _29954_ (.A(net342),
    .B(_23439_),
    .C(_23442_),
    .Y(_23443_));
 sky130_as_sc_hs__nand3_2 _29957_ (.A(net212),
    .B(_23444_),
    .C(_23445_),
    .Y(_23446_));
 sky130_as_sc_hs__nand3_2 _29960_ (.A(net352),
    .B(_23447_),
    .C(_23448_),
    .Y(_23449_));
 sky130_as_sc_hs__nand3_2 _29961_ (.A(net231),
    .B(_23446_),
    .C(_23449_),
    .Y(_23450_));
 sky130_as_sc_hs__nand3_2 _29964_ (.A(net352),
    .B(_23451_),
    .C(_23452_),
    .Y(_23453_));
 sky130_as_sc_hs__nand3_2 _29967_ (.A(net212),
    .B(_23454_),
    .C(_23455_),
    .Y(_23456_));
 sky130_as_sc_hs__nand3_2 _29968_ (.A(net342),
    .B(_23453_),
    .C(_23456_),
    .Y(_23457_));
 sky130_as_sc_hs__nand3_2 _29969_ (.A(net240),
    .B(_23450_),
    .C(_23457_),
    .Y(_23458_));
 sky130_as_sc_hs__nand3_2 _29970_ (.A(net337),
    .B(_23436_),
    .C(_23443_),
    .Y(_23459_));
 sky130_as_sc_hs__nand3_2 _29971_ (.A(net246),
    .B(_23458_),
    .C(_23459_),
    .Y(_23460_));
 sky130_as_sc_hs__and2_2 _29972_ (.A(_23429_),
    .B(_23460_),
    .Y(_23461_));
 sky130_as_sc_hs__inv_2 _29973_ (.Y(_23462_),
    .A(_23461_));
 sky130_as_sc_hs__nand3_2 _29976_ (.A(net213),
    .B(_23463_),
    .C(_23464_),
    .Y(_23465_));
 sky130_as_sc_hs__nand3_2 _29979_ (.A(net353),
    .B(_23466_),
    .C(_23467_),
    .Y(_23468_));
 sky130_as_sc_hs__nand3_2 _29980_ (.A(net231),
    .B(_23465_),
    .C(_23468_),
    .Y(_23469_));
 sky130_as_sc_hs__nand3_2 _29983_ (.A(net213),
    .B(_23470_),
    .C(_23471_),
    .Y(_23472_));
 sky130_as_sc_hs__nand3_2 _29986_ (.A(net353),
    .B(_23473_),
    .C(_23474_),
    .Y(_23475_));
 sky130_as_sc_hs__nand3_2 _29987_ (.A(net342),
    .B(_23472_),
    .C(_23475_),
    .Y(_23476_));
 sky130_as_sc_hs__nand3_2 _29990_ (.A(net213),
    .B(_23477_),
    .C(_23478_),
    .Y(_23479_));
 sky130_as_sc_hs__nand3_2 _29993_ (.A(net353),
    .B(_23480_),
    .C(_23481_),
    .Y(_23482_));
 sky130_as_sc_hs__nand3_2 _29994_ (.A(net231),
    .B(_23479_),
    .C(_23482_),
    .Y(_23483_));
 sky130_as_sc_hs__nand3_2 _29997_ (.A(net353),
    .B(_23484_),
    .C(_23485_),
    .Y(_23486_));
 sky130_as_sc_hs__nand3_2 _30000_ (.A(net213),
    .B(_23487_),
    .C(_23488_),
    .Y(_23489_));
 sky130_as_sc_hs__nand3_2 _30001_ (.A(net342),
    .B(_23486_),
    .C(_23489_),
    .Y(_23490_));
 sky130_as_sc_hs__nand3_2 _30002_ (.A(net240),
    .B(_23483_),
    .C(_23490_),
    .Y(_23491_));
 sky130_as_sc_hs__nand3_2 _30003_ (.A(net337),
    .B(_23469_),
    .C(_23476_),
    .Y(_23492_));
 sky130_as_sc_hs__nand3_2 _30004_ (.A(net336),
    .B(_23491_),
    .C(_23492_),
    .Y(_23493_));
 sky130_as_sc_hs__nand3_2 _30007_ (.A(net214),
    .B(_23494_),
    .C(_23495_),
    .Y(_23496_));
 sky130_as_sc_hs__nand3_2 _30010_ (.A(net353),
    .B(_23497_),
    .C(_23498_),
    .Y(_23499_));
 sky130_as_sc_hs__nand3_2 _30011_ (.A(net231),
    .B(_23496_),
    .C(_23499_),
    .Y(_23500_));
 sky130_as_sc_hs__nand3_2 _30014_ (.A(net214),
    .B(_23501_),
    .C(_23502_),
    .Y(_23503_));
 sky130_as_sc_hs__nand3_2 _30017_ (.A(net353),
    .B(_23504_),
    .C(_23505_),
    .Y(_23506_));
 sky130_as_sc_hs__nand3_2 _30018_ (.A(net342),
    .B(_23503_),
    .C(_23506_),
    .Y(_23507_));
 sky130_as_sc_hs__nand3_2 _30021_ (.A(net213),
    .B(_23508_),
    .C(_23509_),
    .Y(_23510_));
 sky130_as_sc_hs__nand3_2 _30024_ (.A(net353),
    .B(_23511_),
    .C(_23512_),
    .Y(_23513_));
 sky130_as_sc_hs__nand3_2 _30025_ (.A(net231),
    .B(_23510_),
    .C(_23513_),
    .Y(_23514_));
 sky130_as_sc_hs__nand3_2 _30028_ (.A(net354),
    .B(_23515_),
    .C(_23516_),
    .Y(_23517_));
 sky130_as_sc_hs__nand3_2 _30031_ (.A(net213),
    .B(_23518_),
    .C(_23519_),
    .Y(_23520_));
 sky130_as_sc_hs__nand3_2 _30032_ (.A(net342),
    .B(_23517_),
    .C(_23520_),
    .Y(_23521_));
 sky130_as_sc_hs__nand3_2 _30033_ (.A(net240),
    .B(_23514_),
    .C(_23521_),
    .Y(_23522_));
 sky130_as_sc_hs__nand3_2 _30034_ (.A(net337),
    .B(_23500_),
    .C(_23507_),
    .Y(_23523_));
 sky130_as_sc_hs__nand3_2 _30035_ (.A(net246),
    .B(_23522_),
    .C(_23523_),
    .Y(_23524_));
 sky130_as_sc_hs__and2_2 _30036_ (.A(_23493_),
    .B(_23524_),
    .Y(_23525_));
 sky130_as_sc_hs__nand3_2 _30037_ (.A(_23397_),
    .B(_23461_),
    .C(_23525_),
    .Y(_23526_));
 sky130_as_sc_hs__nor2_2 _30038_ (.A(_23334_),
    .B(_23526_),
    .Y(_23527_));
 sky130_as_sc_hs__nand3_2 _30039_ (.A(_23014_),
    .B(_23270_),
    .C(_23527_),
    .Y(_23528_));
 sky130_as_sc_hs__nor2_2 _30040_ (.A(_21723_),
    .B(_23528_),
    .Y(_23529_));
 sky130_as_sc_hs__and2_2 _30041_ (.A(_21723_),
    .B(_23528_),
    .Y(_23530_));
 sky130_as_sc_hs__or2_2 _30042_ (.A(_23529_),
    .B(_23530_),
    .Y(_23531_));
 sky130_as_sc_hs__or2_2 _30044_ (.A(_21659_),
    .B(_21723_),
    .Y(_23533_));
 sky130_as_sc_hs__and2_2 _30045_ (.A(_23532_),
    .B(_23533_),
    .Y(_23534_));
 sky130_as_sc_hs__and2_2 _30046_ (.A(net114),
    .B(net123),
    .Y(_23535_));
 sky130_as_sc_hs__nand3_2 _30049_ (.A(net177),
    .B(_23536_),
    .C(_23537_),
    .Y(_23538_));
 sky130_as_sc_hs__nand3_2 _30052_ (.A(net274),
    .B(_23539_),
    .C(_23540_),
    .Y(_23541_));
 sky130_as_sc_hs__nand3_2 _30053_ (.A(net159),
    .B(_23538_),
    .C(_23541_),
    .Y(_23542_));
 sky130_as_sc_hs__nand3_2 _30056_ (.A(net178),
    .B(_23543_),
    .C(_23544_),
    .Y(_23545_));
 sky130_as_sc_hs__nand3_2 _30059_ (.A(net273),
    .B(_23546_),
    .C(_23547_),
    .Y(_23548_));
 sky130_as_sc_hs__nand3_2 _30060_ (.A(net259),
    .B(_23545_),
    .C(_23548_),
    .Y(_23549_));
 sky130_as_sc_hs__nand3_2 _30063_ (.A(net178),
    .B(_23550_),
    .C(_23551_),
    .Y(_23552_));
 sky130_as_sc_hs__nand3_2 _30066_ (.A(net274),
    .B(_23553_),
    .C(_23554_),
    .Y(_23555_));
 sky130_as_sc_hs__nand3_2 _30067_ (.A(net159),
    .B(_23552_),
    .C(_23555_),
    .Y(_23556_));
 sky130_as_sc_hs__nand3_2 _30070_ (.A(net274),
    .B(_23557_),
    .C(_23558_),
    .Y(_23559_));
 sky130_as_sc_hs__nand3_2 _30073_ (.A(net178),
    .B(_23560_),
    .C(_23561_),
    .Y(_23562_));
 sky130_as_sc_hs__nand3_2 _30074_ (.A(net259),
    .B(_23559_),
    .C(_23562_),
    .Y(_23563_));
 sky130_as_sc_hs__nand3_2 _30075_ (.A(net153),
    .B(_23556_),
    .C(_23563_),
    .Y(_23564_));
 sky130_as_sc_hs__nand3_2 _30076_ (.A(net249),
    .B(_23542_),
    .C(_23549_),
    .Y(_23565_));
 sky130_as_sc_hs__nand3_2 _30077_ (.A(net248),
    .B(_23564_),
    .C(_23565_),
    .Y(_23566_));
 sky130_as_sc_hs__nand3_2 _30080_ (.A(net177),
    .B(_23567_),
    .C(_23568_),
    .Y(_23569_));
 sky130_as_sc_hs__nand3_2 _30083_ (.A(net273),
    .B(_23570_),
    .C(_23571_),
    .Y(_23572_));
 sky130_as_sc_hs__nand3_2 _30084_ (.A(net160),
    .B(_23569_),
    .C(_23572_),
    .Y(_23573_));
 sky130_as_sc_hs__nand3_2 _30087_ (.A(net177),
    .B(_23574_),
    .C(_23575_),
    .Y(_23576_));
 sky130_as_sc_hs__nand3_2 _30090_ (.A(net273),
    .B(_23577_),
    .C(_23578_),
    .Y(_23579_));
 sky130_as_sc_hs__nand3_2 _30091_ (.A(net259),
    .B(_23576_),
    .C(_23579_),
    .Y(_23580_));
 sky130_as_sc_hs__nand3_2 _30094_ (.A(net177),
    .B(_23581_),
    .C(_23582_),
    .Y(_23583_));
 sky130_as_sc_hs__nand3_2 _30097_ (.A(net273),
    .B(_23584_),
    .C(_23585_),
    .Y(_23586_));
 sky130_as_sc_hs__nand3_2 _30098_ (.A(net159),
    .B(_23583_),
    .C(_23586_),
    .Y(_23587_));
 sky130_as_sc_hs__nand3_2 _30101_ (.A(net273),
    .B(_23588_),
    .C(_23589_),
    .Y(_23590_));
 sky130_as_sc_hs__nand3_2 _30104_ (.A(net177),
    .B(_23591_),
    .C(_23592_),
    .Y(_23593_));
 sky130_as_sc_hs__nand3_2 _30105_ (.A(net258),
    .B(_23590_),
    .C(_23593_),
    .Y(_23594_));
 sky130_as_sc_hs__nand3_2 _30106_ (.A(net152),
    .B(_23587_),
    .C(_23594_),
    .Y(_23595_));
 sky130_as_sc_hs__nand3_2 _30107_ (.A(net249),
    .B(_23573_),
    .C(_23580_),
    .Y(_23596_));
 sky130_as_sc_hs__nand3_2 _30108_ (.A(net150),
    .B(_23595_),
    .C(_23596_),
    .Y(_23597_));
 sky130_as_sc_hs__and2_2 _30110_ (.A(_19486_),
    .B(\tholin_riscv.Jimm[12] ),
    .Y(_23599_));
 sky130_as_sc_hs__nor2_2 _30112_ (.A(net411),
    .B(_23600_),
    .Y(_23601_));
 sky130_as_sc_hs__or2_2 _30113_ (.A(net411),
    .B(_23600_),
    .Y(_23602_));
 sky130_as_sc_hs__nor2_2 _30114_ (.A(\tholin_riscv.Jimm[13] ),
    .B(\tholin_riscv.Jimm[12] ),
    .Y(_23603_));
 sky130_as_sc_hs__or2_2 _30115_ (.A(\tholin_riscv.Jimm[13] ),
    .B(\tholin_riscv.Jimm[12] ),
    .Y(_23604_));
 sky130_as_sc_hs__or2_2 _30116_ (.A(net411),
    .B(_23604_),
    .Y(_23605_));
 sky130_as_sc_hs__nor2_2 _30117_ (.A(net411),
    .B(\tholin_riscv.Jimm[13] ),
    .Y(_23606_));
 sky130_as_sc_hs__and2_2 _30118_ (.A(_23598_),
    .B(_23606_),
    .Y(_23607_));
 sky130_as_sc_hs__nand3_2 _30121_ (.A(_20826_),
    .B(_20932_),
    .C(_21037_),
    .Y(_23610_));
 sky130_as_sc_hs__nor2_2 _30122_ (.A(_21140_),
    .B(_23610_),
    .Y(_23611_));
 sky130_as_sc_hs__nand3_2 _30124_ (.A(_21242_),
    .B(_21344_),
    .C(_23611_),
    .Y(_23613_));
 sky130_as_sc_hs__nor2_2 _30125_ (.A(_21343_),
    .B(_21440_),
    .Y(_23614_));
 sky130_as_sc_hs__and2_2 _30126_ (.A(_21534_),
    .B(_23614_),
    .Y(_23615_));
 sky130_as_sc_hs__nand3_2 _30127_ (.A(_21242_),
    .B(_23611_),
    .C(_23615_),
    .Y(_23616_));
 sky130_as_sc_hs__nor2_2 _30128_ (.A(_20106_),
    .B(_23616_),
    .Y(_23617_));
 sky130_as_sc_hs__and2_2 _30129_ (.A(_20191_),
    .B(_23617_),
    .Y(_23618_));
 sky130_as_sc_hs__nand3_2 _30130_ (.A(_20191_),
    .B(_20277_),
    .C(_23617_),
    .Y(_23619_));
 sky130_as_sc_hs__or2_2 _30131_ (.A(_20277_),
    .B(_23618_),
    .Y(_23620_));
 sky130_as_sc_hs__and2_2 _30135_ (.A(_23622_),
    .B(_23623_),
    .Y(_23624_));
 sky130_as_sc_hs__and2_2 _30140_ (.A(_23627_),
    .B(_23628_),
    .Y(_23629_));
 sky130_as_sc_hs__and2_2 _30141_ (.A(net482),
    .B(net480),
    .Y(_23630_));
 sky130_as_sc_hs__or2_2 _30143_ (.A(_21440_),
    .B(_23613_),
    .Y(_23632_));
 sky130_as_sc_hs__and2_2 _30145_ (.A(_23632_),
    .B(_23633_),
    .Y(_23634_));
 sky130_as_sc_hs__nand3_2 _30149_ (.A(_23014_),
    .B(_23204_),
    .C(_23268_),
    .Y(_23638_));
 sky130_as_sc_hs__and2_2 _30154_ (.A(_23641_),
    .B(_23642_),
    .Y(_23643_));
 sky130_as_sc_hs__and2_2 _30155_ (.A(_23636_),
    .B(net478),
    .Y(_23644_));
 sky130_as_sc_hs__or2_2 _30157_ (.A(_22947_),
    .B(_23011_),
    .Y(_23646_));
 sky130_as_sc_hs__and2_2 _30161_ (.A(_23648_),
    .B(_23649_),
    .Y(_23650_));
 sky130_as_sc_hs__and2_2 _30162_ (.A(net483),
    .B(net477),
    .Y(_23651_));
 sky130_as_sc_hs__or2_2 _30163_ (.A(_23078_),
    .B(_23638_),
    .Y(_23652_));
 sky130_as_sc_hs__and2_2 _30168_ (.A(_23655_),
    .B(_23656_),
    .Y(_23657_));
 sky130_as_sc_hs__and2_2 _30169_ (.A(_23636_),
    .B(net475),
    .Y(_23658_));
 sky130_as_sc_hs__or2_2 _30171_ (.A(_23651_),
    .B(_23658_),
    .Y(_23660_));
 sky130_as_sc_hs__or2_2 _30173_ (.A(_23645_),
    .B(_23661_),
    .Y(_23662_));
 sky130_as_sc_hs__and2_2 _30175_ (.A(_23662_),
    .B(_23663_),
    .Y(_23664_));
 sky130_as_sc_hs__or2_2 _30177_ (.A(_23535_),
    .B(_23664_),
    .Y(_23666_));
 sky130_as_sc_hs__and2_2 _30178_ (.A(_23665_),
    .B(_23666_),
    .Y(_23667_));
 sky130_as_sc_hs__or2_2 _30179_ (.A(_23630_),
    .B(_23644_),
    .Y(_23668_));
 sky130_as_sc_hs__or2_2 _30181_ (.A(_21659_),
    .B(_22945_),
    .Y(_23670_));
 sky130_as_sc_hs__or2_2 _30182_ (.A(_22882_),
    .B(_22945_),
    .Y(_23671_));
 sky130_as_sc_hs__and2_2 _30183_ (.A(_22946_),
    .B(_23671_),
    .Y(_23672_));
 sky130_as_sc_hs__and2_2 _30186_ (.A(net482),
    .B(_23674_),
    .Y(_23675_));
 sky130_as_sc_hs__or2_2 _30187_ (.A(_23014_),
    .B(_23268_),
    .Y(_23676_));
 sky130_as_sc_hs__and2_2 _30191_ (.A(_23678_),
    .B(_23679_),
    .Y(_23680_));
 sky130_as_sc_hs__and2_2 _30192_ (.A(_23636_),
    .B(net473),
    .Y(_23681_));
 sky130_as_sc_hs__or2_2 _30194_ (.A(_23669_),
    .B(_23682_),
    .Y(_23683_));
 sky130_as_sc_hs__nand3_2 _30195_ (.A(_23014_),
    .B(_23270_),
    .C(_23525_),
    .Y(_23684_));
 sky130_as_sc_hs__or2_2 _30196_ (.A(_23462_),
    .B(_23684_),
    .Y(_23685_));
 sky130_as_sc_hs__or2_2 _30197_ (.A(_23398_),
    .B(_23685_),
    .Y(_23686_));
 sky130_as_sc_hs__or2_2 _30201_ (.A(_21659_),
    .B(_23334_),
    .Y(_23690_));
 sky130_as_sc_hs__and2_2 _30202_ (.A(_23689_),
    .B(_23690_),
    .Y(_23691_));
 sky130_as_sc_hs__and2_2 _30203_ (.A(net115),
    .B(net121),
    .Y(_23692_));
 sky130_as_sc_hs__and2_2 _30205_ (.A(_23683_),
    .B(_23693_),
    .Y(_23694_));
 sky130_as_sc_hs__and2_2 _30210_ (.A(_20106_),
    .B(_23616_),
    .Y(_23699_));
 sky130_as_sc_hs__nor2_2 _30211_ (.A(_23617_),
    .B(_23699_),
    .Y(_23700_));
 sky130_as_sc_hs__and2_2 _30214_ (.A(net473),
    .B(_23702_),
    .Y(_23703_));
 sky130_as_sc_hs__or2_2 _30215_ (.A(_23667_),
    .B(_23696_),
    .Y(_23704_));
 sky130_as_sc_hs__and2_2 _30216_ (.A(_23697_),
    .B(_23704_),
    .Y(_23705_));
 sky130_as_sc_hs__or2_2 _30220_ (.A(_22171_),
    .B(_22235_),
    .Y(_23709_));
 sky130_as_sc_hs__or2_2 _30222_ (.A(_21660_),
    .B(_23710_),
    .Y(_23711_));
 sky130_as_sc_hs__or2_2 _30225_ (.A(net305),
    .B(\tholin_riscv.regs[24][20] ),
    .Y(_23714_));
 sky130_as_sc_hs__nand3_2 _30226_ (.A(net172),
    .B(_23713_),
    .C(_23714_),
    .Y(_23715_));
 sky130_as_sc_hs__or2_2 _30228_ (.A(net305),
    .B(\tholin_riscv.regs[26][20] ),
    .Y(_23717_));
 sky130_as_sc_hs__nand3_2 _30229_ (.A(net268),
    .B(_23716_),
    .C(_23717_),
    .Y(_23718_));
 sky130_as_sc_hs__nand3_2 _30230_ (.A(net162),
    .B(_23715_),
    .C(_23718_),
    .Y(_23719_));
 sky130_as_sc_hs__or2_2 _30232_ (.A(net324),
    .B(\tholin_riscv.regs[28][20] ),
    .Y(_23721_));
 sky130_as_sc_hs__nand3_2 _30233_ (.A(net180),
    .B(_23720_),
    .C(_23721_),
    .Y(_23722_));
 sky130_as_sc_hs__or2_2 _30235_ (.A(net326),
    .B(\tholin_riscv.regs[30][20] ),
    .Y(_23724_));
 sky130_as_sc_hs__nand3_2 _30236_ (.A(net276),
    .B(_23723_),
    .C(_23724_),
    .Y(_23725_));
 sky130_as_sc_hs__nand3_2 _30237_ (.A(net260),
    .B(_23722_),
    .C(_23725_),
    .Y(_23726_));
 sky130_as_sc_hs__or2_2 _30239_ (.A(net305),
    .B(\tholin_riscv.regs[16][20] ),
    .Y(_23728_));
 sky130_as_sc_hs__nand3_2 _30240_ (.A(net171),
    .B(_23727_),
    .C(_23728_),
    .Y(_23729_));
 sky130_as_sc_hs__or2_2 _30242_ (.A(net305),
    .B(\tholin_riscv.regs[18][20] ),
    .Y(_23731_));
 sky130_as_sc_hs__nand3_2 _30243_ (.A(net269),
    .B(_23730_),
    .C(_23731_),
    .Y(_23732_));
 sky130_as_sc_hs__nand3_2 _30244_ (.A(net162),
    .B(_23729_),
    .C(_23732_),
    .Y(_23733_));
 sky130_as_sc_hs__or2_2 _30246_ (.A(net305),
    .B(\tholin_riscv.regs[22][20] ),
    .Y(_23735_));
 sky130_as_sc_hs__nand3_2 _30247_ (.A(net268),
    .B(_23734_),
    .C(_23735_),
    .Y(_23736_));
 sky130_as_sc_hs__or2_2 _30249_ (.A(net305),
    .B(\tholin_riscv.regs[20][20] ),
    .Y(_23738_));
 sky130_as_sc_hs__nand3_2 _30250_ (.A(net171),
    .B(_23737_),
    .C(_23738_),
    .Y(_23739_));
 sky130_as_sc_hs__nand3_2 _30251_ (.A(net254),
    .B(_23736_),
    .C(_23739_),
    .Y(_23740_));
 sky130_as_sc_hs__nand3_2 _30252_ (.A(net156),
    .B(_23733_),
    .C(_23740_),
    .Y(_23741_));
 sky130_as_sc_hs__nand3_2 _30253_ (.A(net251),
    .B(_23719_),
    .C(_23726_),
    .Y(_23742_));
 sky130_as_sc_hs__nand3_2 _30254_ (.A(net247),
    .B(_23741_),
    .C(_23742_),
    .Y(_23743_));
 sky130_as_sc_hs__or2_2 _30256_ (.A(net303),
    .B(\tholin_riscv.regs[8][20] ),
    .Y(_23745_));
 sky130_as_sc_hs__nand3_2 _30257_ (.A(net171),
    .B(_23744_),
    .C(_23745_),
    .Y(_23746_));
 sky130_as_sc_hs__or2_2 _30259_ (.A(net303),
    .B(\tholin_riscv.regs[10][20] ),
    .Y(_23748_));
 sky130_as_sc_hs__nand3_2 _30260_ (.A(net268),
    .B(_23747_),
    .C(_23748_),
    .Y(_23749_));
 sky130_as_sc_hs__nand3_2 _30261_ (.A(net165),
    .B(_23746_),
    .C(_23749_),
    .Y(_23750_));
 sky130_as_sc_hs__or2_2 _30263_ (.A(net305),
    .B(\tholin_riscv.regs[12][20] ),
    .Y(_23752_));
 sky130_as_sc_hs__nand3_2 _30264_ (.A(net171),
    .B(_23751_),
    .C(_23752_),
    .Y(_23753_));
 sky130_as_sc_hs__or2_2 _30266_ (.A(net306),
    .B(\tholin_riscv.regs[14][20] ),
    .Y(_23755_));
 sky130_as_sc_hs__nand3_2 _30267_ (.A(net268),
    .B(_23754_),
    .C(_23755_),
    .Y(_23756_));
 sky130_as_sc_hs__nand3_2 _30268_ (.A(_00002_),
    .B(_23753_),
    .C(_23756_),
    .Y(_23757_));
 sky130_as_sc_hs__or2_2 _30270_ (.A(net305),
    .B(\tholin_riscv.regs[0][20] ),
    .Y(_23759_));
 sky130_as_sc_hs__nand3_2 _30271_ (.A(net171),
    .B(_23758_),
    .C(_23759_),
    .Y(_23760_));
 sky130_as_sc_hs__or2_2 _30273_ (.A(net303),
    .B(\tholin_riscv.regs[2][20] ),
    .Y(_23762_));
 sky130_as_sc_hs__nand3_2 _30274_ (.A(net268),
    .B(_23761_),
    .C(_23762_),
    .Y(_23763_));
 sky130_as_sc_hs__nand3_2 _30275_ (.A(net165),
    .B(_23760_),
    .C(_23763_),
    .Y(_23764_));
 sky130_as_sc_hs__or2_2 _30277_ (.A(net305),
    .B(\tholin_riscv.regs[6][20] ),
    .Y(_23766_));
 sky130_as_sc_hs__nand3_2 _30278_ (.A(net268),
    .B(_23765_),
    .C(_23766_),
    .Y(_23767_));
 sky130_as_sc_hs__or2_2 _30280_ (.A(net305),
    .B(\tholin_riscv.regs[4][20] ),
    .Y(_23769_));
 sky130_as_sc_hs__nand3_2 _30281_ (.A(net171),
    .B(_23768_),
    .C(_23769_),
    .Y(_23770_));
 sky130_as_sc_hs__nand3_2 _30282_ (.A(net255),
    .B(_23767_),
    .C(_23770_),
    .Y(_23771_));
 sky130_as_sc_hs__nand3_2 _30283_ (.A(net156),
    .B(_23764_),
    .C(_23771_),
    .Y(_23772_));
 sky130_as_sc_hs__nand3_2 _30284_ (.A(net253),
    .B(_23750_),
    .C(_23757_),
    .Y(_23773_));
 sky130_as_sc_hs__nand3_2 _30285_ (.A(net151),
    .B(_23772_),
    .C(_23773_),
    .Y(_23774_));
 sky130_as_sc_hs__inv_2 _30287_ (.Y(_23776_),
    .A(_23775_));
 sky130_as_sc_hs__or2_2 _30289_ (.A(net305),
    .B(\tholin_riscv.regs[24][19] ),
    .Y(_23778_));
 sky130_as_sc_hs__nand3_2 _30290_ (.A(net171),
    .B(_23777_),
    .C(_23778_),
    .Y(_23779_));
 sky130_as_sc_hs__or2_2 _30292_ (.A(net305),
    .B(\tholin_riscv.regs[26][19] ),
    .Y(_23781_));
 sky130_as_sc_hs__nand3_2 _30293_ (.A(net268),
    .B(_23780_),
    .C(_23781_),
    .Y(_23782_));
 sky130_as_sc_hs__nand3_2 _30294_ (.A(net162),
    .B(_23779_),
    .C(_23782_),
    .Y(_23783_));
 sky130_as_sc_hs__or2_2 _30296_ (.A(net306),
    .B(\tholin_riscv.regs[28][19] ),
    .Y(_23785_));
 sky130_as_sc_hs__nand3_2 _30297_ (.A(net172),
    .B(_23784_),
    .C(_23785_),
    .Y(_23786_));
 sky130_as_sc_hs__or2_2 _30299_ (.A(net306),
    .B(\tholin_riscv.regs[30][19] ),
    .Y(_23788_));
 sky130_as_sc_hs__nand3_2 _30300_ (.A(net269),
    .B(_23787_),
    .C(_23788_),
    .Y(_23789_));
 sky130_as_sc_hs__nand3_2 _30301_ (.A(net254),
    .B(_23786_),
    .C(_23789_),
    .Y(_23790_));
 sky130_as_sc_hs__or2_2 _30303_ (.A(net305),
    .B(\tholin_riscv.regs[16][19] ),
    .Y(_23792_));
 sky130_as_sc_hs__nand3_2 _30304_ (.A(net171),
    .B(_23791_),
    .C(_23792_),
    .Y(_23793_));
 sky130_as_sc_hs__or2_2 _30306_ (.A(net305),
    .B(\tholin_riscv.regs[18][19] ),
    .Y(_23795_));
 sky130_as_sc_hs__nand3_2 _30307_ (.A(net268),
    .B(_23794_),
    .C(_23795_),
    .Y(_23796_));
 sky130_as_sc_hs__nand3_2 _30308_ (.A(net162),
    .B(_23793_),
    .C(_23796_),
    .Y(_23797_));
 sky130_as_sc_hs__or2_2 _30310_ (.A(net306),
    .B(\tholin_riscv.regs[22][19] ),
    .Y(_23799_));
 sky130_as_sc_hs__nand3_2 _30311_ (.A(net269),
    .B(_23798_),
    .C(_23799_),
    .Y(_23800_));
 sky130_as_sc_hs__or2_2 _30313_ (.A(net306),
    .B(\tholin_riscv.regs[20][19] ),
    .Y(_23802_));
 sky130_as_sc_hs__nand3_2 _30314_ (.A(net172),
    .B(_23801_),
    .C(_23802_),
    .Y(_23803_));
 sky130_as_sc_hs__nand3_2 _30315_ (.A(net254),
    .B(_23800_),
    .C(_23803_),
    .Y(_23804_));
 sky130_as_sc_hs__nand3_2 _30316_ (.A(net154),
    .B(_23797_),
    .C(_23804_),
    .Y(_23805_));
 sky130_as_sc_hs__nand3_2 _30317_ (.A(net251),
    .B(_23783_),
    .C(_23790_),
    .Y(_23806_));
 sky130_as_sc_hs__nand3_2 _30318_ (.A(net247),
    .B(_23805_),
    .C(_23806_),
    .Y(_23807_));
 sky130_as_sc_hs__or2_2 _30320_ (.A(net321),
    .B(\tholin_riscv.regs[8][19] ),
    .Y(_23809_));
 sky130_as_sc_hs__nand3_2 _30321_ (.A(net182),
    .B(_23808_),
    .C(_23809_),
    .Y(_23810_));
 sky130_as_sc_hs__or2_2 _30323_ (.A(net321),
    .B(\tholin_riscv.regs[10][19] ),
    .Y(_23812_));
 sky130_as_sc_hs__nand3_2 _30324_ (.A(net277),
    .B(_23811_),
    .C(_23812_),
    .Y(_23813_));
 sky130_as_sc_hs__nand3_2 _30325_ (.A(net163),
    .B(_23810_),
    .C(_23813_),
    .Y(_23814_));
 sky130_as_sc_hs__or2_2 _30327_ (.A(net321),
    .B(\tholin_riscv.regs[12][19] ),
    .Y(_23816_));
 sky130_as_sc_hs__nand3_2 _30328_ (.A(net182),
    .B(_23815_),
    .C(_23816_),
    .Y(_23817_));
 sky130_as_sc_hs__or2_2 _30330_ (.A(net321),
    .B(\tholin_riscv.regs[14][19] ),
    .Y(_23819_));
 sky130_as_sc_hs__nand3_2 _30331_ (.A(net277),
    .B(_23818_),
    .C(_23819_),
    .Y(_23820_));
 sky130_as_sc_hs__nand3_2 _30332_ (.A(net260),
    .B(_23817_),
    .C(_23820_),
    .Y(_23821_));
 sky130_as_sc_hs__or2_2 _30334_ (.A(net323),
    .B(\tholin_riscv.regs[0][19] ),
    .Y(_23823_));
 sky130_as_sc_hs__nand3_2 _30335_ (.A(net182),
    .B(_23822_),
    .C(_23823_),
    .Y(_23824_));
 sky130_as_sc_hs__or2_2 _30337_ (.A(net321),
    .B(\tholin_riscv.regs[2][19] ),
    .Y(_23826_));
 sky130_as_sc_hs__nand3_2 _30338_ (.A(net277),
    .B(_23825_),
    .C(_23826_),
    .Y(_23827_));
 sky130_as_sc_hs__nand3_2 _30339_ (.A(net163),
    .B(_23824_),
    .C(_23827_),
    .Y(_23828_));
 sky130_as_sc_hs__or2_2 _30341_ (.A(net333),
    .B(\tholin_riscv.regs[6][19] ),
    .Y(_23830_));
 sky130_as_sc_hs__nand3_2 _30342_ (.A(net277),
    .B(_23829_),
    .C(_23830_),
    .Y(_23831_));
 sky130_as_sc_hs__or2_2 _30344_ (.A(net321),
    .B(\tholin_riscv.regs[4][19] ),
    .Y(_23833_));
 sky130_as_sc_hs__nand3_2 _30345_ (.A(net182),
    .B(_23832_),
    .C(_23833_),
    .Y(_23834_));
 sky130_as_sc_hs__nand3_2 _30346_ (.A(net260),
    .B(_23831_),
    .C(_23834_),
    .Y(_23835_));
 sky130_as_sc_hs__nand3_2 _30347_ (.A(net155),
    .B(_23828_),
    .C(_23835_),
    .Y(_23836_));
 sky130_as_sc_hs__nand3_2 _30348_ (.A(net252),
    .B(_23814_),
    .C(_23821_),
    .Y(_23837_));
 sky130_as_sc_hs__nand3_2 _30349_ (.A(net150),
    .B(_23836_),
    .C(_23837_),
    .Y(_23838_));
 sky130_as_sc_hs__or2_2 _30352_ (.A(net303),
    .B(\tholin_riscv.regs[24][18] ),
    .Y(_23841_));
 sky130_as_sc_hs__nand3_2 _30353_ (.A(net171),
    .B(_23840_),
    .C(_23841_),
    .Y(_23842_));
 sky130_as_sc_hs__or2_2 _30355_ (.A(net303),
    .B(\tholin_riscv.regs[26][18] ),
    .Y(_23844_));
 sky130_as_sc_hs__nand3_2 _30356_ (.A(net268),
    .B(_23843_),
    .C(_23844_),
    .Y(_23845_));
 sky130_as_sc_hs__nand3_2 _30357_ (.A(net162),
    .B(_23842_),
    .C(_23845_),
    .Y(_23846_));
 sky130_as_sc_hs__or2_2 _30359_ (.A(net305),
    .B(\tholin_riscv.regs[28][18] ),
    .Y(_23848_));
 sky130_as_sc_hs__nand3_2 _30360_ (.A(net171),
    .B(_23847_),
    .C(_23848_),
    .Y(_23849_));
 sky130_as_sc_hs__or2_2 _30362_ (.A(net303),
    .B(\tholin_riscv.regs[30][18] ),
    .Y(_23851_));
 sky130_as_sc_hs__nand3_2 _30363_ (.A(net268),
    .B(_23850_),
    .C(_23851_),
    .Y(_23852_));
 sky130_as_sc_hs__nand3_2 _30364_ (.A(net254),
    .B(_23849_),
    .C(_23852_),
    .Y(_23853_));
 sky130_as_sc_hs__or2_2 _30366_ (.A(net303),
    .B(\tholin_riscv.regs[16][18] ),
    .Y(_23855_));
 sky130_as_sc_hs__nand3_2 _30367_ (.A(net171),
    .B(_23854_),
    .C(_23855_),
    .Y(_23856_));
 sky130_as_sc_hs__or2_2 _30369_ (.A(net305),
    .B(\tholin_riscv.regs[18][18] ),
    .Y(_23858_));
 sky130_as_sc_hs__nand3_2 _30370_ (.A(net269),
    .B(_23857_),
    .C(_23858_),
    .Y(_23859_));
 sky130_as_sc_hs__nand3_2 _30371_ (.A(net165),
    .B(_23856_),
    .C(_23859_),
    .Y(_23860_));
 sky130_as_sc_hs__or2_2 _30373_ (.A(net303),
    .B(\tholin_riscv.regs[22][18] ),
    .Y(_23862_));
 sky130_as_sc_hs__nand3_2 _30374_ (.A(net268),
    .B(_23861_),
    .C(_23862_),
    .Y(_23863_));
 sky130_as_sc_hs__or2_2 _30376_ (.A(net304),
    .B(\tholin_riscv.regs[20][18] ),
    .Y(_23865_));
 sky130_as_sc_hs__nand3_2 _30377_ (.A(net171),
    .B(_23864_),
    .C(_23865_),
    .Y(_23866_));
 sky130_as_sc_hs__nand3_2 _30378_ (.A(net254),
    .B(_23863_),
    .C(_23866_),
    .Y(_23867_));
 sky130_as_sc_hs__nand3_2 _30379_ (.A(net154),
    .B(_23860_),
    .C(_23867_),
    .Y(_23868_));
 sky130_as_sc_hs__nand3_2 _30380_ (.A(net251),
    .B(_23846_),
    .C(_23853_),
    .Y(_23869_));
 sky130_as_sc_hs__nand3_2 _30381_ (.A(net247),
    .B(_23868_),
    .C(_23869_),
    .Y(_23870_));
 sky130_as_sc_hs__or2_2 _30383_ (.A(net322),
    .B(\tholin_riscv.regs[8][18] ),
    .Y(_23872_));
 sky130_as_sc_hs__nand3_2 _30384_ (.A(net182),
    .B(_23871_),
    .C(_23872_),
    .Y(_23873_));
 sky130_as_sc_hs__or2_2 _30386_ (.A(net322),
    .B(\tholin_riscv.regs[10][18] ),
    .Y(_23875_));
 sky130_as_sc_hs__nand3_2 _30387_ (.A(net277),
    .B(_23874_),
    .C(_23875_),
    .Y(_23876_));
 sky130_as_sc_hs__nand3_2 _30388_ (.A(net163),
    .B(_23873_),
    .C(_23876_),
    .Y(_23877_));
 sky130_as_sc_hs__or2_2 _30390_ (.A(net322),
    .B(\tholin_riscv.regs[12][18] ),
    .Y(_23879_));
 sky130_as_sc_hs__nand3_2 _30391_ (.A(net182),
    .B(_23878_),
    .C(_23879_),
    .Y(_23880_));
 sky130_as_sc_hs__or2_2 _30393_ (.A(net323),
    .B(\tholin_riscv.regs[14][18] ),
    .Y(_23882_));
 sky130_as_sc_hs__nand3_2 _30394_ (.A(net277),
    .B(_23881_),
    .C(_23882_),
    .Y(_23883_));
 sky130_as_sc_hs__nand3_2 _30395_ (.A(net260),
    .B(_23880_),
    .C(_23883_),
    .Y(_23884_));
 sky130_as_sc_hs__or2_2 _30397_ (.A(net323),
    .B(\tholin_riscv.regs[0][18] ),
    .Y(_23886_));
 sky130_as_sc_hs__nand3_2 _30398_ (.A(net182),
    .B(_23885_),
    .C(_23886_),
    .Y(_23887_));
 sky130_as_sc_hs__or2_2 _30400_ (.A(net323),
    .B(\tholin_riscv.regs[2][18] ),
    .Y(_23889_));
 sky130_as_sc_hs__nand3_2 _30401_ (.A(net277),
    .B(_23888_),
    .C(_23889_),
    .Y(_23890_));
 sky130_as_sc_hs__nand3_2 _30402_ (.A(net163),
    .B(_23887_),
    .C(_23890_),
    .Y(_23891_));
 sky130_as_sc_hs__or2_2 _30404_ (.A(net321),
    .B(\tholin_riscv.regs[6][18] ),
    .Y(_23893_));
 sky130_as_sc_hs__nand3_2 _30405_ (.A(net277),
    .B(_23892_),
    .C(_23893_),
    .Y(_23894_));
 sky130_as_sc_hs__or2_2 _30407_ (.A(net322),
    .B(\tholin_riscv.regs[4][18] ),
    .Y(_23896_));
 sky130_as_sc_hs__nand3_2 _30408_ (.A(net182),
    .B(_23895_),
    .C(_23896_),
    .Y(_23897_));
 sky130_as_sc_hs__nand3_2 _30409_ (.A(net260),
    .B(_23894_),
    .C(_23897_),
    .Y(_23898_));
 sky130_as_sc_hs__nand3_2 _30410_ (.A(net155),
    .B(_23891_),
    .C(_23898_),
    .Y(_23899_));
 sky130_as_sc_hs__nand3_2 _30411_ (.A(net252),
    .B(_23877_),
    .C(_23884_),
    .Y(_23900_));
 sky130_as_sc_hs__nand3_2 _30412_ (.A(net150),
    .B(_23899_),
    .C(_23900_),
    .Y(_23901_));
 sky130_as_sc_hs__inv_2 _30414_ (.Y(_23903_),
    .A(_23902_));
 sky130_as_sc_hs__or2_2 _30416_ (.A(net325),
    .B(\tholin_riscv.regs[24][17] ),
    .Y(_23905_));
 sky130_as_sc_hs__nand3_2 _30417_ (.A(net181),
    .B(_23904_),
    .C(_23905_),
    .Y(_23906_));
 sky130_as_sc_hs__or2_2 _30419_ (.A(net325),
    .B(\tholin_riscv.regs[26][17] ),
    .Y(_23908_));
 sky130_as_sc_hs__nand3_2 _30420_ (.A(net276),
    .B(_23907_),
    .C(_23908_),
    .Y(_23909_));
 sky130_as_sc_hs__nand3_2 _30421_ (.A(net164),
    .B(_23906_),
    .C(_23909_),
    .Y(_23910_));
 sky130_as_sc_hs__or2_2 _30423_ (.A(net325),
    .B(\tholin_riscv.regs[28][17] ),
    .Y(_23912_));
 sky130_as_sc_hs__nand3_2 _30424_ (.A(net181),
    .B(_23911_),
    .C(_23912_),
    .Y(_23913_));
 sky130_as_sc_hs__or2_2 _30426_ (.A(net325),
    .B(\tholin_riscv.regs[30][17] ),
    .Y(_23915_));
 sky130_as_sc_hs__nand3_2 _30427_ (.A(net281),
    .B(_23914_),
    .C(_23915_),
    .Y(_23916_));
 sky130_as_sc_hs__nand3_2 _30428_ (.A(net262),
    .B(_23913_),
    .C(_23916_),
    .Y(_23917_));
 sky130_as_sc_hs__or2_2 _30430_ (.A(net326),
    .B(\tholin_riscv.regs[16][17] ),
    .Y(_23919_));
 sky130_as_sc_hs__nand3_2 _30431_ (.A(net181),
    .B(_23918_),
    .C(_23919_),
    .Y(_23920_));
 sky130_as_sc_hs__or2_2 _30433_ (.A(net326),
    .B(\tholin_riscv.regs[18][17] ),
    .Y(_23922_));
 sky130_as_sc_hs__nand3_2 _30434_ (.A(net276),
    .B(_23921_),
    .C(_23922_),
    .Y(_23923_));
 sky130_as_sc_hs__nand3_2 _30435_ (.A(net164),
    .B(_23920_),
    .C(_23923_),
    .Y(_23924_));
 sky130_as_sc_hs__or2_2 _30437_ (.A(net326),
    .B(\tholin_riscv.regs[22][17] ),
    .Y(_23926_));
 sky130_as_sc_hs__nand3_2 _30438_ (.A(net281),
    .B(_23925_),
    .C(_23926_),
    .Y(_23927_));
 sky130_as_sc_hs__or2_2 _30440_ (.A(net326),
    .B(\tholin_riscv.regs[20][17] ),
    .Y(_23929_));
 sky130_as_sc_hs__nand3_2 _30441_ (.A(net180),
    .B(_23928_),
    .C(_23929_),
    .Y(_23930_));
 sky130_as_sc_hs__nand3_2 _30442_ (.A(net262),
    .B(_23927_),
    .C(_23930_),
    .Y(_23931_));
 sky130_as_sc_hs__nand3_2 _30443_ (.A(net156),
    .B(_23924_),
    .C(_23931_),
    .Y(_23932_));
 sky130_as_sc_hs__nand3_2 _30444_ (.A(net252),
    .B(_23910_),
    .C(_23917_),
    .Y(_23933_));
 sky130_as_sc_hs__nand3_2 _30445_ (.A(net247),
    .B(_23932_),
    .C(_23933_),
    .Y(_23934_));
 sky130_as_sc_hs__or2_2 _30447_ (.A(net327),
    .B(\tholin_riscv.regs[8][17] ),
    .Y(_23936_));
 sky130_as_sc_hs__nand3_2 _30448_ (.A(net183),
    .B(_23935_),
    .C(_23936_),
    .Y(_23937_));
 sky130_as_sc_hs__or2_2 _30450_ (.A(net327),
    .B(\tholin_riscv.regs[10][17] ),
    .Y(_23939_));
 sky130_as_sc_hs__nand3_2 _30451_ (.A(net278),
    .B(_23938_),
    .C(_23939_),
    .Y(_23940_));
 sky130_as_sc_hs__nand3_2 _30452_ (.A(net163),
    .B(_23937_),
    .C(_23940_),
    .Y(_23941_));
 sky130_as_sc_hs__or2_2 _30454_ (.A(net327),
    .B(\tholin_riscv.regs[12][17] ),
    .Y(_23943_));
 sky130_as_sc_hs__nand3_2 _30455_ (.A(net183),
    .B(_23942_),
    .C(_23943_),
    .Y(_23944_));
 sky130_as_sc_hs__or2_2 _30457_ (.A(net327),
    .B(\tholin_riscv.regs[14][17] ),
    .Y(_23946_));
 sky130_as_sc_hs__nand3_2 _30458_ (.A(net278),
    .B(_23945_),
    .C(_23946_),
    .Y(_23947_));
 sky130_as_sc_hs__nand3_2 _30459_ (.A(net261),
    .B(_23944_),
    .C(_23947_),
    .Y(_23948_));
 sky130_as_sc_hs__or2_2 _30461_ (.A(net327),
    .B(\tholin_riscv.regs[0][17] ),
    .Y(_23950_));
 sky130_as_sc_hs__nand3_2 _30462_ (.A(net183),
    .B(_23949_),
    .C(_23950_),
    .Y(_23951_));
 sky130_as_sc_hs__or2_2 _30464_ (.A(net328),
    .B(\tholin_riscv.regs[2][17] ),
    .Y(_23953_));
 sky130_as_sc_hs__nand3_2 _30465_ (.A(net279),
    .B(_23952_),
    .C(_23953_),
    .Y(_23954_));
 sky130_as_sc_hs__nand3_2 _30466_ (.A(net163),
    .B(_23951_),
    .C(_23954_),
    .Y(_23955_));
 sky130_as_sc_hs__or2_2 _30468_ (.A(net327),
    .B(\tholin_riscv.regs[6][17] ),
    .Y(_23957_));
 sky130_as_sc_hs__nand3_2 _30469_ (.A(net278),
    .B(_23956_),
    .C(_23957_),
    .Y(_23958_));
 sky130_as_sc_hs__or2_2 _30471_ (.A(net327),
    .B(\tholin_riscv.regs[4][17] ),
    .Y(_23960_));
 sky130_as_sc_hs__nand3_2 _30472_ (.A(net183),
    .B(_23959_),
    .C(_23960_),
    .Y(_23961_));
 sky130_as_sc_hs__nand3_2 _30473_ (.A(net261),
    .B(_23958_),
    .C(_23961_),
    .Y(_23962_));
 sky130_as_sc_hs__nand3_2 _30474_ (.A(net155),
    .B(_23955_),
    .C(_23962_),
    .Y(_23963_));
 sky130_as_sc_hs__nand3_2 _30475_ (.A(net252),
    .B(_23941_),
    .C(_23948_),
    .Y(_23964_));
 sky130_as_sc_hs__nand3_2 _30476_ (.A(net150),
    .B(_23963_),
    .C(_23964_),
    .Y(_23965_));
 sky130_as_sc_hs__inv_2 _30478_ (.Y(_23967_),
    .A(_23966_));
 sky130_as_sc_hs__and2_2 _30479_ (.A(_20449_),
    .B(_20535_),
    .Y(_23968_));
 sky130_as_sc_hs__nor2_2 _30480_ (.A(_20622_),
    .B(_20707_),
    .Y(_23969_));
 sky130_as_sc_hs__and2_2 _30481_ (.A(_23968_),
    .B(_23969_),
    .Y(_23970_));
 sky130_as_sc_hs__and2_2 _30482_ (.A(_20105_),
    .B(_20191_),
    .Y(_23971_));
 sky130_as_sc_hs__and2_2 _30483_ (.A(_20277_),
    .B(_20363_),
    .Y(_23972_));
 sky130_as_sc_hs__nand3_2 _30484_ (.A(_23970_),
    .B(_23971_),
    .C(_23972_),
    .Y(_23973_));
 sky130_as_sc_hs__nor2_2 _30485_ (.A(_23616_),
    .B(_23973_),
    .Y(_23974_));
 sky130_as_sc_hs__or2_2 _30487_ (.A(net324),
    .B(\tholin_riscv.regs[24][16] ),
    .Y(_23976_));
 sky130_as_sc_hs__nand3_2 _30488_ (.A(net180),
    .B(_23975_),
    .C(_23976_),
    .Y(_23977_));
 sky130_as_sc_hs__or2_2 _30490_ (.A(net326),
    .B(\tholin_riscv.regs[26][16] ),
    .Y(_23979_));
 sky130_as_sc_hs__nand3_2 _30491_ (.A(net276),
    .B(_23978_),
    .C(_23979_),
    .Y(_23980_));
 sky130_as_sc_hs__nand3_2 _30492_ (.A(net164),
    .B(_23977_),
    .C(_23980_),
    .Y(_23981_));
 sky130_as_sc_hs__or2_2 _30494_ (.A(net324),
    .B(\tholin_riscv.regs[28][16] ),
    .Y(_23983_));
 sky130_as_sc_hs__nand3_2 _30495_ (.A(net180),
    .B(_23982_),
    .C(_23983_),
    .Y(_23984_));
 sky130_as_sc_hs__or2_2 _30497_ (.A(net326),
    .B(\tholin_riscv.regs[30][16] ),
    .Y(_23986_));
 sky130_as_sc_hs__nand3_2 _30498_ (.A(net276),
    .B(_23985_),
    .C(_23986_),
    .Y(_23987_));
 sky130_as_sc_hs__nand3_2 _30499_ (.A(net260),
    .B(_23984_),
    .C(_23987_),
    .Y(_23988_));
 sky130_as_sc_hs__or2_2 _30501_ (.A(net326),
    .B(\tholin_riscv.regs[16][16] ),
    .Y(_23990_));
 sky130_as_sc_hs__nand3_2 _30502_ (.A(net180),
    .B(_23989_),
    .C(_23990_),
    .Y(_23991_));
 sky130_as_sc_hs__or2_2 _30504_ (.A(net326),
    .B(\tholin_riscv.regs[18][16] ),
    .Y(_23993_));
 sky130_as_sc_hs__nand3_2 _30505_ (.A(net276),
    .B(_23992_),
    .C(_23993_),
    .Y(_23994_));
 sky130_as_sc_hs__nand3_2 _30506_ (.A(net164),
    .B(_23991_),
    .C(_23994_),
    .Y(_23995_));
 sky130_as_sc_hs__or2_2 _30508_ (.A(net324),
    .B(\tholin_riscv.regs[22][16] ),
    .Y(_23997_));
 sky130_as_sc_hs__nand3_2 _30509_ (.A(net276),
    .B(_23996_),
    .C(_23997_),
    .Y(_23998_));
 sky130_as_sc_hs__or2_2 _30511_ (.A(net324),
    .B(\tholin_riscv.regs[20][16] ),
    .Y(_24000_));
 sky130_as_sc_hs__nand3_2 _30512_ (.A(net180),
    .B(_23999_),
    .C(_24000_),
    .Y(_24001_));
 sky130_as_sc_hs__nand3_2 _30513_ (.A(net260),
    .B(_23998_),
    .C(_24001_),
    .Y(_24002_));
 sky130_as_sc_hs__nand3_2 _30514_ (.A(net154),
    .B(_23995_),
    .C(_24002_),
    .Y(_24003_));
 sky130_as_sc_hs__nand3_2 _30515_ (.A(net253),
    .B(_23981_),
    .C(_23988_),
    .Y(_24004_));
 sky130_as_sc_hs__nand3_2 _30516_ (.A(net247),
    .B(_24003_),
    .C(_24004_),
    .Y(_24005_));
 sky130_as_sc_hs__or2_2 _30518_ (.A(net330),
    .B(\tholin_riscv.regs[8][16] ),
    .Y(_24007_));
 sky130_as_sc_hs__nand3_2 _30519_ (.A(net185),
    .B(_24006_),
    .C(_24007_),
    .Y(_24008_));
 sky130_as_sc_hs__or2_2 _30521_ (.A(net331),
    .B(\tholin_riscv.regs[10][16] ),
    .Y(_24010_));
 sky130_as_sc_hs__nand3_2 _30522_ (.A(net281),
    .B(_24009_),
    .C(_24010_),
    .Y(_24011_));
 sky130_as_sc_hs__nand3_2 _30523_ (.A(net164),
    .B(_24008_),
    .C(_24011_),
    .Y(_24012_));
 sky130_as_sc_hs__or2_2 _30525_ (.A(net330),
    .B(\tholin_riscv.regs[12][16] ),
    .Y(_24014_));
 sky130_as_sc_hs__nand3_2 _30526_ (.A(net185),
    .B(_24013_),
    .C(_24014_),
    .Y(_24015_));
 sky130_as_sc_hs__or2_2 _30528_ (.A(net330),
    .B(\tholin_riscv.regs[14][16] ),
    .Y(_24017_));
 sky130_as_sc_hs__nand3_2 _30529_ (.A(net280),
    .B(_24016_),
    .C(_24017_),
    .Y(_24018_));
 sky130_as_sc_hs__nand3_2 _30530_ (.A(net261),
    .B(_24015_),
    .C(_24018_),
    .Y(_24019_));
 sky130_as_sc_hs__or2_2 _30532_ (.A(net330),
    .B(\tholin_riscv.regs[0][16] ),
    .Y(_24021_));
 sky130_as_sc_hs__nand3_2 _30533_ (.A(net185),
    .B(_24020_),
    .C(_24021_),
    .Y(_24022_));
 sky130_as_sc_hs__or2_2 _30535_ (.A(net330),
    .B(\tholin_riscv.regs[2][16] ),
    .Y(_24024_));
 sky130_as_sc_hs__nand3_2 _30536_ (.A(net280),
    .B(_24023_),
    .C(_24024_),
    .Y(_24025_));
 sky130_as_sc_hs__nand3_2 _30537_ (.A(net165),
    .B(_24022_),
    .C(_24025_),
    .Y(_24026_));
 sky130_as_sc_hs__or2_2 _30539_ (.A(net330),
    .B(\tholin_riscv.regs[6][16] ),
    .Y(_24028_));
 sky130_as_sc_hs__nand3_2 _30540_ (.A(net280),
    .B(_24027_),
    .C(_24028_),
    .Y(_24029_));
 sky130_as_sc_hs__or2_2 _30542_ (.A(net330),
    .B(\tholin_riscv.regs[4][16] ),
    .Y(_24031_));
 sky130_as_sc_hs__nand3_2 _30543_ (.A(net185),
    .B(_24030_),
    .C(_24031_),
    .Y(_24032_));
 sky130_as_sc_hs__nand3_2 _30544_ (.A(net261),
    .B(_24029_),
    .C(_24032_),
    .Y(_24033_));
 sky130_as_sc_hs__nand3_2 _30545_ (.A(net155),
    .B(_24026_),
    .C(_24033_),
    .Y(_24034_));
 sky130_as_sc_hs__nand3_2 _30546_ (.A(net253),
    .B(_24012_),
    .C(_24019_),
    .Y(_24035_));
 sky130_as_sc_hs__nand3_2 _30547_ (.A(net150),
    .B(_24034_),
    .C(_24035_),
    .Y(_24036_));
 sky130_as_sc_hs__nand3_2 _30550_ (.A(_23966_),
    .B(_23974_),
    .C(_24037_),
    .Y(_24039_));
 sky130_as_sc_hs__nor2_2 _30551_ (.A(_23903_),
    .B(_24039_),
    .Y(_24040_));
 sky130_as_sc_hs__nand3_2 _30553_ (.A(_23775_),
    .B(_23839_),
    .C(_24040_),
    .Y(_24042_));
 sky130_as_sc_hs__and2_2 _30558_ (.A(_24045_),
    .B(_24046_),
    .Y(_24047_));
 sky130_as_sc_hs__and2_2 _30559_ (.A(_23712_),
    .B(net470),
    .Y(_24048_));
 sky130_as_sc_hs__and2_2 _30561_ (.A(_21977_),
    .B(_22170_),
    .Y(_24050_));
 sky130_as_sc_hs__nor2_2 _30562_ (.A(_22171_),
    .B(_24050_),
    .Y(_24051_));
 sky130_as_sc_hs__or2_2 _30566_ (.A(net324),
    .B(\tholin_riscv.regs[24][21] ),
    .Y(_24055_));
 sky130_as_sc_hs__nand3_2 _30567_ (.A(net180),
    .B(_24054_),
    .C(_24055_),
    .Y(_24056_));
 sky130_as_sc_hs__or2_2 _30569_ (.A(net324),
    .B(\tholin_riscv.regs[26][21] ),
    .Y(_24058_));
 sky130_as_sc_hs__nand3_2 _30570_ (.A(net276),
    .B(_24057_),
    .C(_24058_),
    .Y(_24059_));
 sky130_as_sc_hs__nand3_2 _30571_ (.A(net164),
    .B(_24056_),
    .C(_24059_),
    .Y(_24060_));
 sky130_as_sc_hs__or2_2 _30573_ (.A(net324),
    .B(\tholin_riscv.regs[28][21] ),
    .Y(_24062_));
 sky130_as_sc_hs__nand3_2 _30574_ (.A(net180),
    .B(_24061_),
    .C(_24062_),
    .Y(_24063_));
 sky130_as_sc_hs__or2_2 _30576_ (.A(net324),
    .B(\tholin_riscv.regs[30][21] ),
    .Y(_24065_));
 sky130_as_sc_hs__nand3_2 _30577_ (.A(net276),
    .B(_24064_),
    .C(_24065_),
    .Y(_24066_));
 sky130_as_sc_hs__nand3_2 _30578_ (.A(net260),
    .B(_24063_),
    .C(_24066_),
    .Y(_24067_));
 sky130_as_sc_hs__or2_2 _30580_ (.A(net324),
    .B(\tholin_riscv.regs[16][21] ),
    .Y(_24069_));
 sky130_as_sc_hs__nand3_2 _30581_ (.A(net180),
    .B(_24068_),
    .C(_24069_),
    .Y(_24070_));
 sky130_as_sc_hs__or2_2 _30583_ (.A(net324),
    .B(\tholin_riscv.regs[18][21] ),
    .Y(_24072_));
 sky130_as_sc_hs__nand3_2 _30584_ (.A(net276),
    .B(_24071_),
    .C(_24072_),
    .Y(_24073_));
 sky130_as_sc_hs__nand3_2 _30585_ (.A(net164),
    .B(_24070_),
    .C(_24073_),
    .Y(_24074_));
 sky130_as_sc_hs__or2_2 _30587_ (.A(net325),
    .B(\tholin_riscv.regs[22][21] ),
    .Y(_24076_));
 sky130_as_sc_hs__nand3_2 _30588_ (.A(net276),
    .B(_24075_),
    .C(_24076_),
    .Y(_24077_));
 sky130_as_sc_hs__or2_2 _30590_ (.A(net325),
    .B(\tholin_riscv.regs[20][21] ),
    .Y(_24079_));
 sky130_as_sc_hs__nand3_2 _30591_ (.A(net181),
    .B(_24078_),
    .C(_24079_),
    .Y(_24080_));
 sky130_as_sc_hs__nand3_2 _30592_ (.A(net260),
    .B(_24077_),
    .C(_24080_),
    .Y(_24081_));
 sky130_as_sc_hs__nand3_2 _30593_ (.A(net155),
    .B(_24074_),
    .C(_24081_),
    .Y(_24082_));
 sky130_as_sc_hs__nand3_2 _30594_ (.A(net252),
    .B(_24060_),
    .C(_24067_),
    .Y(_24083_));
 sky130_as_sc_hs__nand3_2 _30595_ (.A(net247),
    .B(_24082_),
    .C(_24083_),
    .Y(_24084_));
 sky130_as_sc_hs__or2_2 _30597_ (.A(net327),
    .B(\tholin_riscv.regs[8][21] ),
    .Y(_24086_));
 sky130_as_sc_hs__nand3_2 _30598_ (.A(net183),
    .B(_24085_),
    .C(_24086_),
    .Y(_24087_));
 sky130_as_sc_hs__or2_2 _30600_ (.A(net327),
    .B(\tholin_riscv.regs[10][21] ),
    .Y(_24089_));
 sky130_as_sc_hs__nand3_2 _30601_ (.A(net278),
    .B(_24088_),
    .C(_24089_),
    .Y(_24090_));
 sky130_as_sc_hs__nand3_2 _30602_ (.A(net165),
    .B(_24087_),
    .C(_24090_),
    .Y(_24091_));
 sky130_as_sc_hs__or2_2 _30604_ (.A(net329),
    .B(\tholin_riscv.regs[12][21] ),
    .Y(_24093_));
 sky130_as_sc_hs__nand3_2 _30605_ (.A(net183),
    .B(_24092_),
    .C(_24093_),
    .Y(_24094_));
 sky130_as_sc_hs__or2_2 _30607_ (.A(net329),
    .B(\tholin_riscv.regs[14][21] ),
    .Y(_24096_));
 sky130_as_sc_hs__nand3_2 _30608_ (.A(net278),
    .B(_24095_),
    .C(_24096_),
    .Y(_24097_));
 sky130_as_sc_hs__nand3_2 _30609_ (.A(net261),
    .B(_24094_),
    .C(_24097_),
    .Y(_24098_));
 sky130_as_sc_hs__or2_2 _30611_ (.A(net329),
    .B(\tholin_riscv.regs[0][21] ),
    .Y(_24100_));
 sky130_as_sc_hs__nand3_2 _30612_ (.A(net184),
    .B(_24099_),
    .C(_24100_),
    .Y(_24101_));
 sky130_as_sc_hs__or2_2 _30614_ (.A(net327),
    .B(\tholin_riscv.regs[2][21] ),
    .Y(_24103_));
 sky130_as_sc_hs__nand3_2 _30615_ (.A(net279),
    .B(_24102_),
    .C(_24103_),
    .Y(_24104_));
 sky130_as_sc_hs__nand3_2 _30616_ (.A(net163),
    .B(_24101_),
    .C(_24104_),
    .Y(_24105_));
 sky130_as_sc_hs__or2_2 _30618_ (.A(net327),
    .B(\tholin_riscv.regs[6][21] ),
    .Y(_24107_));
 sky130_as_sc_hs__nand3_2 _30619_ (.A(net278),
    .B(_24106_),
    .C(_24107_),
    .Y(_24108_));
 sky130_as_sc_hs__or2_2 _30621_ (.A(net329),
    .B(\tholin_riscv.regs[4][21] ),
    .Y(_24110_));
 sky130_as_sc_hs__nand3_2 _30622_ (.A(net183),
    .B(_24109_),
    .C(_24110_),
    .Y(_24111_));
 sky130_as_sc_hs__nand3_2 _30623_ (.A(net261),
    .B(_24108_),
    .C(_24111_),
    .Y(_24112_));
 sky130_as_sc_hs__nand3_2 _30624_ (.A(net155),
    .B(_24105_),
    .C(_24112_),
    .Y(_24113_));
 sky130_as_sc_hs__nand3_2 _30625_ (.A(net252),
    .B(_24091_),
    .C(_24098_),
    .Y(_24114_));
 sky130_as_sc_hs__nand3_2 _30626_ (.A(net151),
    .B(_24113_),
    .C(_24114_),
    .Y(_24115_));
 sky130_as_sc_hs__inv_2 _30628_ (.Y(_24117_),
    .A(_24116_));
 sky130_as_sc_hs__or2_2 _30629_ (.A(_24042_),
    .B(_24117_),
    .Y(_24118_));
 sky130_as_sc_hs__and2_2 _30634_ (.A(_24121_),
    .B(_24122_),
    .Y(_24123_));
 sky130_as_sc_hs__and2_2 _30635_ (.A(_24053_),
    .B(net468),
    .Y(_24124_));
 sky130_as_sc_hs__and2_2 _30636_ (.A(_21659_),
    .B(_22169_),
    .Y(_24125_));
 sky130_as_sc_hs__or2_2 _30637_ (.A(_22040_),
    .B(_24125_),
    .Y(_24126_));
 sky130_as_sc_hs__and2_2 _30639_ (.A(_24126_),
    .B(_24127_),
    .Y(_24128_));
 sky130_as_sc_hs__or2_2 _30641_ (.A(net297),
    .B(\tholin_riscv.regs[24][22] ),
    .Y(_24130_));
 sky130_as_sc_hs__nand3_2 _30642_ (.A(net169),
    .B(_24129_),
    .C(_24130_),
    .Y(_24131_));
 sky130_as_sc_hs__or2_2 _30644_ (.A(net297),
    .B(\tholin_riscv.regs[26][22] ),
    .Y(_24133_));
 sky130_as_sc_hs__nand3_2 _30645_ (.A(net266),
    .B(_24132_),
    .C(_24133_),
    .Y(_24134_));
 sky130_as_sc_hs__nand3_2 _30646_ (.A(net162),
    .B(_24131_),
    .C(_24134_),
    .Y(_24135_));
 sky130_as_sc_hs__or2_2 _30648_ (.A(net304),
    .B(\tholin_riscv.regs[28][22] ),
    .Y(_24137_));
 sky130_as_sc_hs__nand3_2 _30649_ (.A(net171),
    .B(_24136_),
    .C(_24137_),
    .Y(_24138_));
 sky130_as_sc_hs__or2_2 _30651_ (.A(net304),
    .B(\tholin_riscv.regs[30][22] ),
    .Y(_24140_));
 sky130_as_sc_hs__nand3_2 _30652_ (.A(net268),
    .B(_24139_),
    .C(_24140_),
    .Y(_24141_));
 sky130_as_sc_hs__nand3_2 _30653_ (.A(net254),
    .B(_24138_),
    .C(_24141_),
    .Y(_24142_));
 sky130_as_sc_hs__or2_2 _30655_ (.A(net304),
    .B(\tholin_riscv.regs[16][22] ),
    .Y(_24144_));
 sky130_as_sc_hs__nand3_2 _30656_ (.A(net171),
    .B(_24143_),
    .C(_24144_),
    .Y(_24145_));
 sky130_as_sc_hs__or2_2 _30658_ (.A(net304),
    .B(\tholin_riscv.regs[18][22] ),
    .Y(_24147_));
 sky130_as_sc_hs__nand3_2 _30659_ (.A(net268),
    .B(_24146_),
    .C(_24147_),
    .Y(_24148_));
 sky130_as_sc_hs__nand3_2 _30660_ (.A(net162),
    .B(_24145_),
    .C(_24148_),
    .Y(_24149_));
 sky130_as_sc_hs__or2_2 _30662_ (.A(net298),
    .B(\tholin_riscv.regs[22][22] ),
    .Y(_24151_));
 sky130_as_sc_hs__nand3_2 _30663_ (.A(net266),
    .B(_24150_),
    .C(_24151_),
    .Y(_24152_));
 sky130_as_sc_hs__or2_2 _30665_ (.A(net298),
    .B(\tholin_riscv.regs[20][22] ),
    .Y(_24154_));
 sky130_as_sc_hs__nand3_2 _30666_ (.A(net168),
    .B(_24153_),
    .C(_24154_),
    .Y(_24155_));
 sky130_as_sc_hs__nand3_2 _30667_ (.A(net255),
    .B(_24152_),
    .C(_24155_),
    .Y(_24156_));
 sky130_as_sc_hs__nand3_2 _30668_ (.A(net154),
    .B(_24149_),
    .C(_24156_),
    .Y(_24157_));
 sky130_as_sc_hs__nand3_2 _30669_ (.A(net251),
    .B(_24135_),
    .C(_24142_),
    .Y(_24158_));
 sky130_as_sc_hs__nand3_2 _30670_ (.A(net247),
    .B(_24157_),
    .C(_24158_),
    .Y(_24159_));
 sky130_as_sc_hs__or2_2 _30672_ (.A(net322),
    .B(\tholin_riscv.regs[8][22] ),
    .Y(_24161_));
 sky130_as_sc_hs__nand3_2 _30673_ (.A(net180),
    .B(_24160_),
    .C(_24161_),
    .Y(_24162_));
 sky130_as_sc_hs__or2_2 _30675_ (.A(net322),
    .B(\tholin_riscv.regs[10][22] ),
    .Y(_24164_));
 sky130_as_sc_hs__nand3_2 _30676_ (.A(net276),
    .B(_24163_),
    .C(_24164_),
    .Y(_24165_));
 sky130_as_sc_hs__nand3_2 _30677_ (.A(net162),
    .B(_24162_),
    .C(_24165_),
    .Y(_24166_));
 sky130_as_sc_hs__or2_2 _30679_ (.A(net324),
    .B(\tholin_riscv.regs[12][22] ),
    .Y(_24168_));
 sky130_as_sc_hs__nand3_2 _30680_ (.A(net180),
    .B(_24167_),
    .C(_24168_),
    .Y(_24169_));
 sky130_as_sc_hs__or2_2 _30682_ (.A(net324),
    .B(\tholin_riscv.regs[14][22] ),
    .Y(_24171_));
 sky130_as_sc_hs__nand3_2 _30683_ (.A(net276),
    .B(_24170_),
    .C(_24171_),
    .Y(_24172_));
 sky130_as_sc_hs__nand3_2 _30684_ (.A(net260),
    .B(_24169_),
    .C(_24172_),
    .Y(_24173_));
 sky130_as_sc_hs__or2_2 _30686_ (.A(net322),
    .B(\tholin_riscv.regs[0][22] ),
    .Y(_24175_));
 sky130_as_sc_hs__nand3_2 _30687_ (.A(net180),
    .B(_24174_),
    .C(_24175_),
    .Y(_24176_));
 sky130_as_sc_hs__or2_2 _30689_ (.A(net324),
    .B(\tholin_riscv.regs[2][22] ),
    .Y(_24178_));
 sky130_as_sc_hs__nand3_2 _30690_ (.A(net276),
    .B(_24177_),
    .C(_24178_),
    .Y(_24179_));
 sky130_as_sc_hs__nand3_2 _30691_ (.A(net164),
    .B(_24176_),
    .C(_24179_),
    .Y(_24180_));
 sky130_as_sc_hs__or2_2 _30693_ (.A(net324),
    .B(\tholin_riscv.regs[6][22] ),
    .Y(_24182_));
 sky130_as_sc_hs__nand3_2 _30694_ (.A(net276),
    .B(_24181_),
    .C(_24182_),
    .Y(_24183_));
 sky130_as_sc_hs__or2_2 _30696_ (.A(net324),
    .B(\tholin_riscv.regs[4][22] ),
    .Y(_24185_));
 sky130_as_sc_hs__nand3_2 _30697_ (.A(net180),
    .B(_24184_),
    .C(_24185_),
    .Y(_24186_));
 sky130_as_sc_hs__nand3_2 _30698_ (.A(net262),
    .B(_24183_),
    .C(_24186_),
    .Y(_24187_));
 sky130_as_sc_hs__nand3_2 _30699_ (.A(net156),
    .B(_24180_),
    .C(_24187_),
    .Y(_24188_));
 sky130_as_sc_hs__nand3_2 _30700_ (.A(net253),
    .B(_24166_),
    .C(_24173_),
    .Y(_24189_));
 sky130_as_sc_hs__nand3_2 _30701_ (.A(net151),
    .B(_24188_),
    .C(_24189_),
    .Y(_24190_));
 sky130_as_sc_hs__inv_2 _30703_ (.Y(_24192_),
    .A(_24191_));
 sky130_as_sc_hs__or2_2 _30705_ (.A(_24118_),
    .B(_24192_),
    .Y(_24194_));
 sky130_as_sc_hs__and2_2 _30709_ (.A(_24196_),
    .B(_24197_),
    .Y(_24198_));
 sky130_as_sc_hs__nand3_2 _30710_ (.A(net90),
    .B(_24196_),
    .C(_24197_),
    .Y(_24199_));
 sky130_as_sc_hs__nand3_2 _30711_ (.A(_24124_),
    .B(net90),
    .C(net466),
    .Y(_24200_));
 sky130_as_sc_hs__nand2b_2 _30712_ (.B(_24199_),
    .Y(_24201_),
    .A(_24124_));
 sky130_as_sc_hs__and2_2 _30713_ (.A(_24200_),
    .B(_24201_),
    .Y(_24202_));
 sky130_as_sc_hs__or2_2 _30715_ (.A(_24048_),
    .B(_24202_),
    .Y(_24204_));
 sky130_as_sc_hs__and2_2 _30716_ (.A(_24203_),
    .B(_24204_),
    .Y(_24205_));
 sky130_as_sc_hs__or2_2 _30717_ (.A(_23839_),
    .B(_24040_),
    .Y(_24206_));
 sky130_as_sc_hs__and2_2 _30721_ (.A(_24208_),
    .B(_24209_),
    .Y(_24210_));
 sky130_as_sc_hs__and2_2 _30722_ (.A(_23712_),
    .B(net464),
    .Y(_24211_));
 sky130_as_sc_hs__nand3_2 _30726_ (.A(_21659_),
    .B(_22238_),
    .C(_24213_),
    .Y(_24215_));
 sky130_as_sc_hs__and2_2 _30728_ (.A(_23903_),
    .B(_24039_),
    .Y(_24217_));
 sky130_as_sc_hs__or2_2 _30729_ (.A(_24040_),
    .B(_24217_),
    .Y(_24218_));
 sky130_as_sc_hs__and2_2 _30732_ (.A(_24219_),
    .B(_24220_),
    .Y(_24221_));
 sky130_as_sc_hs__and2_2 _30733_ (.A(_24216_),
    .B(net462),
    .Y(_24222_));
 sky130_as_sc_hs__nand3_2 _30736_ (.A(_22171_),
    .B(_22237_),
    .C(_22365_),
    .Y(_24225_));
 sky130_as_sc_hs__nand3_2 _30739_ (.A(_21659_),
    .B(_24225_),
    .C(_24226_),
    .Y(_24228_));
 sky130_as_sc_hs__and2_2 _30745_ (.A(_24232_),
    .B(_24233_),
    .Y(_24234_));
 sky130_as_sc_hs__and2_2 _30746_ (.A(_24229_),
    .B(net461),
    .Y(_24235_));
 sky130_as_sc_hs__or2_2 _30747_ (.A(_24211_),
    .B(_24222_),
    .Y(_24236_));
 sky130_as_sc_hs__and2_2 _30748_ (.A(_24223_),
    .B(_24236_),
    .Y(_24237_));
 sky130_as_sc_hs__or2_2 _30751_ (.A(_22104_),
    .B(_22168_),
    .Y(_24240_));
 sky130_as_sc_hs__and2_2 _30755_ (.A(_24242_),
    .B(_24243_),
    .Y(_24244_));
 sky130_as_sc_hs__nand3_2 _30756_ (.A(_24196_),
    .B(_24197_),
    .C(net458),
    .Y(_24245_));
 sky130_as_sc_hs__or2_2 _30758_ (.A(_24245_),
    .B(_24246_),
    .Y(_24247_));
 sky130_as_sc_hs__and2_2 _30759_ (.A(net470),
    .B(_24053_),
    .Y(_24248_));
 sky130_as_sc_hs__and2_2 _30761_ (.A(_24247_),
    .B(_24249_),
    .Y(_24250_));
 sky130_as_sc_hs__nand3_2 _30766_ (.A(_21659_),
    .B(_22367_),
    .C(_24254_),
    .Y(_24255_));
 sky130_as_sc_hs__and2_2 _30768_ (.A(net461),
    .B(_24256_),
    .Y(_24257_));
 sky130_as_sc_hs__and2_2 _30769_ (.A(net462),
    .B(_24229_),
    .Y(_24258_));
 sky130_as_sc_hs__and2_2 _30770_ (.A(net464),
    .B(_24216_),
    .Y(_24259_));
 sky130_as_sc_hs__or2_2 _30772_ (.A(_24258_),
    .B(_24259_),
    .Y(_24261_));
 sky130_as_sc_hs__and2_2 _30773_ (.A(_24260_),
    .B(_24261_),
    .Y(_24262_));
 sky130_as_sc_hs__or2_2 _30775_ (.A(_24257_),
    .B(_24262_),
    .Y(_24264_));
 sky130_as_sc_hs__and2_2 _30776_ (.A(_24263_),
    .B(_24264_),
    .Y(_24265_));
 sky130_as_sc_hs__or2_2 _30778_ (.A(_24252_),
    .B(_24265_),
    .Y(_24267_));
 sky130_as_sc_hs__and2_2 _30779_ (.A(_24266_),
    .B(_24267_),
    .Y(_24268_));
 sky130_as_sc_hs__or2_2 _30781_ (.A(_24239_),
    .B(_24268_),
    .Y(_24270_));
 sky130_as_sc_hs__and2_2 _30782_ (.A(_24269_),
    .B(_24270_),
    .Y(_24271_));
 sky130_as_sc_hs__or2_2 _30784_ (.A(net200),
    .B(\tholin_riscv.regs[25][25] ),
    .Y(_24273_));
 sky130_as_sc_hs__or2_2 _30785_ (.A(net325),
    .B(\tholin_riscv.regs[24][25] ),
    .Y(_24274_));
 sky130_as_sc_hs__nand3_2 _30786_ (.A(net181),
    .B(_24273_),
    .C(_24274_),
    .Y(_24275_));
 sky130_as_sc_hs__or2_2 _30787_ (.A(net200),
    .B(\tholin_riscv.regs[27][25] ),
    .Y(_24276_));
 sky130_as_sc_hs__or2_2 _30788_ (.A(net332),
    .B(\tholin_riscv.regs[26][25] ),
    .Y(_24277_));
 sky130_as_sc_hs__nand3_2 _30789_ (.A(net280),
    .B(_24276_),
    .C(_24277_),
    .Y(_24278_));
 sky130_as_sc_hs__nand3_2 _30790_ (.A(net164),
    .B(_24275_),
    .C(_24278_),
    .Y(_24279_));
 sky130_as_sc_hs__or2_2 _30791_ (.A(net196),
    .B(\tholin_riscv.regs[29][25] ),
    .Y(_24280_));
 sky130_as_sc_hs__or2_2 _30792_ (.A(net325),
    .B(\tholin_riscv.regs[28][25] ),
    .Y(_24281_));
 sky130_as_sc_hs__nand3_2 _30793_ (.A(net181),
    .B(_24280_),
    .C(_24281_),
    .Y(_24282_));
 sky130_as_sc_hs__or2_2 _30794_ (.A(net196),
    .B(\tholin_riscv.regs[31][25] ),
    .Y(_24283_));
 sky130_as_sc_hs__or2_2 _30795_ (.A(net325),
    .B(\tholin_riscv.regs[30][25] ),
    .Y(_24284_));
 sky130_as_sc_hs__nand3_2 _30796_ (.A(net281),
    .B(_24283_),
    .C(_24284_),
    .Y(_24285_));
 sky130_as_sc_hs__nand3_2 _30797_ (.A(net260),
    .B(_24282_),
    .C(_24285_),
    .Y(_24286_));
 sky130_as_sc_hs__or2_2 _30798_ (.A(net199),
    .B(\tholin_riscv.regs[17][25] ),
    .Y(_24287_));
 sky130_as_sc_hs__or2_2 _30799_ (.A(net331),
    .B(\tholin_riscv.regs[16][25] ),
    .Y(_24288_));
 sky130_as_sc_hs__nand3_2 _30800_ (.A(net185),
    .B(_24287_),
    .C(_24288_),
    .Y(_24289_));
 sky130_as_sc_hs__or2_2 _30801_ (.A(net199),
    .B(\tholin_riscv.regs[19][25] ),
    .Y(_24290_));
 sky130_as_sc_hs__or2_2 _30802_ (.A(net331),
    .B(\tholin_riscv.regs[18][25] ),
    .Y(_24291_));
 sky130_as_sc_hs__nand3_2 _30803_ (.A(net280),
    .B(_24290_),
    .C(_24291_),
    .Y(_24292_));
 sky130_as_sc_hs__nand3_2 _30804_ (.A(net164),
    .B(_24289_),
    .C(_24292_),
    .Y(_24293_));
 sky130_as_sc_hs__or2_2 _30805_ (.A(net199),
    .B(\tholin_riscv.regs[23][25] ),
    .Y(_24294_));
 sky130_as_sc_hs__or2_2 _30806_ (.A(net332),
    .B(\tholin_riscv.regs[22][25] ),
    .Y(_24295_));
 sky130_as_sc_hs__nand3_2 _30807_ (.A(net280),
    .B(_24294_),
    .C(_24295_),
    .Y(_24296_));
 sky130_as_sc_hs__or2_2 _30808_ (.A(net199),
    .B(\tholin_riscv.regs[21][25] ),
    .Y(_24297_));
 sky130_as_sc_hs__or2_2 _30809_ (.A(net331),
    .B(\tholin_riscv.regs[20][25] ),
    .Y(_24298_));
 sky130_as_sc_hs__nand3_2 _30810_ (.A(net185),
    .B(_24297_),
    .C(_24298_),
    .Y(_24299_));
 sky130_as_sc_hs__nand3_2 _30811_ (.A(net262),
    .B(_24296_),
    .C(_24299_),
    .Y(_24300_));
 sky130_as_sc_hs__nand3_2 _30812_ (.A(net155),
    .B(_24293_),
    .C(_24300_),
    .Y(_24301_));
 sky130_as_sc_hs__nand3_2 _30813_ (.A(net252),
    .B(_24279_),
    .C(_24286_),
    .Y(_24302_));
 sky130_as_sc_hs__nor2_2 _30815_ (.A(net151),
    .B(_24303_),
    .Y(_24304_));
 sky130_as_sc_hs__or2_2 _30816_ (.A(net187),
    .B(\tholin_riscv.regs[9][25] ),
    .Y(_24305_));
 sky130_as_sc_hs__or2_2 _30817_ (.A(net286),
    .B(\tholin_riscv.regs[8][25] ),
    .Y(_24306_));
 sky130_as_sc_hs__nand3_2 _30818_ (.A(net166),
    .B(_24305_),
    .C(_24306_),
    .Y(_24307_));
 sky130_as_sc_hs__or2_2 _30819_ (.A(net187),
    .B(\tholin_riscv.regs[11][25] ),
    .Y(_24308_));
 sky130_as_sc_hs__or2_2 _30820_ (.A(net286),
    .B(\tholin_riscv.regs[10][25] ),
    .Y(_24309_));
 sky130_as_sc_hs__nand3_2 _30821_ (.A(net263),
    .B(_24308_),
    .C(_24309_),
    .Y(_24310_));
 sky130_as_sc_hs__nand3_2 _30822_ (.A(net157),
    .B(_24307_),
    .C(_24310_),
    .Y(_24311_));
 sky130_as_sc_hs__or2_2 _30823_ (.A(net187),
    .B(\tholin_riscv.regs[13][25] ),
    .Y(_24312_));
 sky130_as_sc_hs__or2_2 _30824_ (.A(net308),
    .B(\tholin_riscv.regs[12][25] ),
    .Y(_24313_));
 sky130_as_sc_hs__nand3_2 _30825_ (.A(net166),
    .B(_24312_),
    .C(_24313_),
    .Y(_24314_));
 sky130_as_sc_hs__or2_2 _30826_ (.A(net187),
    .B(\tholin_riscv.regs[15][25] ),
    .Y(_24315_));
 sky130_as_sc_hs__or2_2 _30827_ (.A(net286),
    .B(\tholin_riscv.regs[14][25] ),
    .Y(_24316_));
 sky130_as_sc_hs__nand3_2 _30828_ (.A(net263),
    .B(_24315_),
    .C(_24316_),
    .Y(_24317_));
 sky130_as_sc_hs__nand3_2 _30829_ (.A(net256),
    .B(_24314_),
    .C(_24317_),
    .Y(_24318_));
 sky130_as_sc_hs__or2_2 _30830_ (.A(net187),
    .B(\tholin_riscv.regs[1][25] ),
    .Y(_24319_));
 sky130_as_sc_hs__or2_2 _30831_ (.A(net308),
    .B(\tholin_riscv.regs[0][25] ),
    .Y(_24320_));
 sky130_as_sc_hs__nand3_2 _30832_ (.A(net174),
    .B(_24319_),
    .C(_24320_),
    .Y(_24321_));
 sky130_as_sc_hs__or2_2 _30833_ (.A(net187),
    .B(\tholin_riscv.regs[3][25] ),
    .Y(_24322_));
 sky130_as_sc_hs__or2_2 _30834_ (.A(net308),
    .B(\tholin_riscv.regs[2][25] ),
    .Y(_24323_));
 sky130_as_sc_hs__nand3_2 _30835_ (.A(net270),
    .B(_24322_),
    .C(_24323_),
    .Y(_24324_));
 sky130_as_sc_hs__nand3_2 _30836_ (.A(net157),
    .B(_24321_),
    .C(_24324_),
    .Y(_24325_));
 sky130_as_sc_hs__or2_2 _30837_ (.A(net187),
    .B(\tholin_riscv.regs[7][25] ),
    .Y(_24326_));
 sky130_as_sc_hs__or2_2 _30838_ (.A(net308),
    .B(\tholin_riscv.regs[6][25] ),
    .Y(_24327_));
 sky130_as_sc_hs__nand3_2 _30839_ (.A(net270),
    .B(_24326_),
    .C(_24327_),
    .Y(_24328_));
 sky130_as_sc_hs__or2_2 _30840_ (.A(net187),
    .B(\tholin_riscv.regs[5][25] ),
    .Y(_24329_));
 sky130_as_sc_hs__or2_2 _30841_ (.A(net308),
    .B(\tholin_riscv.regs[4][25] ),
    .Y(_24330_));
 sky130_as_sc_hs__nand3_2 _30842_ (.A(net174),
    .B(_24329_),
    .C(_24330_),
    .Y(_24331_));
 sky130_as_sc_hs__nand3_2 _30843_ (.A(net257),
    .B(_24328_),
    .C(_24331_),
    .Y(_24332_));
 sky130_as_sc_hs__nand3_2 _30844_ (.A(net153),
    .B(_24325_),
    .C(_24332_),
    .Y(_24333_));
 sky130_as_sc_hs__nand3_2 _30845_ (.A(net250),
    .B(_24311_),
    .C(_24318_),
    .Y(_24334_));
 sky130_as_sc_hs__and2_2 _30846_ (.A(_24333_),
    .B(_24334_),
    .Y(_24335_));
 sky130_as_sc_hs__and2_2 _30847_ (.A(net151),
    .B(_24335_),
    .Y(_24336_));
 sky130_as_sc_hs__nor2_2 _30848_ (.A(_24304_),
    .B(_24336_),
    .Y(_24337_));
 sky130_as_sc_hs__or2_2 _30849_ (.A(_24304_),
    .B(_24336_),
    .Y(_24338_));
 sky130_as_sc_hs__and2_2 _30850_ (.A(_23839_),
    .B(_23902_),
    .Y(_24339_));
 sky130_as_sc_hs__nand3_2 _30851_ (.A(_23966_),
    .B(_24037_),
    .C(_24339_),
    .Y(_24340_));
 sky130_as_sc_hs__or2_2 _30853_ (.A(net298),
    .B(\tholin_riscv.regs[24][23] ),
    .Y(_24342_));
 sky130_as_sc_hs__nand3_2 _30854_ (.A(net169),
    .B(_24341_),
    .C(_24342_),
    .Y(_24343_));
 sky130_as_sc_hs__or2_2 _30856_ (.A(net298),
    .B(\tholin_riscv.regs[26][23] ),
    .Y(_24345_));
 sky130_as_sc_hs__nand3_2 _30857_ (.A(net266),
    .B(_24344_),
    .C(_24345_),
    .Y(_24346_));
 sky130_as_sc_hs__nand3_2 _30858_ (.A(net162),
    .B(_24343_),
    .C(_24346_),
    .Y(_24347_));
 sky130_as_sc_hs__or2_2 _30860_ (.A(net298),
    .B(\tholin_riscv.regs[28][23] ),
    .Y(_24349_));
 sky130_as_sc_hs__nand3_2 _30861_ (.A(net168),
    .B(_24348_),
    .C(_24349_),
    .Y(_24350_));
 sky130_as_sc_hs__or2_2 _30863_ (.A(net298),
    .B(\tholin_riscv.regs[30][23] ),
    .Y(_24352_));
 sky130_as_sc_hs__nand3_2 _30864_ (.A(net265),
    .B(_24351_),
    .C(_24352_),
    .Y(_24353_));
 sky130_as_sc_hs__nand3_2 _30865_ (.A(net255),
    .B(_24350_),
    .C(_24353_),
    .Y(_24354_));
 sky130_as_sc_hs__or2_2 _30867_ (.A(net294),
    .B(\tholin_riscv.regs[16][23] ),
    .Y(_24356_));
 sky130_as_sc_hs__nand3_2 _30868_ (.A(net168),
    .B(_24355_),
    .C(_24356_),
    .Y(_24357_));
 sky130_as_sc_hs__or2_2 _30870_ (.A(net294),
    .B(\tholin_riscv.regs[18][23] ),
    .Y(_24359_));
 sky130_as_sc_hs__nand3_2 _30871_ (.A(net265),
    .B(_24358_),
    .C(_24359_),
    .Y(_24360_));
 sky130_as_sc_hs__nand3_2 _30872_ (.A(net161),
    .B(_24357_),
    .C(_24360_),
    .Y(_24361_));
 sky130_as_sc_hs__or2_2 _30874_ (.A(net294),
    .B(\tholin_riscv.regs[22][23] ),
    .Y(_24363_));
 sky130_as_sc_hs__nand3_2 _30875_ (.A(net265),
    .B(_24362_),
    .C(_24363_),
    .Y(_24364_));
 sky130_as_sc_hs__or2_2 _30877_ (.A(net294),
    .B(\tholin_riscv.regs[20][23] ),
    .Y(_24366_));
 sky130_as_sc_hs__nand3_2 _30878_ (.A(net168),
    .B(_24365_),
    .C(_24366_),
    .Y(_24367_));
 sky130_as_sc_hs__nand3_2 _30879_ (.A(net255),
    .B(_24364_),
    .C(_24367_),
    .Y(_24368_));
 sky130_as_sc_hs__nand3_2 _30880_ (.A(net154),
    .B(_24361_),
    .C(_24368_),
    .Y(_24369_));
 sky130_as_sc_hs__nand3_2 _30881_ (.A(net251),
    .B(_24347_),
    .C(_24354_),
    .Y(_24370_));
 sky130_as_sc_hs__nand3_2 _30882_ (.A(net247),
    .B(_24369_),
    .C(_24370_),
    .Y(_24371_));
 sky130_as_sc_hs__or2_2 _30884_ (.A(net300),
    .B(\tholin_riscv.regs[8][23] ),
    .Y(_24373_));
 sky130_as_sc_hs__nand3_2 _30885_ (.A(net170),
    .B(_24372_),
    .C(_24373_),
    .Y(_24374_));
 sky130_as_sc_hs__or2_2 _30887_ (.A(net299),
    .B(\tholin_riscv.regs[10][23] ),
    .Y(_24376_));
 sky130_as_sc_hs__nand3_2 _30888_ (.A(net267),
    .B(_24375_),
    .C(_24376_),
    .Y(_24377_));
 sky130_as_sc_hs__nand3_2 _30889_ (.A(net161),
    .B(_24374_),
    .C(_24377_),
    .Y(_24378_));
 sky130_as_sc_hs__or2_2 _30891_ (.A(net303),
    .B(\tholin_riscv.regs[12][23] ),
    .Y(_24380_));
 sky130_as_sc_hs__nand3_2 _30892_ (.A(net171),
    .B(_24379_),
    .C(_24380_),
    .Y(_24381_));
 sky130_as_sc_hs__or2_2 _30894_ (.A(net303),
    .B(\tholin_riscv.regs[14][23] ),
    .Y(_24383_));
 sky130_as_sc_hs__nand3_2 _30895_ (.A(net268),
    .B(_24382_),
    .C(_24383_),
    .Y(_24384_));
 sky130_as_sc_hs__nand3_2 _30896_ (.A(net256),
    .B(_24381_),
    .C(_24384_),
    .Y(_24385_));
 sky130_as_sc_hs__or2_2 _30898_ (.A(net300),
    .B(\tholin_riscv.regs[0][23] ),
    .Y(_24387_));
 sky130_as_sc_hs__nand3_2 _30899_ (.A(net170),
    .B(_24386_),
    .C(_24387_),
    .Y(_24388_));
 sky130_as_sc_hs__or2_2 _30901_ (.A(net300),
    .B(\tholin_riscv.regs[2][23] ),
    .Y(_24390_));
 sky130_as_sc_hs__nand3_2 _30902_ (.A(net267),
    .B(_24389_),
    .C(_24390_),
    .Y(_24391_));
 sky130_as_sc_hs__nand3_2 _30903_ (.A(net161),
    .B(_24388_),
    .C(_24391_),
    .Y(_24392_));
 sky130_as_sc_hs__or2_2 _30905_ (.A(net300),
    .B(\tholin_riscv.regs[6][23] ),
    .Y(_24394_));
 sky130_as_sc_hs__nand3_2 _30906_ (.A(net267),
    .B(_24393_),
    .C(_24394_),
    .Y(_24395_));
 sky130_as_sc_hs__or2_2 _30908_ (.A(net303),
    .B(\tholin_riscv.regs[4][23] ),
    .Y(_24397_));
 sky130_as_sc_hs__nand3_2 _30909_ (.A(net168),
    .B(_24396_),
    .C(_24397_),
    .Y(_24398_));
 sky130_as_sc_hs__nand3_2 _30910_ (.A(net254),
    .B(_24395_),
    .C(_24398_),
    .Y(_24399_));
 sky130_as_sc_hs__nand3_2 _30911_ (.A(net156),
    .B(_24392_),
    .C(_24399_),
    .Y(_24400_));
 sky130_as_sc_hs__nand3_2 _30912_ (.A(net251),
    .B(_24378_),
    .C(_24385_),
    .Y(_24401_));
 sky130_as_sc_hs__nand3_2 _30913_ (.A(net151),
    .B(_24400_),
    .C(_24401_),
    .Y(_24402_));
 sky130_as_sc_hs__inv_2 _30915_ (.Y(_24404_),
    .A(_24403_));
 sky130_as_sc_hs__and2_2 _30916_ (.A(_24191_),
    .B(_24403_),
    .Y(_24405_));
 sky130_as_sc_hs__nand3_2 _30917_ (.A(_23775_),
    .B(_24116_),
    .C(_24405_),
    .Y(_24406_));
 sky130_as_sc_hs__nor2_2 _30918_ (.A(_24340_),
    .B(_24406_),
    .Y(_24407_));
 sky130_as_sc_hs__or2_2 _30920_ (.A(net197),
    .B(\tholin_riscv.regs[25][24] ),
    .Y(_24409_));
 sky130_as_sc_hs__or2_2 _30921_ (.A(net328),
    .B(\tholin_riscv.regs[24][24] ),
    .Y(_24410_));
 sky130_as_sc_hs__nand3_2 _30922_ (.A(net184),
    .B(_24409_),
    .C(_24410_),
    .Y(_24411_));
 sky130_as_sc_hs__or2_2 _30923_ (.A(net197),
    .B(\tholin_riscv.regs[27][24] ),
    .Y(_24412_));
 sky130_as_sc_hs__or2_2 _30924_ (.A(net328),
    .B(\tholin_riscv.regs[26][24] ),
    .Y(_24413_));
 sky130_as_sc_hs__nand3_2 _30925_ (.A(net279),
    .B(_24412_),
    .C(_24413_),
    .Y(_24414_));
 sky130_as_sc_hs__nand3_2 _30926_ (.A(net163),
    .B(_24411_),
    .C(_24414_),
    .Y(_24415_));
 sky130_as_sc_hs__or2_2 _30927_ (.A(net197),
    .B(\tholin_riscv.regs[29][24] ),
    .Y(_24416_));
 sky130_as_sc_hs__or2_2 _30928_ (.A(net328),
    .B(\tholin_riscv.regs[28][24] ),
    .Y(_24417_));
 sky130_as_sc_hs__nand3_2 _30929_ (.A(net183),
    .B(_24416_),
    .C(_24417_),
    .Y(_24418_));
 sky130_as_sc_hs__or2_2 _30930_ (.A(net197),
    .B(\tholin_riscv.regs[31][24] ),
    .Y(_24419_));
 sky130_as_sc_hs__or2_2 _30931_ (.A(net328),
    .B(\tholin_riscv.regs[30][24] ),
    .Y(_24420_));
 sky130_as_sc_hs__nand3_2 _30932_ (.A(net278),
    .B(_24419_),
    .C(_24420_),
    .Y(_24421_));
 sky130_as_sc_hs__nand3_2 _30933_ (.A(net261),
    .B(_24418_),
    .C(_24421_),
    .Y(_24422_));
 sky130_as_sc_hs__or2_2 _30934_ (.A(net197),
    .B(\tholin_riscv.regs[17][24] ),
    .Y(_24423_));
 sky130_as_sc_hs__or2_2 _30935_ (.A(net319),
    .B(\tholin_riscv.regs[16][24] ),
    .Y(_24424_));
 sky130_as_sc_hs__nand3_2 _30936_ (.A(net183),
    .B(_24423_),
    .C(_24424_),
    .Y(_24425_));
 sky130_as_sc_hs__or2_2 _30937_ (.A(net197),
    .B(\tholin_riscv.regs[19][24] ),
    .Y(_24426_));
 sky130_as_sc_hs__or2_2 _30938_ (.A(net328),
    .B(\tholin_riscv.regs[18][24] ),
    .Y(_24427_));
 sky130_as_sc_hs__nand3_2 _30939_ (.A(net279),
    .B(_24426_),
    .C(_24427_),
    .Y(_24428_));
 sky130_as_sc_hs__nand3_2 _30940_ (.A(net163),
    .B(_24425_),
    .C(_24428_),
    .Y(_24429_));
 sky130_as_sc_hs__or2_2 _30941_ (.A(net197),
    .B(\tholin_riscv.regs[23][24] ),
    .Y(_24430_));
 sky130_as_sc_hs__or2_2 _30942_ (.A(net328),
    .B(\tholin_riscv.regs[22][24] ),
    .Y(_24431_));
 sky130_as_sc_hs__nand3_2 _30943_ (.A(net279),
    .B(_24430_),
    .C(_24431_),
    .Y(_24432_));
 sky130_as_sc_hs__or2_2 _30944_ (.A(net197),
    .B(\tholin_riscv.regs[21][24] ),
    .Y(_24433_));
 sky130_as_sc_hs__or2_2 _30945_ (.A(net328),
    .B(\tholin_riscv.regs[20][24] ),
    .Y(_24434_));
 sky130_as_sc_hs__nand3_2 _30946_ (.A(net183),
    .B(_24433_),
    .C(_24434_),
    .Y(_24435_));
 sky130_as_sc_hs__nand3_2 _30947_ (.A(net261),
    .B(_24432_),
    .C(_24435_),
    .Y(_24436_));
 sky130_as_sc_hs__nand3_2 _30948_ (.A(net155),
    .B(_24429_),
    .C(_24436_),
    .Y(_24437_));
 sky130_as_sc_hs__nand3_2 _30949_ (.A(net252),
    .B(_24415_),
    .C(_24422_),
    .Y(_24438_));
 sky130_as_sc_hs__nand3_2 _30950_ (.A(net247),
    .B(_24437_),
    .C(_24438_),
    .Y(_24439_));
 sky130_as_sc_hs__or2_2 _30951_ (.A(net194),
    .B(\tholin_riscv.regs[9][24] ),
    .Y(_24440_));
 sky130_as_sc_hs__or2_2 _30952_ (.A(net320),
    .B(\tholin_riscv.regs[8][24] ),
    .Y(_24441_));
 sky130_as_sc_hs__nand3_2 _30953_ (.A(net177),
    .B(_24440_),
    .C(_24441_),
    .Y(_24442_));
 sky130_as_sc_hs__or2_2 _30954_ (.A(net193),
    .B(\tholin_riscv.regs[11][24] ),
    .Y(_24443_));
 sky130_as_sc_hs__or2_2 _30955_ (.A(net316),
    .B(\tholin_riscv.regs[10][24] ),
    .Y(_24444_));
 sky130_as_sc_hs__nand3_2 _30956_ (.A(net273),
    .B(_24443_),
    .C(_24444_),
    .Y(_24445_));
 sky130_as_sc_hs__nand3_2 _30957_ (.A(net158),
    .B(_24442_),
    .C(_24445_),
    .Y(_24446_));
 sky130_as_sc_hs__or2_2 _30958_ (.A(net193),
    .B(\tholin_riscv.regs[13][24] ),
    .Y(_24447_));
 sky130_as_sc_hs__or2_2 _30959_ (.A(net316),
    .B(\tholin_riscv.regs[12][24] ),
    .Y(_24448_));
 sky130_as_sc_hs__nand3_2 _30960_ (.A(net179),
    .B(_24447_),
    .C(_24448_),
    .Y(_24449_));
 sky130_as_sc_hs__or2_2 _30961_ (.A(net194),
    .B(\tholin_riscv.regs[15][24] ),
    .Y(_24450_));
 sky130_as_sc_hs__or2_2 _30962_ (.A(net319),
    .B(\tholin_riscv.regs[14][24] ),
    .Y(_24451_));
 sky130_as_sc_hs__nand3_2 _30963_ (.A(net273),
    .B(_24450_),
    .C(_24451_),
    .Y(_24452_));
 sky130_as_sc_hs__nand3_2 _30964_ (.A(net258),
    .B(_24449_),
    .C(_24452_),
    .Y(_24453_));
 sky130_as_sc_hs__or2_2 _30965_ (.A(net192),
    .B(\tholin_riscv.regs[1][24] ),
    .Y(_24454_));
 sky130_as_sc_hs__or2_2 _30966_ (.A(net317),
    .B(\tholin_riscv.regs[0][24] ),
    .Y(_24455_));
 sky130_as_sc_hs__nand3_2 _30967_ (.A(net179),
    .B(_24454_),
    .C(_24455_),
    .Y(_24456_));
 sky130_as_sc_hs__or2_2 _30968_ (.A(net192),
    .B(\tholin_riscv.regs[3][24] ),
    .Y(_24457_));
 sky130_as_sc_hs__or2_2 _30969_ (.A(net317),
    .B(\tholin_riscv.regs[2][24] ),
    .Y(_24458_));
 sky130_as_sc_hs__nand3_2 _30970_ (.A(net272),
    .B(_24457_),
    .C(_24458_),
    .Y(_24459_));
 sky130_as_sc_hs__nand3_2 _30971_ (.A(net158),
    .B(_24456_),
    .C(_24459_),
    .Y(_24460_));
 sky130_as_sc_hs__or2_2 _30972_ (.A(net191),
    .B(\tholin_riscv.regs[7][24] ),
    .Y(_24461_));
 sky130_as_sc_hs__or2_2 _30973_ (.A(net317),
    .B(\tholin_riscv.regs[6][24] ),
    .Y(_24462_));
 sky130_as_sc_hs__nand3_2 _30974_ (.A(net272),
    .B(_24461_),
    .C(_24462_),
    .Y(_24463_));
 sky130_as_sc_hs__or2_2 _30975_ (.A(net192),
    .B(\tholin_riscv.regs[5][24] ),
    .Y(_24464_));
 sky130_as_sc_hs__or2_2 _30976_ (.A(net317),
    .B(\tholin_riscv.regs[4][24] ),
    .Y(_24465_));
 sky130_as_sc_hs__nand3_2 _30977_ (.A(net179),
    .B(_24464_),
    .C(_24465_),
    .Y(_24466_));
 sky130_as_sc_hs__nand3_2 _30978_ (.A(net258),
    .B(_24463_),
    .C(_24466_),
    .Y(_24467_));
 sky130_as_sc_hs__nand3_2 _30979_ (.A(net152),
    .B(_24460_),
    .C(_24467_),
    .Y(_24468_));
 sky130_as_sc_hs__nand3_2 _30980_ (.A(net249),
    .B(_24446_),
    .C(_24453_),
    .Y(_24469_));
 sky130_as_sc_hs__nand3_2 _30981_ (.A(net150),
    .B(_24468_),
    .C(_24469_),
    .Y(_24470_));
 sky130_as_sc_hs__inv_2 _30983_ (.Y(_24472_),
    .A(_24471_));
 sky130_as_sc_hs__nand3_2 _30984_ (.A(_23974_),
    .B(_24407_),
    .C(_24471_),
    .Y(_24473_));
 sky130_as_sc_hs__nor2_2 _30985_ (.A(_24337_),
    .B(_24473_),
    .Y(_24474_));
 sky130_as_sc_hs__and2_2 _30986_ (.A(_24337_),
    .B(_24473_),
    .Y(_24475_));
 sky130_as_sc_hs__or2_2 _30987_ (.A(_24474_),
    .B(_24475_),
    .Y(_24476_));
 sky130_as_sc_hs__and2_2 _30990_ (.A(_24477_),
    .B(_24478_),
    .Y(_24479_));
 sky130_as_sc_hs__and2_2 _30991_ (.A(net112),
    .B(net456),
    .Y(_24480_));
 sky130_as_sc_hs__and2_2 _30992_ (.A(net470),
    .B(_24216_),
    .Y(_24481_));
 sky130_as_sc_hs__nand3_2 _30994_ (.A(_24053_),
    .B(_24196_),
    .C(_24197_),
    .Y(_24483_));
 sky130_as_sc_hs__or2_2 _30996_ (.A(_24482_),
    .B(_24483_),
    .Y(_24485_));
 sky130_as_sc_hs__and2_2 _30997_ (.A(_24484_),
    .B(_24485_),
    .Y(_24486_));
 sky130_as_sc_hs__or2_2 _30999_ (.A(_24481_),
    .B(_24486_),
    .Y(_24488_));
 sky130_as_sc_hs__and2_2 _31000_ (.A(_24487_),
    .B(_24488_),
    .Y(_24489_));
 sky130_as_sc_hs__or2_2 _31002_ (.A(_24480_),
    .B(_24489_),
    .Y(_24491_));
 sky130_as_sc_hs__and2_2 _31003_ (.A(_24490_),
    .B(_24491_),
    .Y(_24492_));
 sky130_as_sc_hs__nor2_2 _31007_ (.A(_22367_),
    .B(_22622_),
    .Y(_24496_));
 sky130_as_sc_hs__or2_2 _31008_ (.A(_22367_),
    .B(_22622_),
    .Y(_24497_));
 sky130_as_sc_hs__or2_2 _31011_ (.A(_21660_),
    .B(_24499_),
    .Y(_24500_));
 sky130_as_sc_hs__and2_2 _31013_ (.A(net460),
    .B(_24501_),
    .Y(_24502_));
 sky130_as_sc_hs__and2_2 _31014_ (.A(net462),
    .B(_24256_),
    .Y(_24503_));
 sky130_as_sc_hs__and2_2 _31015_ (.A(net464),
    .B(_24229_),
    .Y(_24504_));
 sky130_as_sc_hs__or2_2 _31017_ (.A(_24503_),
    .B(_24504_),
    .Y(_24506_));
 sky130_as_sc_hs__and2_2 _31018_ (.A(_24505_),
    .B(_24506_),
    .Y(_24507_));
 sky130_as_sc_hs__or2_2 _31020_ (.A(_24502_),
    .B(_24507_),
    .Y(_24509_));
 sky130_as_sc_hs__and2_2 _31021_ (.A(_24508_),
    .B(_24509_),
    .Y(_24510_));
 sky130_as_sc_hs__or2_2 _31023_ (.A(_24494_),
    .B(_24510_),
    .Y(_24512_));
 sky130_as_sc_hs__and2_2 _31024_ (.A(_24511_),
    .B(_24512_),
    .Y(_24513_));
 sky130_as_sc_hs__or2_2 _31026_ (.A(_24493_),
    .B(_24513_),
    .Y(_24515_));
 sky130_as_sc_hs__and2_2 _31027_ (.A(_24514_),
    .B(_24515_),
    .Y(_24516_));
 sky130_as_sc_hs__or2_2 _31029_ (.A(_24492_),
    .B(_24516_),
    .Y(_24518_));
 sky130_as_sc_hs__or2_2 _31031_ (.A(_24272_),
    .B(_24519_),
    .Y(_24520_));
 sky130_as_sc_hs__and2_2 _31033_ (.A(_24520_),
    .B(_24521_),
    .Y(_24522_));
 sky130_as_sc_hs__or2_2 _31034_ (.A(_23607_),
    .B(_24037_),
    .Y(_24523_));
 sky130_as_sc_hs__or2_2 _31035_ (.A(_23974_),
    .B(_24037_),
    .Y(_24524_));
 sky130_as_sc_hs__and2_2 _31036_ (.A(_24038_),
    .B(_24524_),
    .Y(_24525_));
 sky130_as_sc_hs__and2_2 _31039_ (.A(_24256_),
    .B(_24527_),
    .Y(_24528_));
 sky130_as_sc_hs__nor2_2 _31040_ (.A(_20364_),
    .B(_23619_),
    .Y(_24529_));
 sky130_as_sc_hs__nand3_2 _31042_ (.A(_20449_),
    .B(_20535_),
    .C(_24529_),
    .Y(_24531_));
 sky130_as_sc_hs__nor2_2 _31043_ (.A(_20622_),
    .B(_24531_),
    .Y(_24532_));
 sky130_as_sc_hs__nor2b_2 _31044_ (.A(_24532_),
    .Y(_24533_),
    .B(_20707_));
 sky130_as_sc_hs__or2_2 _31045_ (.A(_23974_),
    .B(_24533_),
    .Y(_24534_));
 sky130_as_sc_hs__or2_2 _31047_ (.A(_20707_),
    .B(_23607_),
    .Y(_24536_));
 sky130_as_sc_hs__and2_2 _31048_ (.A(_24535_),
    .B(_24536_),
    .Y(_24537_));
 sky130_as_sc_hs__nand3_2 _31049_ (.A(_24501_),
    .B(_24535_),
    .C(_24536_),
    .Y(_24538_));
 sky130_as_sc_hs__nand3_2 _31050_ (.A(_24501_),
    .B(_24528_),
    .C(_24537_),
    .Y(_24539_));
 sky130_as_sc_hs__or2_2 _31055_ (.A(_21660_),
    .B(_24543_),
    .Y(_24544_));
 sky130_as_sc_hs__and2_2 _31057_ (.A(_20622_),
    .B(_24531_),
    .Y(_24546_));
 sky130_as_sc_hs__or2_2 _31058_ (.A(_24532_),
    .B(_24546_),
    .Y(_24547_));
 sky130_as_sc_hs__or2_2 _31060_ (.A(_20622_),
    .B(_23607_),
    .Y(_24549_));
 sky130_as_sc_hs__and2_2 _31061_ (.A(_24548_),
    .B(_24549_),
    .Y(_24550_));
 sky130_as_sc_hs__and2_2 _31062_ (.A(_24545_),
    .B(net87),
    .Y(_24551_));
 sky130_as_sc_hs__nand2b_2 _31063_ (.B(_24538_),
    .Y(_24552_),
    .A(_24528_));
 sky130_as_sc_hs__and2_2 _31064_ (.A(_24539_),
    .B(_24552_),
    .Y(_24553_));
 sky130_as_sc_hs__nand3_2 _31067_ (.A(_22494_),
    .B(_22559_),
    .C(_24496_),
    .Y(_24556_));
 sky130_as_sc_hs__and2_2 _31072_ (.A(_24559_),
    .B(_24560_),
    .Y(_24561_));
 sky130_as_sc_hs__and2_2 _31073_ (.A(net87),
    .B(net455),
    .Y(_24562_));
 sky130_as_sc_hs__nand3_2 _31074_ (.A(_24535_),
    .B(_24536_),
    .C(_24545_),
    .Y(_24563_));
 sky130_as_sc_hs__or2_2 _31076_ (.A(_24563_),
    .B(_24564_),
    .Y(_24565_));
 sky130_as_sc_hs__and2_2 _31078_ (.A(_24565_),
    .B(_24566_),
    .Y(_24567_));
 sky130_as_sc_hs__or2_2 _31080_ (.A(_24562_),
    .B(_24567_),
    .Y(_24569_));
 sky130_as_sc_hs__and2_2 _31081_ (.A(_24568_),
    .B(_24569_),
    .Y(_24570_));
 sky130_as_sc_hs__or2_2 _31083_ (.A(_24555_),
    .B(_24570_),
    .Y(_24572_));
 sky130_as_sc_hs__and2_2 _31084_ (.A(_24571_),
    .B(_24572_),
    .Y(_24573_));
 sky130_as_sc_hs__nor2_2 _31085_ (.A(_22430_),
    .B(_24556_),
    .Y(_24574_));
 sky130_as_sc_hs__or2_2 _31087_ (.A(_22879_),
    .B(_24574_),
    .Y(_24576_));
 sky130_as_sc_hs__and2_2 _31091_ (.A(_24578_),
    .B(_24579_),
    .Y(_24580_));
 sky130_as_sc_hs__or2_2 _31092_ (.A(_20449_),
    .B(_24529_),
    .Y(_24581_));
 sky130_as_sc_hs__and2_2 _31096_ (.A(_24583_),
    .B(_24584_),
    .Y(_24585_));
 sky130_as_sc_hs__and2_2 _31097_ (.A(net453),
    .B(net450),
    .Y(_24586_));
 sky130_as_sc_hs__and2_2 _31098_ (.A(_22430_),
    .B(_24556_),
    .Y(_24587_));
 sky130_as_sc_hs__or2_2 _31099_ (.A(_24574_),
    .B(_24587_),
    .Y(_24588_));
 sky130_as_sc_hs__or2_2 _31101_ (.A(_21659_),
    .B(_22430_),
    .Y(_24590_));
 sky130_as_sc_hs__and2_2 _31102_ (.A(_24589_),
    .B(_24590_),
    .Y(_24591_));
 sky130_as_sc_hs__and2_2 _31107_ (.A(_24594_),
    .B(_24595_),
    .Y(_24596_));
 sky130_as_sc_hs__and2_2 _31108_ (.A(net85),
    .B(net448),
    .Y(_24597_));
 sky130_as_sc_hs__or2_2 _31110_ (.A(_24586_),
    .B(_24597_),
    .Y(_24599_));
 sky130_as_sc_hs__and2_2 _31111_ (.A(_24598_),
    .B(_24599_),
    .Y(_24600_));
 sky130_as_sc_hs__and2_2 _31116_ (.A(net87),
    .B(net86),
    .Y(_24605_));
 sky130_as_sc_hs__nand3_2 _31117_ (.A(_24535_),
    .B(_24536_),
    .C(net455),
    .Y(_24606_));
 sky130_as_sc_hs__or2_2 _31119_ (.A(_24606_),
    .B(_24607_),
    .Y(_24608_));
 sky130_as_sc_hs__and2_2 _31121_ (.A(_24608_),
    .B(_24609_),
    .Y(_24610_));
 sky130_as_sc_hs__or2_2 _31123_ (.A(_24605_),
    .B(_24610_),
    .Y(_24612_));
 sky130_as_sc_hs__and2_2 _31124_ (.A(_24611_),
    .B(_24612_),
    .Y(_24613_));
 sky130_as_sc_hs__or2_2 _31126_ (.A(_24604_),
    .B(_24613_),
    .Y(_24615_));
 sky130_as_sc_hs__and2_2 _31127_ (.A(_24614_),
    .B(_24615_),
    .Y(_24616_));
 sky130_as_sc_hs__nand3_2 _31128_ (.A(_22815_),
    .B(_22879_),
    .C(_24574_),
    .Y(_24617_));
 sky130_as_sc_hs__and2_2 _31133_ (.A(_24620_),
    .B(_24621_),
    .Y(_24622_));
 sky130_as_sc_hs__and2_2 _31134_ (.A(net450),
    .B(net447),
    .Y(_24623_));
 sky130_as_sc_hs__and2_2 _31135_ (.A(net453),
    .B(net448),
    .Y(_24624_));
 sky130_as_sc_hs__or2_2 _31137_ (.A(_24623_),
    .B(_24624_),
    .Y(_24626_));
 sky130_as_sc_hs__and2_2 _31138_ (.A(_24625_),
    .B(_24626_),
    .Y(_24627_));
 sky130_as_sc_hs__or2_2 _31140_ (.A(_24616_),
    .B(_24627_),
    .Y(_24629_));
 sky130_as_sc_hs__and2_2 _31141_ (.A(_24628_),
    .B(_24629_),
    .Y(_24630_));
 sky130_as_sc_hs__or2_2 _31143_ (.A(_24603_),
    .B(_24630_),
    .Y(_24632_));
 sky130_as_sc_hs__and2_2 _31144_ (.A(_24631_),
    .B(_24632_),
    .Y(_24633_));
 sky130_as_sc_hs__or2_2 _31146_ (.A(_24602_),
    .B(_24633_),
    .Y(_24635_));
 sky130_as_sc_hs__and2_2 _31147_ (.A(_24634_),
    .B(_24635_),
    .Y(_24636_));
 sky130_as_sc_hs__and2_2 _31150_ (.A(net458),
    .B(net456),
    .Y(_24639_));
 sky130_as_sc_hs__and2_2 _31151_ (.A(net470),
    .B(_24229_),
    .Y(_24640_));
 sky130_as_sc_hs__nand3_2 _31153_ (.A(_23712_),
    .B(_24196_),
    .C(_24197_),
    .Y(_24642_));
 sky130_as_sc_hs__or2_2 _31155_ (.A(_24641_),
    .B(_24642_),
    .Y(_24644_));
 sky130_as_sc_hs__and2_2 _31156_ (.A(_24643_),
    .B(_24644_),
    .Y(_24645_));
 sky130_as_sc_hs__or2_2 _31158_ (.A(_24640_),
    .B(_24645_),
    .Y(_24647_));
 sky130_as_sc_hs__and2_2 _31159_ (.A(_24646_),
    .B(_24647_),
    .Y(_24648_));
 sky130_as_sc_hs__or2_2 _31161_ (.A(_24639_),
    .B(_24648_),
    .Y(_24650_));
 sky130_as_sc_hs__or2_2 _31163_ (.A(_24490_),
    .B(_24651_),
    .Y(_24652_));
 sky130_as_sc_hs__and2_2 _31165_ (.A(_24652_),
    .B(_24653_),
    .Y(_24654_));
 sky130_as_sc_hs__and2_2 _31168_ (.A(net461),
    .B(_24545_),
    .Y(_24657_));
 sky130_as_sc_hs__and2_2 _31169_ (.A(net462),
    .B(_24501_),
    .Y(_24658_));
 sky130_as_sc_hs__and2_2 _31170_ (.A(net464),
    .B(_24256_),
    .Y(_24659_));
 sky130_as_sc_hs__or2_2 _31172_ (.A(_24658_),
    .B(_24659_),
    .Y(_24661_));
 sky130_as_sc_hs__and2_2 _31173_ (.A(_24660_),
    .B(_24661_),
    .Y(_24662_));
 sky130_as_sc_hs__or2_2 _31175_ (.A(_24657_),
    .B(_24662_),
    .Y(_24664_));
 sky130_as_sc_hs__and2_2 _31176_ (.A(_24663_),
    .B(_24664_),
    .Y(_24665_));
 sky130_as_sc_hs__or2_2 _31178_ (.A(_24656_),
    .B(_24665_),
    .Y(_24667_));
 sky130_as_sc_hs__and2_2 _31179_ (.A(_24666_),
    .B(_24667_),
    .Y(_24668_));
 sky130_as_sc_hs__or2_2 _31181_ (.A(_24655_),
    .B(_24668_),
    .Y(_24670_));
 sky130_as_sc_hs__and2_2 _31182_ (.A(_24669_),
    .B(_24670_),
    .Y(_24671_));
 sky130_as_sc_hs__or2_2 _31184_ (.A(_24654_),
    .B(_24671_),
    .Y(_24673_));
 sky130_as_sc_hs__or2_2 _31186_ (.A(_24517_),
    .B(_24674_),
    .Y(_24675_));
 sky130_as_sc_hs__and2_2 _31188_ (.A(_24675_),
    .B(_24676_),
    .Y(_24677_));
 sky130_as_sc_hs__and2_2 _31192_ (.A(net87),
    .B(net453),
    .Y(_24681_));
 sky130_as_sc_hs__nand3_2 _31193_ (.A(_24535_),
    .B(_24536_),
    .C(net86),
    .Y(_24682_));
 sky130_as_sc_hs__or2_2 _31195_ (.A(_24682_),
    .B(_24683_),
    .Y(_24684_));
 sky130_as_sc_hs__and2_2 _31197_ (.A(_24684_),
    .B(_24685_),
    .Y(_24686_));
 sky130_as_sc_hs__or2_2 _31199_ (.A(_24681_),
    .B(_24686_),
    .Y(_24688_));
 sky130_as_sc_hs__and2_2 _31200_ (.A(_24687_),
    .B(_24688_),
    .Y(_24689_));
 sky130_as_sc_hs__or2_2 _31202_ (.A(_24680_),
    .B(_24689_),
    .Y(_24691_));
 sky130_as_sc_hs__and2_2 _31203_ (.A(_24690_),
    .B(_24691_),
    .Y(_24692_));
 sky130_as_sc_hs__or2_2 _31204_ (.A(_22687_),
    .B(_24617_),
    .Y(_24693_));
 sky130_as_sc_hs__or2_2 _31208_ (.A(_21659_),
    .B(_22687_),
    .Y(_24697_));
 sky130_as_sc_hs__and2_2 _31209_ (.A(_24696_),
    .B(_24697_),
    .Y(_24698_));
 sky130_as_sc_hs__and2_2 _31210_ (.A(net450),
    .B(net79),
    .Y(_24699_));
 sky130_as_sc_hs__and2_2 _31211_ (.A(net448),
    .B(net447),
    .Y(_24700_));
 sky130_as_sc_hs__or2_2 _31213_ (.A(_24699_),
    .B(_24700_),
    .Y(_24702_));
 sky130_as_sc_hs__and2_2 _31214_ (.A(_24701_),
    .B(_24702_),
    .Y(_24703_));
 sky130_as_sc_hs__or2_2 _31216_ (.A(_24692_),
    .B(_24703_),
    .Y(_24705_));
 sky130_as_sc_hs__and2_2 _31217_ (.A(_24704_),
    .B(_24705_),
    .Y(_24706_));
 sky130_as_sc_hs__or2_2 _31219_ (.A(_24679_),
    .B(_24706_),
    .Y(_24708_));
 sky130_as_sc_hs__and2_2 _31220_ (.A(_24707_),
    .B(_24708_),
    .Y(_24709_));
 sky130_as_sc_hs__or2_2 _31222_ (.A(_24678_),
    .B(_24709_),
    .Y(_24711_));
 sky130_as_sc_hs__and2_2 _31223_ (.A(_24710_),
    .B(_24711_),
    .Y(_24712_));
 sky130_as_sc_hs__or2_2 _31225_ (.A(_24677_),
    .B(_24712_),
    .Y(_24714_));
 sky130_as_sc_hs__and2_2 _31226_ (.A(_24713_),
    .B(_24714_),
    .Y(_24715_));
 sky130_as_sc_hs__or2_2 _31228_ (.A(_24638_),
    .B(_24715_),
    .Y(_24717_));
 sky130_as_sc_hs__and2_2 _31229_ (.A(_24716_),
    .B(_24717_),
    .Y(_24718_));
 sky130_as_sc_hs__and2_2 _31230_ (.A(_20364_),
    .B(_23619_),
    .Y(_24719_));
 sky130_as_sc_hs__or2_2 _31231_ (.A(_24529_),
    .B(_24719_),
    .Y(_24720_));
 sky130_as_sc_hs__and2_2 _31234_ (.A(_24721_),
    .B(_24722_),
    .Y(_24723_));
 sky130_as_sc_hs__and2_2 _31235_ (.A(net78),
    .B(net444),
    .Y(_24724_));
 sky130_as_sc_hs__or2_2 _31237_ (.A(_20191_),
    .B(_23617_),
    .Y(_24726_));
 sky130_as_sc_hs__nor2b_2 _31238_ (.A(_23618_),
    .Y(_24727_),
    .B(_24726_));
 sky130_as_sc_hs__and2_2 _31241_ (.A(_23674_),
    .B(_24729_),
    .Y(_24730_));
 sky130_as_sc_hs__or2_2 _31243_ (.A(_24724_),
    .B(_24730_),
    .Y(_24732_));
 sky130_as_sc_hs__or2_2 _31245_ (.A(_24598_),
    .B(_24733_),
    .Y(_24734_));
 sky130_as_sc_hs__and2_2 _31248_ (.A(net447),
    .B(net444),
    .Y(_24737_));
 sky130_as_sc_hs__and2_2 _31249_ (.A(_22751_),
    .B(_24693_),
    .Y(_24738_));
 sky130_as_sc_hs__or2_2 _31250_ (.A(_22882_),
    .B(_24738_),
    .Y(_24739_));
 sky130_as_sc_hs__and2_2 _31253_ (.A(_24740_),
    .B(_24741_),
    .Y(_24742_));
 sky130_as_sc_hs__and2_2 _31254_ (.A(_24729_),
    .B(net442),
    .Y(_24743_));
 sky130_as_sc_hs__or2_2 _31256_ (.A(_24736_),
    .B(_24744_),
    .Y(_24745_));
 sky130_as_sc_hs__and2_2 _31258_ (.A(_24745_),
    .B(_24746_),
    .Y(_24747_));
 sky130_as_sc_hs__and2_2 _31259_ (.A(net455),
    .B(net448),
    .Y(_24748_));
 sky130_as_sc_hs__and2_2 _31260_ (.A(net450),
    .B(net86),
    .Y(_24749_));
 sky130_as_sc_hs__or2_2 _31262_ (.A(_24737_),
    .B(_24743_),
    .Y(_24751_));
 sky130_as_sc_hs__or2_2 _31264_ (.A(_24750_),
    .B(_24752_),
    .Y(_24753_));
 sky130_as_sc_hs__and2_2 _31265_ (.A(net78),
    .B(_24729_),
    .Y(_24754_));
 sky130_as_sc_hs__and2_2 _31266_ (.A(net452),
    .B(net444),
    .Y(_24755_));
 sky130_as_sc_hs__or2_2 _31270_ (.A(_24756_),
    .B(_24758_),
    .Y(_24759_));
 sky130_as_sc_hs__or2_2 _31273_ (.A(_24747_),
    .B(_24760_),
    .Y(_24762_));
 sky130_as_sc_hs__and2_2 _31274_ (.A(_24761_),
    .B(_24762_),
    .Y(_24763_));
 sky130_as_sc_hs__and2_2 _31277_ (.A(_23613_),
    .B(_24765_),
    .Y(_24766_));
 sky130_as_sc_hs__and2_2 _31280_ (.A(net473),
    .B(_24768_),
    .Y(_24769_));
 sky130_as_sc_hs__and2_2 _31283_ (.A(_23616_),
    .B(_24771_),
    .Y(_24772_));
 sky130_as_sc_hs__and2_2 _31286_ (.A(net477),
    .B(_24774_),
    .Y(_24775_));
 sky130_as_sc_hs__and2_2 _31291_ (.A(_24778_),
    .B(_24779_),
    .Y(_24780_));
 sky130_as_sc_hs__and2_2 _31292_ (.A(net458),
    .B(net441),
    .Y(_24781_));
 sky130_as_sc_hs__or2_2 _31294_ (.A(_24775_),
    .B(_24781_),
    .Y(_24783_));
 sky130_as_sc_hs__and2_2 _31295_ (.A(_24782_),
    .B(_24783_),
    .Y(_24784_));
 sky130_as_sc_hs__or2_2 _31297_ (.A(_24769_),
    .B(_24784_),
    .Y(_24786_));
 sky130_as_sc_hs__and2_2 _31298_ (.A(_24785_),
    .B(_24786_),
    .Y(_24787_));
 sky130_as_sc_hs__and2_2 _31299_ (.A(net481),
    .B(_24774_),
    .Y(_24788_));
 sky130_as_sc_hs__and2_2 _31300_ (.A(net112),
    .B(net441),
    .Y(_24789_));
 sky130_as_sc_hs__and2_2 _31302_ (.A(_21787_),
    .B(_23012_),
    .Y(_24791_));
 sky130_as_sc_hs__or2_2 _31303_ (.A(_23014_),
    .B(_24791_),
    .Y(_24792_));
 sky130_as_sc_hs__and2_2 _31306_ (.A(_24793_),
    .B(_24794_),
    .Y(_24795_));
 sky130_as_sc_hs__and2_2 _31307_ (.A(_24768_),
    .B(net439),
    .Y(_24796_));
 sky130_as_sc_hs__or2_2 _31308_ (.A(_24788_),
    .B(_24789_),
    .Y(_24797_));
 sky130_as_sc_hs__and2_2 _31309_ (.A(_24790_),
    .B(_24797_),
    .Y(_24798_));
 sky130_as_sc_hs__or2_2 _31313_ (.A(_24787_),
    .B(_24800_),
    .Y(_24802_));
 sky130_as_sc_hs__and2_2 _31314_ (.A(_24801_),
    .B(_24802_),
    .Y(_24803_));
 sky130_as_sc_hs__and2_2 _31316_ (.A(_21140_),
    .B(_23610_),
    .Y(_24805_));
 sky130_as_sc_hs__nor2_2 _31317_ (.A(_23611_),
    .B(_24805_),
    .Y(_24806_));
 sky130_as_sc_hs__and2_2 _31320_ (.A(net475),
    .B(_24808_),
    .Y(_24809_));
 sky130_as_sc_hs__or2_2 _31321_ (.A(_21242_),
    .B(_23607_),
    .Y(_24810_));
 sky130_as_sc_hs__or2_2 _31322_ (.A(_21242_),
    .B(_23611_),
    .Y(_24811_));
 sky130_as_sc_hs__and2_2 _31323_ (.A(_23612_),
    .B(_24811_),
    .Y(_24812_));
 sky130_as_sc_hs__and2_2 _31326_ (.A(net479),
    .B(_24814_),
    .Y(_24815_));
 sky130_as_sc_hs__and2_2 _31331_ (.A(_24818_),
    .B(_24819_),
    .Y(_24820_));
 sky130_as_sc_hs__nand3_2 _31332_ (.A(net91),
    .B(_24818_),
    .C(_24819_),
    .Y(_24821_));
 sky130_as_sc_hs__nand3_2 _31333_ (.A(net90),
    .B(_24815_),
    .C(net437),
    .Y(_24822_));
 sky130_as_sc_hs__nand2b_2 _31334_ (.B(_24821_),
    .Y(_24823_),
    .A(_24815_));
 sky130_as_sc_hs__and2_2 _31335_ (.A(_24822_),
    .B(_24823_),
    .Y(_24824_));
 sky130_as_sc_hs__nand3_2 _31336_ (.A(_24809_),
    .B(_24822_),
    .C(_24823_),
    .Y(_24825_));
 sky130_as_sc_hs__or2_2 _31337_ (.A(_24809_),
    .B(_24824_),
    .Y(_24826_));
 sky130_as_sc_hs__and2_2 _31338_ (.A(_24825_),
    .B(_24826_),
    .Y(_24827_));
 sky130_as_sc_hs__or2_2 _31340_ (.A(_24803_),
    .B(_24827_),
    .Y(_24829_));
 sky130_as_sc_hs__and2_2 _31341_ (.A(_24828_),
    .B(_24829_),
    .Y(_24830_));
 sky130_as_sc_hs__and2_2 _31345_ (.A(net481),
    .B(_24729_),
    .Y(_24834_));
 sky130_as_sc_hs__nand3_2 _31346_ (.A(net445),
    .B(_24740_),
    .C(_24741_),
    .Y(_24835_));
 sky130_as_sc_hs__or2_2 _31347_ (.A(net197),
    .B(\tholin_riscv.regs[25][26] ),
    .Y(_24836_));
 sky130_as_sc_hs__or2_2 _31348_ (.A(net329),
    .B(\tholin_riscv.regs[24][26] ),
    .Y(_24837_));
 sky130_as_sc_hs__nand3_2 _31349_ (.A(net184),
    .B(_24836_),
    .C(_24837_),
    .Y(_24838_));
 sky130_as_sc_hs__or2_2 _31350_ (.A(net197),
    .B(\tholin_riscv.regs[27][26] ),
    .Y(_24839_));
 sky130_as_sc_hs__or2_2 _31351_ (.A(net329),
    .B(\tholin_riscv.regs[26][26] ),
    .Y(_24840_));
 sky130_as_sc_hs__nand3_2 _31352_ (.A(net279),
    .B(_24839_),
    .C(_24840_),
    .Y(_24841_));
 sky130_as_sc_hs__nand3_2 _31353_ (.A(net163),
    .B(_24838_),
    .C(_24841_),
    .Y(_24842_));
 sky130_as_sc_hs__or2_2 _31354_ (.A(net197),
    .B(\tholin_riscv.regs[29][26] ),
    .Y(_24843_));
 sky130_as_sc_hs__or2_2 _31355_ (.A(net329),
    .B(\tholin_riscv.regs[28][26] ),
    .Y(_24844_));
 sky130_as_sc_hs__nand3_2 _31356_ (.A(net184),
    .B(_24843_),
    .C(_24844_),
    .Y(_24845_));
 sky130_as_sc_hs__or2_2 _31357_ (.A(net199),
    .B(\tholin_riscv.regs[31][26] ),
    .Y(_24846_));
 sky130_as_sc_hs__or2_2 _31358_ (.A(net328),
    .B(\tholin_riscv.regs[30][26] ),
    .Y(_24847_));
 sky130_as_sc_hs__nand3_2 _31359_ (.A(net281),
    .B(_24846_),
    .C(_24847_),
    .Y(_24848_));
 sky130_as_sc_hs__nand3_2 _31360_ (.A(net261),
    .B(_24845_),
    .C(_24848_),
    .Y(_24849_));
 sky130_as_sc_hs__or2_2 _31361_ (.A(net199),
    .B(\tholin_riscv.regs[17][26] ),
    .Y(_24850_));
 sky130_as_sc_hs__or2_2 _31362_ (.A(net331),
    .B(\tholin_riscv.regs[16][26] ),
    .Y(_24851_));
 sky130_as_sc_hs__nand3_2 _31363_ (.A(net185),
    .B(_24850_),
    .C(_24851_),
    .Y(_24852_));
 sky130_as_sc_hs__or2_2 _31364_ (.A(net199),
    .B(\tholin_riscv.regs[19][26] ),
    .Y(_24853_));
 sky130_as_sc_hs__or2_2 _31365_ (.A(net331),
    .B(\tholin_riscv.regs[18][26] ),
    .Y(_24854_));
 sky130_as_sc_hs__nand3_2 _31366_ (.A(net281),
    .B(_24853_),
    .C(_24854_),
    .Y(_24855_));
 sky130_as_sc_hs__nand3_2 _31367_ (.A(net164),
    .B(_24852_),
    .C(_24855_),
    .Y(_24856_));
 sky130_as_sc_hs__or2_2 _31368_ (.A(net199),
    .B(\tholin_riscv.regs[23][26] ),
    .Y(_24857_));
 sky130_as_sc_hs__or2_2 _31369_ (.A(net331),
    .B(\tholin_riscv.regs[22][26] ),
    .Y(_24858_));
 sky130_as_sc_hs__nand3_2 _31370_ (.A(net281),
    .B(_24857_),
    .C(_24858_),
    .Y(_24859_));
 sky130_as_sc_hs__or2_2 _31371_ (.A(net199),
    .B(\tholin_riscv.regs[21][26] ),
    .Y(_24860_));
 sky130_as_sc_hs__or2_2 _31372_ (.A(net331),
    .B(\tholin_riscv.regs[20][26] ),
    .Y(_24861_));
 sky130_as_sc_hs__nand3_2 _31373_ (.A(net185),
    .B(_24860_),
    .C(_24861_),
    .Y(_24862_));
 sky130_as_sc_hs__nand3_2 _31374_ (.A(net261),
    .B(_24859_),
    .C(_24862_),
    .Y(_24863_));
 sky130_as_sc_hs__nand3_2 _31375_ (.A(net155),
    .B(_24856_),
    .C(_24863_),
    .Y(_24864_));
 sky130_as_sc_hs__nand3_2 _31376_ (.A(net252),
    .B(_24842_),
    .C(_24849_),
    .Y(_24865_));
 sky130_as_sc_hs__nand3_2 _31377_ (.A(net247),
    .B(_24864_),
    .C(_24865_),
    .Y(_24866_));
 sky130_as_sc_hs__or2_2 _31378_ (.A(net191),
    .B(\tholin_riscv.regs[9][26] ),
    .Y(_24867_));
 sky130_as_sc_hs__or2_2 _31379_ (.A(net316),
    .B(\tholin_riscv.regs[8][26] ),
    .Y(_24868_));
 sky130_as_sc_hs__nand3_2 _31380_ (.A(net179),
    .B(_24867_),
    .C(_24868_),
    .Y(_24869_));
 sky130_as_sc_hs__or2_2 _31381_ (.A(net191),
    .B(\tholin_riscv.regs[11][26] ),
    .Y(_24870_));
 sky130_as_sc_hs__or2_2 _31382_ (.A(net317),
    .B(\tholin_riscv.regs[10][26] ),
    .Y(_24871_));
 sky130_as_sc_hs__nand3_2 _31383_ (.A(net272),
    .B(_24870_),
    .C(_24871_),
    .Y(_24872_));
 sky130_as_sc_hs__nand3_2 _31384_ (.A(net158),
    .B(_24869_),
    .C(_24872_),
    .Y(_24873_));
 sky130_as_sc_hs__or2_2 _31385_ (.A(net192),
    .B(\tholin_riscv.regs[13][26] ),
    .Y(_24874_));
 sky130_as_sc_hs__or2_2 _31386_ (.A(net316),
    .B(\tholin_riscv.regs[12][26] ),
    .Y(_24875_));
 sky130_as_sc_hs__nand3_2 _31387_ (.A(net179),
    .B(_24874_),
    .C(_24875_),
    .Y(_24876_));
 sky130_as_sc_hs__or2_2 _31388_ (.A(net191),
    .B(\tholin_riscv.regs[15][26] ),
    .Y(_24877_));
 sky130_as_sc_hs__or2_2 _31389_ (.A(net317),
    .B(\tholin_riscv.regs[14][26] ),
    .Y(_24878_));
 sky130_as_sc_hs__nand3_2 _31390_ (.A(net272),
    .B(_24877_),
    .C(_24878_),
    .Y(_24879_));
 sky130_as_sc_hs__nand3_2 _31391_ (.A(net258),
    .B(_24876_),
    .C(_24879_),
    .Y(_24880_));
 sky130_as_sc_hs__or2_2 _31392_ (.A(net192),
    .B(\tholin_riscv.regs[1][26] ),
    .Y(_24881_));
 sky130_as_sc_hs__or2_2 _31393_ (.A(net317),
    .B(\tholin_riscv.regs[0][26] ),
    .Y(_24882_));
 sky130_as_sc_hs__nand3_2 _31394_ (.A(net176),
    .B(_24881_),
    .C(_24882_),
    .Y(_24883_));
 sky130_as_sc_hs__or2_2 _31395_ (.A(net192),
    .B(\tholin_riscv.regs[3][26] ),
    .Y(_24884_));
 sky130_as_sc_hs__or2_2 _31396_ (.A(net317),
    .B(\tholin_riscv.regs[2][26] ),
    .Y(_24885_));
 sky130_as_sc_hs__nand3_2 _31397_ (.A(net272),
    .B(_24884_),
    .C(_24885_),
    .Y(_24886_));
 sky130_as_sc_hs__nand3_2 _31398_ (.A(net158),
    .B(_24883_),
    .C(_24886_),
    .Y(_24887_));
 sky130_as_sc_hs__or2_2 _31399_ (.A(net192),
    .B(\tholin_riscv.regs[7][26] ),
    .Y(_24888_));
 sky130_as_sc_hs__or2_2 _31400_ (.A(net317),
    .B(\tholin_riscv.regs[6][26] ),
    .Y(_24889_));
 sky130_as_sc_hs__nand3_2 _31401_ (.A(net272),
    .B(_24888_),
    .C(_24889_),
    .Y(_24890_));
 sky130_as_sc_hs__or2_2 _31402_ (.A(net192),
    .B(\tholin_riscv.regs[5][26] ),
    .Y(_24891_));
 sky130_as_sc_hs__or2_2 _31403_ (.A(net317),
    .B(\tholin_riscv.regs[4][26] ),
    .Y(_24892_));
 sky130_as_sc_hs__nand3_2 _31404_ (.A(net179),
    .B(_24891_),
    .C(_24892_),
    .Y(_24893_));
 sky130_as_sc_hs__nand3_2 _31405_ (.A(net258),
    .B(_24890_),
    .C(_24893_),
    .Y(_24894_));
 sky130_as_sc_hs__nand3_2 _31406_ (.A(net152),
    .B(_24887_),
    .C(_24894_),
    .Y(_24895_));
 sky130_as_sc_hs__nand3_2 _31407_ (.A(net249),
    .B(_24873_),
    .C(_24880_),
    .Y(_24896_));
 sky130_as_sc_hs__nand3_2 _31408_ (.A(net150),
    .B(_24895_),
    .C(_24896_),
    .Y(_24897_));
 sky130_as_sc_hs__or2_2 _31411_ (.A(_24474_),
    .B(_24898_),
    .Y(_24900_));
 sky130_as_sc_hs__and2_2 _31415_ (.A(_24902_),
    .B(_24903_),
    .Y(_24904_));
 sky130_as_sc_hs__or2_2 _31417_ (.A(_24835_),
    .B(_24905_),
    .Y(_24906_));
 sky130_as_sc_hs__and2_2 _31419_ (.A(_24906_),
    .B(_24907_),
    .Y(_24908_));
 sky130_as_sc_hs__or2_2 _31421_ (.A(_24834_),
    .B(_24908_),
    .Y(_24910_));
 sky130_as_sc_hs__or2_2 _31423_ (.A(_24625_),
    .B(_24911_),
    .Y(_24912_));
 sky130_as_sc_hs__or2_2 _31426_ (.A(_24731_),
    .B(_24914_),
    .Y(_24915_));
 sky130_as_sc_hs__and2_2 _31428_ (.A(_24915_),
    .B(_24916_),
    .Y(_24917_));
 sky130_as_sc_hs__or2_2 _31431_ (.A(_24917_),
    .B(_24918_),
    .Y(_24920_));
 sky130_as_sc_hs__and2_2 _31432_ (.A(_24919_),
    .B(_24920_),
    .Y(_24921_));
 sky130_as_sc_hs__and2_2 _31434_ (.A(net479),
    .B(_24768_),
    .Y(_24923_));
 sky130_as_sc_hs__and2_2 _31435_ (.A(_24774_),
    .B(net439),
    .Y(_24924_));
 sky130_as_sc_hs__and2_2 _31436_ (.A(net91),
    .B(net441),
    .Y(_24925_));
 sky130_as_sc_hs__or2_2 _31438_ (.A(_24924_),
    .B(_24925_),
    .Y(_24927_));
 sky130_as_sc_hs__and2_2 _31439_ (.A(_24926_),
    .B(_24927_),
    .Y(_24928_));
 sky130_as_sc_hs__or2_2 _31441_ (.A(_24923_),
    .B(_24928_),
    .Y(_24930_));
 sky130_as_sc_hs__and2_2 _31442_ (.A(_24929_),
    .B(_24930_),
    .Y(_24931_));
 sky130_as_sc_hs__or2_2 _31444_ (.A(_24922_),
    .B(_24931_),
    .Y(_24933_));
 sky130_as_sc_hs__and2_2 _31445_ (.A(_24932_),
    .B(_24933_),
    .Y(_24934_));
 sky130_as_sc_hs__and2_2 _31446_ (.A(_23141_),
    .B(_23652_),
    .Y(_24935_));
 sky130_as_sc_hs__or2_2 _31447_ (.A(_23271_),
    .B(_24935_),
    .Y(_24936_));
 sky130_as_sc_hs__or2_2 _31449_ (.A(_21659_),
    .B(_23141_),
    .Y(_24938_));
 sky130_as_sc_hs__and2_2 _31450_ (.A(_24937_),
    .B(_24938_),
    .Y(_24939_));
 sky130_as_sc_hs__and2_2 _31451_ (.A(_24808_),
    .B(net84),
    .Y(_24940_));
 sky130_as_sc_hs__and2_2 _31452_ (.A(net475),
    .B(_24814_),
    .Y(_24941_));
 sky130_as_sc_hs__nand3_2 _31453_ (.A(_24053_),
    .B(_24818_),
    .C(_24819_),
    .Y(_24942_));
 sky130_as_sc_hs__nand3_2 _31454_ (.A(_24053_),
    .B(net437),
    .C(_24941_),
    .Y(_24943_));
 sky130_as_sc_hs__nand2b_2 _31455_ (.B(_24942_),
    .Y(_24944_),
    .A(_24941_));
 sky130_as_sc_hs__and2_2 _31456_ (.A(_24943_),
    .B(_24944_),
    .Y(_24945_));
 sky130_as_sc_hs__nand3_2 _31457_ (.A(_24940_),
    .B(_24943_),
    .C(_24944_),
    .Y(_24946_));
 sky130_as_sc_hs__or2_2 _31458_ (.A(_24940_),
    .B(_24945_),
    .Y(_24947_));
 sky130_as_sc_hs__and2_2 _31459_ (.A(_24946_),
    .B(_24947_),
    .Y(_24948_));
 sky130_as_sc_hs__or2_2 _31461_ (.A(_24934_),
    .B(_24948_),
    .Y(_24950_));
 sky130_as_sc_hs__and2_2 _31462_ (.A(_24949_),
    .B(_24950_),
    .Y(_24951_));
 sky130_as_sc_hs__or2_2 _31464_ (.A(_24921_),
    .B(_24951_),
    .Y(_24953_));
 sky130_as_sc_hs__and2_2 _31465_ (.A(_24952_),
    .B(_24953_),
    .Y(_24954_));
 sky130_as_sc_hs__or2_2 _31467_ (.A(_24833_),
    .B(_24954_),
    .Y(_24956_));
 sky130_as_sc_hs__and2_2 _31468_ (.A(_24955_),
    .B(_24956_),
    .Y(_24957_));
 sky130_as_sc_hs__or2_2 _31470_ (.A(_24832_),
    .B(_24957_),
    .Y(_24959_));
 sky130_as_sc_hs__and2_2 _31471_ (.A(_24958_),
    .B(_24959_),
    .Y(_24960_));
 sky130_as_sc_hs__or2_2 _31476_ (.A(net200),
    .B(\tholin_riscv.regs[25][27] ),
    .Y(_24965_));
 sky130_as_sc_hs__or2_2 _31477_ (.A(net330),
    .B(\tholin_riscv.regs[24][27] ),
    .Y(_24966_));
 sky130_as_sc_hs__nand3_2 _31478_ (.A(net185),
    .B(_24965_),
    .C(_24966_),
    .Y(_24967_));
 sky130_as_sc_hs__or2_2 _31479_ (.A(net200),
    .B(\tholin_riscv.regs[27][27] ),
    .Y(_24968_));
 sky130_as_sc_hs__or2_2 _31480_ (.A(net330),
    .B(\tholin_riscv.regs[26][27] ),
    .Y(_24969_));
 sky130_as_sc_hs__nand3_2 _31481_ (.A(net280),
    .B(_24968_),
    .C(_24969_),
    .Y(_24970_));
 sky130_as_sc_hs__nand3_2 _31482_ (.A(net164),
    .B(_24967_),
    .C(_24970_),
    .Y(_24971_));
 sky130_as_sc_hs__or2_2 _31483_ (.A(net200),
    .B(\tholin_riscv.regs[29][27] ),
    .Y(_24972_));
 sky130_as_sc_hs__or2_2 _31484_ (.A(net330),
    .B(\tholin_riscv.regs[28][27] ),
    .Y(_24973_));
 sky130_as_sc_hs__nand3_2 _31485_ (.A(net185),
    .B(_24972_),
    .C(_24973_),
    .Y(_24974_));
 sky130_as_sc_hs__or2_2 _31486_ (.A(net200),
    .B(\tholin_riscv.regs[31][27] ),
    .Y(_24975_));
 sky130_as_sc_hs__or2_2 _31487_ (.A(net332),
    .B(\tholin_riscv.regs[30][27] ),
    .Y(_24976_));
 sky130_as_sc_hs__nand3_2 _31488_ (.A(net280),
    .B(_24975_),
    .C(_24976_),
    .Y(_24977_));
 sky130_as_sc_hs__nand3_2 _31489_ (.A(net262),
    .B(_24974_),
    .C(_24977_),
    .Y(_24978_));
 sky130_as_sc_hs__or2_2 _31490_ (.A(net200),
    .B(\tholin_riscv.regs[17][27] ),
    .Y(_24979_));
 sky130_as_sc_hs__or2_2 _31491_ (.A(net330),
    .B(\tholin_riscv.regs[16][27] ),
    .Y(_24980_));
 sky130_as_sc_hs__nand3_2 _31492_ (.A(net185),
    .B(_24979_),
    .C(_24980_),
    .Y(_24981_));
 sky130_as_sc_hs__or2_2 _31493_ (.A(net200),
    .B(\tholin_riscv.regs[19][27] ),
    .Y(_24982_));
 sky130_as_sc_hs__or2_2 _31494_ (.A(net330),
    .B(\tholin_riscv.regs[18][27] ),
    .Y(_24983_));
 sky130_as_sc_hs__nand3_2 _31495_ (.A(net280),
    .B(_24982_),
    .C(_24983_),
    .Y(_24984_));
 sky130_as_sc_hs__nand3_2 _31496_ (.A(net164),
    .B(_24981_),
    .C(_24984_),
    .Y(_24985_));
 sky130_as_sc_hs__or2_2 _31497_ (.A(net200),
    .B(\tholin_riscv.regs[23][27] ),
    .Y(_24986_));
 sky130_as_sc_hs__or2_2 _31498_ (.A(net332),
    .B(\tholin_riscv.regs[22][27] ),
    .Y(_24987_));
 sky130_as_sc_hs__nand3_2 _31499_ (.A(net280),
    .B(_24986_),
    .C(_24987_),
    .Y(_24988_));
 sky130_as_sc_hs__or2_2 _31500_ (.A(net200),
    .B(\tholin_riscv.regs[21][27] ),
    .Y(_24989_));
 sky130_as_sc_hs__or2_2 _31501_ (.A(net332),
    .B(\tholin_riscv.regs[20][27] ),
    .Y(_24990_));
 sky130_as_sc_hs__nand3_2 _31502_ (.A(net185),
    .B(_24989_),
    .C(_24990_),
    .Y(_24991_));
 sky130_as_sc_hs__nand3_2 _31503_ (.A(net262),
    .B(_24988_),
    .C(_24991_),
    .Y(_24992_));
 sky130_as_sc_hs__nand3_2 _31504_ (.A(net155),
    .B(_24985_),
    .C(_24992_),
    .Y(_24993_));
 sky130_as_sc_hs__nand3_2 _31505_ (.A(net252),
    .B(_24971_),
    .C(_24978_),
    .Y(_24994_));
 sky130_as_sc_hs__nand3_2 _31506_ (.A(net248),
    .B(_24993_),
    .C(_24994_),
    .Y(_24995_));
 sky130_as_sc_hs__or2_2 _31507_ (.A(net191),
    .B(\tholin_riscv.regs[9][27] ),
    .Y(_24996_));
 sky130_as_sc_hs__or2_2 _31508_ (.A(net316),
    .B(\tholin_riscv.regs[8][27] ),
    .Y(_24997_));
 sky130_as_sc_hs__nand3_2 _31509_ (.A(net176),
    .B(_24996_),
    .C(_24997_),
    .Y(_24998_));
 sky130_as_sc_hs__or2_2 _31510_ (.A(net191),
    .B(\tholin_riscv.regs[11][27] ),
    .Y(_24999_));
 sky130_as_sc_hs__or2_2 _31511_ (.A(net316),
    .B(\tholin_riscv.regs[10][27] ),
    .Y(_25000_));
 sky130_as_sc_hs__nand3_2 _31512_ (.A(net275),
    .B(_24999_),
    .C(_25000_),
    .Y(_25001_));
 sky130_as_sc_hs__nand3_2 _31513_ (.A(net158),
    .B(_24998_),
    .C(_25001_),
    .Y(_25002_));
 sky130_as_sc_hs__or2_2 _31514_ (.A(net191),
    .B(\tholin_riscv.regs[13][27] ),
    .Y(_25003_));
 sky130_as_sc_hs__or2_2 _31515_ (.A(net316),
    .B(\tholin_riscv.regs[12][27] ),
    .Y(_25004_));
 sky130_as_sc_hs__nand3_2 _31516_ (.A(net176),
    .B(_25003_),
    .C(_25004_),
    .Y(_25005_));
 sky130_as_sc_hs__or2_2 _31517_ (.A(net195),
    .B(\tholin_riscv.regs[15][27] ),
    .Y(_25006_));
 sky130_as_sc_hs__or2_2 _31518_ (.A(net314),
    .B(\tholin_riscv.regs[14][27] ),
    .Y(_25007_));
 sky130_as_sc_hs__nand3_2 _31519_ (.A(net272),
    .B(_25006_),
    .C(_25007_),
    .Y(_25008_));
 sky130_as_sc_hs__nand3_2 _31520_ (.A(net258),
    .B(_25005_),
    .C(_25008_),
    .Y(_25009_));
 sky130_as_sc_hs__or2_2 _31521_ (.A(net191),
    .B(\tholin_riscv.regs[1][27] ),
    .Y(_25010_));
 sky130_as_sc_hs__or2_2 _31522_ (.A(net316),
    .B(\tholin_riscv.regs[0][27] ),
    .Y(_25011_));
 sky130_as_sc_hs__nand3_2 _31523_ (.A(net176),
    .B(_25010_),
    .C(_25011_),
    .Y(_25012_));
 sky130_as_sc_hs__or2_2 _31524_ (.A(net195),
    .B(\tholin_riscv.regs[3][27] ),
    .Y(_25013_));
 sky130_as_sc_hs__or2_2 _31525_ (.A(net314),
    .B(\tholin_riscv.regs[2][27] ),
    .Y(_25014_));
 sky130_as_sc_hs__nand3_2 _31526_ (.A(net272),
    .B(_25013_),
    .C(_25014_),
    .Y(_25015_));
 sky130_as_sc_hs__nand3_2 _31527_ (.A(net158),
    .B(_25012_),
    .C(_25015_),
    .Y(_25016_));
 sky130_as_sc_hs__or2_2 _31528_ (.A(net195),
    .B(\tholin_riscv.regs[7][27] ),
    .Y(_25017_));
 sky130_as_sc_hs__or2_2 _31529_ (.A(net314),
    .B(\tholin_riscv.regs[6][27] ),
    .Y(_25018_));
 sky130_as_sc_hs__nand3_2 _31530_ (.A(net272),
    .B(_25017_),
    .C(_25018_),
    .Y(_25019_));
 sky130_as_sc_hs__or2_2 _31531_ (.A(net195),
    .B(\tholin_riscv.regs[5][27] ),
    .Y(_25020_));
 sky130_as_sc_hs__or2_2 _31532_ (.A(net314),
    .B(\tholin_riscv.regs[4][27] ),
    .Y(_25021_));
 sky130_as_sc_hs__nand3_2 _31533_ (.A(net176),
    .B(_25020_),
    .C(_25021_),
    .Y(_25022_));
 sky130_as_sc_hs__nand3_2 _31534_ (.A(net258),
    .B(_25019_),
    .C(_25022_),
    .Y(_25023_));
 sky130_as_sc_hs__nand3_2 _31535_ (.A(net152),
    .B(_25016_),
    .C(_25023_),
    .Y(_25024_));
 sky130_as_sc_hs__nand3_2 _31536_ (.A(net249),
    .B(_25002_),
    .C(_25009_),
    .Y(_25025_));
 sky130_as_sc_hs__nand3_2 _31537_ (.A(net150),
    .B(_25024_),
    .C(_25025_),
    .Y(_25026_));
 sky130_as_sc_hs__inv_2 _31539_ (.Y(_25028_),
    .A(_25027_));
 sky130_as_sc_hs__and2_2 _31540_ (.A(_24898_),
    .B(_25027_),
    .Y(_25029_));
 sky130_as_sc_hs__and2_2 _31546_ (.A(_25033_),
    .B(_25034_),
    .Y(_25035_));
 sky130_as_sc_hs__and2_2 _31547_ (.A(net112),
    .B(_25035_),
    .Y(_25036_));
 sky130_as_sc_hs__and2_2 _31548_ (.A(net90),
    .B(net456),
    .Y(_25037_));
 sky130_as_sc_hs__or2_2 _31550_ (.A(_25036_),
    .B(_25037_),
    .Y(_25039_));
 sky130_as_sc_hs__and2_2 _31551_ (.A(_25038_),
    .B(_25039_),
    .Y(_25040_));
 sky130_as_sc_hs__and2_2 _31552_ (.A(net470),
    .B(_24256_),
    .Y(_25041_));
 sky130_as_sc_hs__nand3_2 _31553_ (.A(_24196_),
    .B(_24197_),
    .C(_24216_),
    .Y(_25042_));
 sky130_as_sc_hs__or2_2 _31555_ (.A(_25042_),
    .B(_25043_),
    .Y(_25044_));
 sky130_as_sc_hs__and2_2 _31557_ (.A(_25044_),
    .B(_25045_),
    .Y(_25046_));
 sky130_as_sc_hs__or2_2 _31559_ (.A(_25041_),
    .B(_25046_),
    .Y(_25048_));
 sky130_as_sc_hs__and2_2 _31560_ (.A(_25047_),
    .B(_25048_),
    .Y(_25049_));
 sky130_as_sc_hs__or2_2 _31562_ (.A(_25040_),
    .B(_25049_),
    .Y(_25051_));
 sky130_as_sc_hs__or2_2 _31564_ (.A(_24649_),
    .B(_25052_),
    .Y(_25053_));
 sky130_as_sc_hs__and2_2 _31566_ (.A(_25053_),
    .B(_25054_),
    .Y(_25055_));
 sky130_as_sc_hs__and2_2 _31569_ (.A(net461),
    .B(net455),
    .Y(_25058_));
 sky130_as_sc_hs__and2_2 _31570_ (.A(net462),
    .B(_24545_),
    .Y(_25059_));
 sky130_as_sc_hs__and2_2 _31571_ (.A(net464),
    .B(_24501_),
    .Y(_25060_));
 sky130_as_sc_hs__or2_2 _31573_ (.A(_25059_),
    .B(_25060_),
    .Y(_25062_));
 sky130_as_sc_hs__and2_2 _31574_ (.A(_25061_),
    .B(_25062_),
    .Y(_25063_));
 sky130_as_sc_hs__or2_2 _31576_ (.A(_25058_),
    .B(_25063_),
    .Y(_25065_));
 sky130_as_sc_hs__and2_2 _31577_ (.A(_25064_),
    .B(_25065_),
    .Y(_25066_));
 sky130_as_sc_hs__or2_2 _31579_ (.A(_25057_),
    .B(_25066_),
    .Y(_25068_));
 sky130_as_sc_hs__and2_2 _31580_ (.A(_25067_),
    .B(_25068_),
    .Y(_25069_));
 sky130_as_sc_hs__or2_2 _31582_ (.A(_25056_),
    .B(_25069_),
    .Y(_25071_));
 sky130_as_sc_hs__and2_2 _31583_ (.A(_25070_),
    .B(_25071_),
    .Y(_25072_));
 sky130_as_sc_hs__or2_2 _31585_ (.A(_25055_),
    .B(_25072_),
    .Y(_25074_));
 sky130_as_sc_hs__and2_2 _31586_ (.A(_25073_),
    .B(_25074_),
    .Y(_25075_));
 sky130_as_sc_hs__or2_2 _31588_ (.A(_24964_),
    .B(_25075_),
    .Y(_25077_));
 sky130_as_sc_hs__and2_2 _31589_ (.A(_25076_),
    .B(_25077_),
    .Y(_25078_));
 sky130_as_sc_hs__and2_2 _31592_ (.A(_24550_),
    .B(net447),
    .Y(_25081_));
 sky130_as_sc_hs__nand3_2 _31593_ (.A(_24535_),
    .B(_24536_),
    .C(net453),
    .Y(_25082_));
 sky130_as_sc_hs__or2_2 _31595_ (.A(_25082_),
    .B(_25083_),
    .Y(_25084_));
 sky130_as_sc_hs__and2_2 _31597_ (.A(_25084_),
    .B(_25085_),
    .Y(_25086_));
 sky130_as_sc_hs__or2_2 _31599_ (.A(_25081_),
    .B(_25086_),
    .Y(_25088_));
 sky130_as_sc_hs__and2_2 _31600_ (.A(_25087_),
    .B(_25088_),
    .Y(_25089_));
 sky130_as_sc_hs__or2_2 _31603_ (.A(_25089_),
    .B(_25090_),
    .Y(_25092_));
 sky130_as_sc_hs__and2_2 _31604_ (.A(_25091_),
    .B(_25092_),
    .Y(_25093_));
 sky130_as_sc_hs__and2_2 _31605_ (.A(net448),
    .B(net79),
    .Y(_25094_));
 sky130_as_sc_hs__and2_2 _31606_ (.A(net450),
    .B(net443),
    .Y(_25095_));
 sky130_as_sc_hs__or2_2 _31608_ (.A(_25094_),
    .B(_25095_),
    .Y(_25097_));
 sky130_as_sc_hs__and2_2 _31609_ (.A(_25096_),
    .B(_25097_),
    .Y(_25098_));
 sky130_as_sc_hs__or2_2 _31611_ (.A(_25093_),
    .B(_25098_),
    .Y(_25100_));
 sky130_as_sc_hs__and2_2 _31612_ (.A(_25099_),
    .B(_25100_),
    .Y(_25101_));
 sky130_as_sc_hs__or2_2 _31614_ (.A(_25080_),
    .B(_25101_),
    .Y(_25103_));
 sky130_as_sc_hs__and2_2 _31615_ (.A(_25102_),
    .B(_25103_),
    .Y(_25104_));
 sky130_as_sc_hs__or2_2 _31617_ (.A(_25079_),
    .B(_25104_),
    .Y(_25106_));
 sky130_as_sc_hs__and2_2 _31618_ (.A(_25105_),
    .B(_25106_),
    .Y(_25107_));
 sky130_as_sc_hs__or2_2 _31620_ (.A(_25078_),
    .B(_25107_),
    .Y(_25109_));
 sky130_as_sc_hs__and2_2 _31621_ (.A(_25108_),
    .B(_25109_),
    .Y(_25110_));
 sky130_as_sc_hs__or2_2 _31623_ (.A(_24963_),
    .B(_25110_),
    .Y(_25112_));
 sky130_as_sc_hs__and2_2 _31624_ (.A(_25111_),
    .B(_25112_),
    .Y(_25113_));
 sky130_as_sc_hs__and2_2 _31628_ (.A(net477),
    .B(_24729_),
    .Y(_25117_));
 sky130_as_sc_hs__and2_2 _31629_ (.A(_23674_),
    .B(net445),
    .Y(_25118_));
 sky130_as_sc_hs__and2_2 _31630_ (.A(net459),
    .B(net435),
    .Y(_25119_));
 sky130_as_sc_hs__or2_2 _31632_ (.A(_25118_),
    .B(_25119_),
    .Y(_25121_));
 sky130_as_sc_hs__and2_2 _31633_ (.A(_25120_),
    .B(_25121_),
    .Y(_25122_));
 sky130_as_sc_hs__or2_2 _31635_ (.A(_25117_),
    .B(_25122_),
    .Y(_25124_));
 sky130_as_sc_hs__or2_2 _31637_ (.A(_24701_),
    .B(_25125_),
    .Y(_25126_));
 sky130_as_sc_hs__and2_2 _31639_ (.A(_25126_),
    .B(_25127_),
    .Y(_25128_));
 sky130_as_sc_hs__or2_2 _31641_ (.A(_25116_),
    .B(_25128_),
    .Y(_25130_));
 sky130_as_sc_hs__and2_2 _31642_ (.A(_25129_),
    .B(_25130_),
    .Y(_25131_));
 sky130_as_sc_hs__or2_2 _31645_ (.A(_25131_),
    .B(_25132_),
    .Y(_25134_));
 sky130_as_sc_hs__and2_2 _31646_ (.A(_25133_),
    .B(_25134_),
    .Y(_25135_));
 sky130_as_sc_hs__or2_2 _31647_ (.A(_23271_),
    .B(_23525_),
    .Y(_25136_));
 sky130_as_sc_hs__and2_2 _31651_ (.A(_25138_),
    .B(_25139_),
    .Y(_25140_));
 sky130_as_sc_hs__and2_2 _31652_ (.A(_24808_),
    .B(net432),
    .Y(_25141_));
 sky130_as_sc_hs__and2_2 _31653_ (.A(_24814_),
    .B(net84),
    .Y(_25142_));
 sky130_as_sc_hs__nand3_2 _31654_ (.A(_23712_),
    .B(_24818_),
    .C(_24819_),
    .Y(_25143_));
 sky130_as_sc_hs__nand3_2 _31655_ (.A(_23712_),
    .B(net437),
    .C(_25142_),
    .Y(_25144_));
 sky130_as_sc_hs__nand2b_2 _31656_ (.B(_25143_),
    .Y(_25145_),
    .A(_25142_));
 sky130_as_sc_hs__and2_2 _31657_ (.A(_25144_),
    .B(_25145_),
    .Y(_25146_));
 sky130_as_sc_hs__nand3_2 _31658_ (.A(_25141_),
    .B(_25144_),
    .C(_25145_),
    .Y(_25147_));
 sky130_as_sc_hs__or2_2 _31659_ (.A(_25141_),
    .B(_25146_),
    .Y(_25148_));
 sky130_as_sc_hs__and2_2 _31660_ (.A(_25147_),
    .B(_25148_),
    .Y(_25149_));
 sky130_as_sc_hs__and2_2 _31661_ (.A(net475),
    .B(_24768_),
    .Y(_25150_));
 sky130_as_sc_hs__and2_2 _31662_ (.A(net473),
    .B(_24774_),
    .Y(_25151_));
 sky130_as_sc_hs__and2_2 _31663_ (.A(_24053_),
    .B(net441),
    .Y(_25152_));
 sky130_as_sc_hs__or2_2 _31665_ (.A(_25151_),
    .B(_25152_),
    .Y(_25154_));
 sky130_as_sc_hs__and2_2 _31666_ (.A(_25153_),
    .B(_25154_),
    .Y(_25155_));
 sky130_as_sc_hs__or2_2 _31668_ (.A(_25150_),
    .B(_25155_),
    .Y(_25157_));
 sky130_as_sc_hs__and2_2 _31669_ (.A(_25156_),
    .B(_25157_),
    .Y(_25158_));
 sky130_as_sc_hs__or2_2 _31672_ (.A(_25158_),
    .B(_25159_),
    .Y(_25161_));
 sky130_as_sc_hs__and2_2 _31673_ (.A(_25160_),
    .B(_25161_),
    .Y(_25162_));
 sky130_as_sc_hs__or2_2 _31675_ (.A(_25149_),
    .B(_25162_),
    .Y(_25164_));
 sky130_as_sc_hs__and2_2 _31676_ (.A(_25163_),
    .B(_25164_),
    .Y(_25165_));
 sky130_as_sc_hs__or2_2 _31678_ (.A(_25135_),
    .B(_25165_),
    .Y(_25167_));
 sky130_as_sc_hs__and2_2 _31679_ (.A(_25166_),
    .B(_25167_),
    .Y(_25168_));
 sky130_as_sc_hs__or2_2 _31681_ (.A(_25115_),
    .B(_25168_),
    .Y(_25170_));
 sky130_as_sc_hs__and2_2 _31682_ (.A(_25169_),
    .B(_25170_),
    .Y(_25171_));
 sky130_as_sc_hs__or2_2 _31684_ (.A(_25114_),
    .B(_25171_),
    .Y(_25173_));
 sky130_as_sc_hs__and2_2 _31685_ (.A(_25172_),
    .B(_25173_),
    .Y(_25174_));
 sky130_as_sc_hs__or2_2 _31687_ (.A(_25113_),
    .B(_25174_),
    .Y(_25176_));
 sky130_as_sc_hs__and2_2 _31688_ (.A(_25175_),
    .B(_25176_),
    .Y(_25177_));
 sky130_as_sc_hs__or2_2 _31690_ (.A(_24962_),
    .B(_25177_),
    .Y(_25179_));
 sky130_as_sc_hs__and2_2 _31691_ (.A(_25178_),
    .B(_25179_),
    .Y(_25180_));
 sky130_as_sc_hs__and2_2 _31692_ (.A(_23674_),
    .B(_24774_),
    .Y(_25181_));
 sky130_as_sc_hs__and2_2 _31693_ (.A(net477),
    .B(_24768_),
    .Y(_25182_));
 sky130_as_sc_hs__or2_2 _31695_ (.A(_24796_),
    .B(_24798_),
    .Y(_25184_));
 sky130_as_sc_hs__or2_2 _31697_ (.A(_25183_),
    .B(_25185_),
    .Y(_25186_));
 sky130_as_sc_hs__and2_2 _31699_ (.A(_25186_),
    .B(_25187_),
    .Y(_25188_));
 sky130_as_sc_hs__and2_2 _31700_ (.A(net479),
    .B(_24808_),
    .Y(_25189_));
 sky130_as_sc_hs__and2_2 _31701_ (.A(net473),
    .B(_24814_),
    .Y(_25190_));
 sky130_as_sc_hs__nand3_2 _31702_ (.A(net459),
    .B(_24818_),
    .C(_24819_),
    .Y(_25191_));
 sky130_as_sc_hs__nand3_2 _31703_ (.A(net459),
    .B(net437),
    .C(_25190_),
    .Y(_25192_));
 sky130_as_sc_hs__nand2b_2 _31704_ (.B(_25191_),
    .Y(_25193_),
    .A(_25190_));
 sky130_as_sc_hs__and2_2 _31705_ (.A(_25192_),
    .B(_25193_),
    .Y(_25194_));
 sky130_as_sc_hs__or2_2 _31707_ (.A(_25189_),
    .B(_25194_),
    .Y(_25196_));
 sky130_as_sc_hs__and2_2 _31708_ (.A(_25195_),
    .B(_25196_),
    .Y(_25197_));
 sky130_as_sc_hs__and2_2 _31714_ (.A(_23609_),
    .B(_25202_),
    .Y(_25203_));
 sky130_as_sc_hs__and2_2 _31717_ (.A(net432),
    .B(_25205_),
    .Y(_25206_));
 sky130_as_sc_hs__and2_2 _31720_ (.A(_23610_),
    .B(_25208_),
    .Y(_25209_));
 sky130_as_sc_hs__and2_2 _31723_ (.A(net84),
    .B(_25211_),
    .Y(_25212_));
 sky130_as_sc_hs__or2_2 _31725_ (.A(_25206_),
    .B(_25212_),
    .Y(_25214_));
 sky130_as_sc_hs__and2_2 _31726_ (.A(_25213_),
    .B(_25214_),
    .Y(_25215_));
 sky130_as_sc_hs__or2_2 _31728_ (.A(_25200_),
    .B(_25215_),
    .Y(_25217_));
 sky130_as_sc_hs__and2_2 _31730_ (.A(net84),
    .B(_25205_),
    .Y(_25219_));
 sky130_as_sc_hs__and2_2 _31731_ (.A(net475),
    .B(_25211_),
    .Y(_25220_));
 sky130_as_sc_hs__or2_2 _31733_ (.A(_25218_),
    .B(_25221_),
    .Y(_25222_));
 sky130_as_sc_hs__and2_2 _31735_ (.A(_25222_),
    .B(_25223_),
    .Y(_25224_));
 sky130_as_sc_hs__and2_2 _31737_ (.A(net439),
    .B(_24814_),
    .Y(_25226_));
 sky130_as_sc_hs__nand3_2 _31738_ (.A(net112),
    .B(_24818_),
    .C(_24819_),
    .Y(_25227_));
 sky130_as_sc_hs__nand3_2 _31739_ (.A(net112),
    .B(net437),
    .C(_25226_),
    .Y(_25228_));
 sky130_as_sc_hs__and2_2 _31740_ (.A(net473),
    .B(_24808_),
    .Y(_25229_));
 sky130_as_sc_hs__nand2b_2 _31741_ (.B(_25227_),
    .Y(_25230_),
    .A(_25226_));
 sky130_as_sc_hs__and2_2 _31742_ (.A(_25228_),
    .B(_25230_),
    .Y(_25231_));
 sky130_as_sc_hs__or2_2 _31745_ (.A(_25219_),
    .B(_25220_),
    .Y(_25234_));
 sky130_as_sc_hs__and2_2 _31746_ (.A(_25221_),
    .B(_25234_),
    .Y(_25235_));
 sky130_as_sc_hs__and2_2 _31748_ (.A(net479),
    .B(_25211_),
    .Y(_25237_));
 sky130_as_sc_hs__and2_2 _31749_ (.A(net475),
    .B(_25205_),
    .Y(_25238_));
 sky130_as_sc_hs__or2_2 _31751_ (.A(_25233_),
    .B(_25235_),
    .Y(_25240_));
 sky130_as_sc_hs__or2_2 _31753_ (.A(_25239_),
    .B(_25241_),
    .Y(_25242_));
 sky130_as_sc_hs__or2_2 _31755_ (.A(_25199_),
    .B(_25224_),
    .Y(_25244_));
 sky130_as_sc_hs__and2_2 _31756_ (.A(_25225_),
    .B(_25244_),
    .Y(_25245_));
 sky130_as_sc_hs__nand3_2 _31757_ (.A(_25225_),
    .B(_25243_),
    .C(_25244_),
    .Y(_25246_));
 sky130_as_sc_hs__and2_2 _31766_ (.A(_25253_),
    .B(_25254_),
    .Y(_25255_));
 sky130_as_sc_hs__and2_2 _31767_ (.A(_25205_),
    .B(net430),
    .Y(_25256_));
 sky130_as_sc_hs__and2_2 _31768_ (.A(net432),
    .B(_25211_),
    .Y(_25257_));
 sky130_as_sc_hs__or2_2 _31770_ (.A(_25256_),
    .B(_25257_),
    .Y(_25259_));
 sky130_as_sc_hs__and2_2 _31771_ (.A(_25258_),
    .B(_25259_),
    .Y(_25260_));
 sky130_as_sc_hs__or2_2 _31773_ (.A(_25250_),
    .B(_25260_),
    .Y(_25262_));
 sky130_as_sc_hs__or2_2 _31775_ (.A(_25213_),
    .B(_25263_),
    .Y(_25264_));
 sky130_as_sc_hs__and2_2 _31777_ (.A(_25264_),
    .B(_25265_),
    .Y(_25266_));
 sky130_as_sc_hs__or2_2 _31779_ (.A(_25249_),
    .B(_25266_),
    .Y(_25268_));
 sky130_as_sc_hs__and2_2 _31780_ (.A(_25267_),
    .B(_25268_),
    .Y(_25269_));
 sky130_as_sc_hs__or2_2 _31782_ (.A(_25248_),
    .B(_25269_),
    .Y(_25271_));
 sky130_as_sc_hs__and2_2 _31783_ (.A(_25270_),
    .B(_25271_),
    .Y(_25272_));
 sky130_as_sc_hs__or2_2 _31785_ (.A(_25247_),
    .B(_25272_),
    .Y(_25274_));
 sky130_as_sc_hs__and2_2 _31786_ (.A(_25273_),
    .B(_25274_),
    .Y(_25275_));
 sky130_as_sc_hs__and2_2 _31787_ (.A(net477),
    .B(_23702_),
    .Y(_25276_));
 sky130_as_sc_hs__and2_2 _31792_ (.A(_25279_),
    .B(_25280_),
    .Y(_25281_));
 sky130_as_sc_hs__and2_2 _31793_ (.A(net114),
    .B(net428),
    .Y(_25282_));
 sky130_as_sc_hs__or2_2 _31794_ (.A(_23675_),
    .B(_23681_),
    .Y(_25283_));
 sky130_as_sc_hs__and2_2 _31796_ (.A(net482),
    .B(net442),
    .Y(_25285_));
 sky130_as_sc_hs__and2_2 _31797_ (.A(_23636_),
    .B(net438),
    .Y(_25286_));
 sky130_as_sc_hs__or2_2 _31799_ (.A(_25284_),
    .B(_25287_),
    .Y(_25288_));
 sky130_as_sc_hs__and2_2 _31801_ (.A(_25288_),
    .B(_25289_),
    .Y(_25290_));
 sky130_as_sc_hs__or2_2 _31803_ (.A(_25282_),
    .B(_25290_),
    .Y(_25292_));
 sky130_as_sc_hs__and2_2 _31804_ (.A(_25291_),
    .B(_25292_),
    .Y(_25293_));
 sky130_as_sc_hs__or2_2 _31805_ (.A(_25285_),
    .B(_25286_),
    .Y(_25294_));
 sky130_as_sc_hs__and2_2 _31807_ (.A(_23636_),
    .B(net476),
    .Y(_25296_));
 sky130_as_sc_hs__and2_2 _31808_ (.A(net482),
    .B(net78),
    .Y(_25297_));
 sky130_as_sc_hs__or2_2 _31810_ (.A(_25295_),
    .B(_25298_),
    .Y(_25299_));
 sky130_as_sc_hs__and2_2 _31811_ (.A(net115),
    .B(net430),
    .Y(_25300_));
 sky130_as_sc_hs__and2_2 _31813_ (.A(_25299_),
    .B(_25301_),
    .Y(_25302_));
 sky130_as_sc_hs__or2_2 _31817_ (.A(_25293_),
    .B(_25304_),
    .Y(_25306_));
 sky130_as_sc_hs__and2_2 _31818_ (.A(_25305_),
    .B(_25306_),
    .Y(_25307_));
 sky130_as_sc_hs__or2_2 _31820_ (.A(_25276_),
    .B(_25307_),
    .Y(_25309_));
 sky130_as_sc_hs__and2_2 _31821_ (.A(_25308_),
    .B(_25309_),
    .Y(_25310_));
 sky130_as_sc_hs__and2_2 _31829_ (.A(_25205_),
    .B(net428),
    .Y(_25318_));
 sky130_as_sc_hs__and2_2 _31830_ (.A(_25211_),
    .B(net430),
    .Y(_25319_));
 sky130_as_sc_hs__or2_2 _31832_ (.A(_25318_),
    .B(_25319_),
    .Y(_25321_));
 sky130_as_sc_hs__and2_2 _31833_ (.A(_25320_),
    .B(_25321_),
    .Y(_25322_));
 sky130_as_sc_hs__or2_2 _31835_ (.A(_25317_),
    .B(_25322_),
    .Y(_25324_));
 sky130_as_sc_hs__or2_2 _31837_ (.A(_25258_),
    .B(_25325_),
    .Y(_25326_));
 sky130_as_sc_hs__and2_2 _31839_ (.A(_25326_),
    .B(_25327_),
    .Y(_25328_));
 sky130_as_sc_hs__or2_2 _31841_ (.A(_25316_),
    .B(_25328_),
    .Y(_25330_));
 sky130_as_sc_hs__and2_2 _31842_ (.A(_25329_),
    .B(_25330_),
    .Y(_25331_));
 sky130_as_sc_hs__or2_2 _31844_ (.A(_25315_),
    .B(_25331_),
    .Y(_25333_));
 sky130_as_sc_hs__and2_2 _31845_ (.A(_25332_),
    .B(_25333_),
    .Y(_25334_));
 sky130_as_sc_hs__or2_2 _31847_ (.A(_25314_),
    .B(_25334_),
    .Y(_25336_));
 sky130_as_sc_hs__and2_2 _31848_ (.A(_25335_),
    .B(_25336_),
    .Y(_25337_));
 sky130_as_sc_hs__and2_2 _31849_ (.A(_23702_),
    .B(net439),
    .Y(_25338_));
 sky130_as_sc_hs__or2_2 _31850_ (.A(_23692_),
    .B(_23694_),
    .Y(_25339_));
 sky130_as_sc_hs__and2_2 _31851_ (.A(_23695_),
    .B(_25339_),
    .Y(_25340_));
 sky130_as_sc_hs__or2_2 _31854_ (.A(_25340_),
    .B(_25341_),
    .Y(_25343_));
 sky130_as_sc_hs__and2_2 _31855_ (.A(_25342_),
    .B(_25343_),
    .Y(_25344_));
 sky130_as_sc_hs__or2_2 _31857_ (.A(_25338_),
    .B(_25344_),
    .Y(_25346_));
 sky130_as_sc_hs__and2_2 _31858_ (.A(_25345_),
    .B(_25346_),
    .Y(_25347_));
 sky130_as_sc_hs__or2_2 _31860_ (.A(_25337_),
    .B(_25347_),
    .Y(_25349_));
 sky130_as_sc_hs__and2_2 _31861_ (.A(_25348_),
    .B(_25349_),
    .Y(_25350_));
 sky130_as_sc_hs__or2_2 _31863_ (.A(_25313_),
    .B(_25350_),
    .Y(_25352_));
 sky130_as_sc_hs__and2_2 _31864_ (.A(_25351_),
    .B(_25352_),
    .Y(_25353_));
 sky130_as_sc_hs__or2_2 _31866_ (.A(_25312_),
    .B(_25353_),
    .Y(_25355_));
 sky130_as_sc_hs__and2_2 _31867_ (.A(_25354_),
    .B(_25355_),
    .Y(_25356_));
 sky130_as_sc_hs__and2_2 _31873_ (.A(net458),
    .B(_25035_),
    .Y(_25362_));
 sky130_as_sc_hs__and2_2 _31874_ (.A(_24053_),
    .B(net456),
    .Y(_25363_));
 sky130_as_sc_hs__or2_2 _31876_ (.A(_25362_),
    .B(_25363_),
    .Y(_25365_));
 sky130_as_sc_hs__or2_2 _31878_ (.A(_25038_),
    .B(_25366_),
    .Y(_25367_));
 sky130_as_sc_hs__and2_2 _31880_ (.A(_25367_),
    .B(_25368_),
    .Y(_25369_));
 sky130_as_sc_hs__and2_2 _31881_ (.A(net470),
    .B(_24501_),
    .Y(_25370_));
 sky130_as_sc_hs__nand3_2 _31882_ (.A(_24196_),
    .B(_24197_),
    .C(_24229_),
    .Y(_25371_));
 sky130_as_sc_hs__or2_2 _31884_ (.A(_25371_),
    .B(_25372_),
    .Y(_25373_));
 sky130_as_sc_hs__and2_2 _31886_ (.A(_25373_),
    .B(_25374_),
    .Y(_25375_));
 sky130_as_sc_hs__or2_2 _31888_ (.A(_25370_),
    .B(_25375_),
    .Y(_25377_));
 sky130_as_sc_hs__and2_2 _31889_ (.A(_25376_),
    .B(_25377_),
    .Y(_25378_));
 sky130_as_sc_hs__or2_2 _31891_ (.A(_25369_),
    .B(_25378_),
    .Y(_25380_));
 sky130_as_sc_hs__or2_2 _31893_ (.A(_25050_),
    .B(_25381_),
    .Y(_25382_));
 sky130_as_sc_hs__and2_2 _31895_ (.A(_25382_),
    .B(_25383_),
    .Y(_25384_));
 sky130_as_sc_hs__and2_2 _31898_ (.A(net461),
    .B(net86),
    .Y(_25387_));
 sky130_as_sc_hs__and2_2 _31899_ (.A(net464),
    .B(_24545_),
    .Y(_25388_));
 sky130_as_sc_hs__and2_2 _31900_ (.A(net462),
    .B(net455),
    .Y(_25389_));
 sky130_as_sc_hs__or2_2 _31901_ (.A(_25388_),
    .B(_25389_),
    .Y(_25390_));
 sky130_as_sc_hs__and2_2 _31903_ (.A(_25390_),
    .B(_25391_),
    .Y(_25392_));
 sky130_as_sc_hs__or2_2 _31905_ (.A(_25387_),
    .B(_25392_),
    .Y(_25394_));
 sky130_as_sc_hs__and2_2 _31906_ (.A(_25393_),
    .B(_25394_),
    .Y(_25395_));
 sky130_as_sc_hs__or2_2 _31908_ (.A(_25386_),
    .B(_25395_),
    .Y(_25397_));
 sky130_as_sc_hs__and2_2 _31909_ (.A(_25396_),
    .B(_25397_),
    .Y(_25398_));
 sky130_as_sc_hs__or2_2 _31911_ (.A(_25385_),
    .B(_25398_),
    .Y(_25400_));
 sky130_as_sc_hs__and2_2 _31912_ (.A(_25399_),
    .B(_25400_),
    .Y(_25401_));
 sky130_as_sc_hs__or2_2 _31914_ (.A(_25384_),
    .B(_25401_),
    .Y(_25403_));
 sky130_as_sc_hs__and2_2 _31915_ (.A(_25402_),
    .B(_25403_),
    .Y(_25404_));
 sky130_as_sc_hs__or2_2 _31917_ (.A(_25361_),
    .B(_25404_),
    .Y(_25406_));
 sky130_as_sc_hs__and2_2 _31918_ (.A(_25405_),
    .B(_25406_),
    .Y(_25407_));
 sky130_as_sc_hs__and2_2 _31921_ (.A(net87),
    .B(net79),
    .Y(_25410_));
 sky130_as_sc_hs__nand3_2 _31922_ (.A(_24535_),
    .B(_24536_),
    .C(net447),
    .Y(_25411_));
 sky130_as_sc_hs__or2_2 _31924_ (.A(_25411_),
    .B(_25412_),
    .Y(_25413_));
 sky130_as_sc_hs__and2_2 _31926_ (.A(_25413_),
    .B(_25414_),
    .Y(_25415_));
 sky130_as_sc_hs__or2_2 _31928_ (.A(_25410_),
    .B(_25415_),
    .Y(_25417_));
 sky130_as_sc_hs__and2_2 _31929_ (.A(_25416_),
    .B(_25417_),
    .Y(_25418_));
 sky130_as_sc_hs__or2_2 _31932_ (.A(_25418_),
    .B(_25419_),
    .Y(_25421_));
 sky130_as_sc_hs__and2_2 _31933_ (.A(_25420_),
    .B(_25421_),
    .Y(_25422_));
 sky130_as_sc_hs__and2_2 _31934_ (.A(_23674_),
    .B(net450),
    .Y(_25423_));
 sky130_as_sc_hs__nand3_2 _31935_ (.A(net449),
    .B(_24740_),
    .C(_24741_),
    .Y(_25424_));
 sky130_as_sc_hs__or2_2 _31936_ (.A(net200),
    .B(\tholin_riscv.regs[25][28] ),
    .Y(_25425_));
 sky130_as_sc_hs__or2_2 _31937_ (.A(net331),
    .B(\tholin_riscv.regs[24][28] ),
    .Y(_25426_));
 sky130_as_sc_hs__nand3_2 _31938_ (.A(net186),
    .B(_25425_),
    .C(_25426_),
    .Y(_25427_));
 sky130_as_sc_hs__or2_2 _31939_ (.A(net199),
    .B(\tholin_riscv.regs[27][28] ),
    .Y(_25428_));
 sky130_as_sc_hs__or2_2 _31940_ (.A(net331),
    .B(\tholin_riscv.regs[26][28] ),
    .Y(_25429_));
 sky130_as_sc_hs__nand3_2 _31941_ (.A(net280),
    .B(_25428_),
    .C(_25429_),
    .Y(_25430_));
 sky130_as_sc_hs__nand3_2 _31942_ (.A(net164),
    .B(_25427_),
    .C(_25430_),
    .Y(_25431_));
 sky130_as_sc_hs__or2_2 _31943_ (.A(net199),
    .B(\tholin_riscv.regs[29][28] ),
    .Y(_25432_));
 sky130_as_sc_hs__or2_2 _31944_ (.A(net331),
    .B(\tholin_riscv.regs[28][28] ),
    .Y(_25433_));
 sky130_as_sc_hs__nand3_2 _31945_ (.A(net185),
    .B(_25432_),
    .C(_25433_),
    .Y(_25434_));
 sky130_as_sc_hs__or2_2 _31946_ (.A(net199),
    .B(\tholin_riscv.regs[31][28] ),
    .Y(_25435_));
 sky130_as_sc_hs__or2_2 _31947_ (.A(net331),
    .B(\tholin_riscv.regs[30][28] ),
    .Y(_25436_));
 sky130_as_sc_hs__nand3_2 _31948_ (.A(net280),
    .B(_25435_),
    .C(_25436_),
    .Y(_25437_));
 sky130_as_sc_hs__nand3_2 _31949_ (.A(net262),
    .B(_25434_),
    .C(_25437_),
    .Y(_25438_));
 sky130_as_sc_hs__or2_2 _31950_ (.A(net199),
    .B(\tholin_riscv.regs[17][28] ),
    .Y(_25439_));
 sky130_as_sc_hs__or2_2 _31951_ (.A(net331),
    .B(\tholin_riscv.regs[16][28] ),
    .Y(_25440_));
 sky130_as_sc_hs__nand3_2 _31952_ (.A(net185),
    .B(_25439_),
    .C(_25440_),
    .Y(_25441_));
 sky130_as_sc_hs__or2_2 _31953_ (.A(net199),
    .B(\tholin_riscv.regs[19][28] ),
    .Y(_25442_));
 sky130_as_sc_hs__or2_2 _31954_ (.A(net331),
    .B(\tholin_riscv.regs[18][28] ),
    .Y(_25443_));
 sky130_as_sc_hs__nand3_2 _31955_ (.A(net280),
    .B(_25442_),
    .C(_25443_),
    .Y(_25444_));
 sky130_as_sc_hs__nand3_2 _31956_ (.A(net165),
    .B(_25441_),
    .C(_25444_),
    .Y(_25445_));
 sky130_as_sc_hs__or2_2 _31957_ (.A(net199),
    .B(\tholin_riscv.regs[23][28] ),
    .Y(_25446_));
 sky130_as_sc_hs__or2_2 _31958_ (.A(net331),
    .B(\tholin_riscv.regs[22][28] ),
    .Y(_25447_));
 sky130_as_sc_hs__nand3_2 _31959_ (.A(net280),
    .B(_25446_),
    .C(_25447_),
    .Y(_25448_));
 sky130_as_sc_hs__or2_2 _31960_ (.A(net199),
    .B(\tholin_riscv.regs[21][28] ),
    .Y(_25449_));
 sky130_as_sc_hs__or2_2 _31961_ (.A(net330),
    .B(\tholin_riscv.regs[20][28] ),
    .Y(_25450_));
 sky130_as_sc_hs__nand3_2 _31962_ (.A(net185),
    .B(_25449_),
    .C(_25450_),
    .Y(_25451_));
 sky130_as_sc_hs__nand3_2 _31963_ (.A(net262),
    .B(_25448_),
    .C(_25451_),
    .Y(_25452_));
 sky130_as_sc_hs__nand3_2 _31964_ (.A(net155),
    .B(_25445_),
    .C(_25452_),
    .Y(_25453_));
 sky130_as_sc_hs__nand3_2 _31965_ (.A(net252),
    .B(_25431_),
    .C(_25438_),
    .Y(_25454_));
 sky130_as_sc_hs__nand3_2 _31966_ (.A(_00004_),
    .B(_25453_),
    .C(_25454_),
    .Y(_25455_));
 sky130_as_sc_hs__or2_2 _31967_ (.A(net191),
    .B(\tholin_riscv.regs[9][28] ),
    .Y(_25456_));
 sky130_as_sc_hs__or2_2 _31968_ (.A(net316),
    .B(\tholin_riscv.regs[8][28] ),
    .Y(_25457_));
 sky130_as_sc_hs__nand3_2 _31969_ (.A(net176),
    .B(_25456_),
    .C(_25457_),
    .Y(_25458_));
 sky130_as_sc_hs__or2_2 _31970_ (.A(net191),
    .B(\tholin_riscv.regs[11][28] ),
    .Y(_25459_));
 sky130_as_sc_hs__or2_2 _31971_ (.A(net316),
    .B(\tholin_riscv.regs[10][28] ),
    .Y(_25460_));
 sky130_as_sc_hs__nand3_2 _31972_ (.A(net275),
    .B(_25459_),
    .C(_25460_),
    .Y(_25461_));
 sky130_as_sc_hs__nand3_2 _31973_ (.A(net158),
    .B(_25458_),
    .C(_25461_),
    .Y(_25462_));
 sky130_as_sc_hs__or2_2 _31974_ (.A(net191),
    .B(\tholin_riscv.regs[13][28] ),
    .Y(_25463_));
 sky130_as_sc_hs__or2_2 _31975_ (.A(net316),
    .B(\tholin_riscv.regs[12][28] ),
    .Y(_25464_));
 sky130_as_sc_hs__nand3_2 _31976_ (.A(net176),
    .B(_25463_),
    .C(_25464_),
    .Y(_25465_));
 sky130_as_sc_hs__or2_2 _31977_ (.A(net191),
    .B(\tholin_riscv.regs[15][28] ),
    .Y(_25466_));
 sky130_as_sc_hs__or2_2 _31978_ (.A(net316),
    .B(\tholin_riscv.regs[14][28] ),
    .Y(_25467_));
 sky130_as_sc_hs__nand3_2 _31979_ (.A(net275),
    .B(_25466_),
    .C(_25467_),
    .Y(_25468_));
 sky130_as_sc_hs__nand3_2 _31980_ (.A(net258),
    .B(_25465_),
    .C(_25468_),
    .Y(_25469_));
 sky130_as_sc_hs__or2_2 _31981_ (.A(net191),
    .B(\tholin_riscv.regs[1][28] ),
    .Y(_25470_));
 sky130_as_sc_hs__or2_2 _31982_ (.A(net316),
    .B(\tholin_riscv.regs[0][28] ),
    .Y(_25471_));
 sky130_as_sc_hs__nand3_2 _31983_ (.A(net176),
    .B(_25470_),
    .C(_25471_),
    .Y(_25472_));
 sky130_as_sc_hs__or2_2 _31984_ (.A(net191),
    .B(\tholin_riscv.regs[3][28] ),
    .Y(_25473_));
 sky130_as_sc_hs__or2_2 _31985_ (.A(net316),
    .B(\tholin_riscv.regs[2][28] ),
    .Y(_25474_));
 sky130_as_sc_hs__nand3_2 _31986_ (.A(net275),
    .B(_25473_),
    .C(_25474_),
    .Y(_25475_));
 sky130_as_sc_hs__nand3_2 _31987_ (.A(net158),
    .B(_25472_),
    .C(_25475_),
    .Y(_25476_));
 sky130_as_sc_hs__or2_2 _31988_ (.A(net191),
    .B(\tholin_riscv.regs[7][28] ),
    .Y(_25477_));
 sky130_as_sc_hs__or2_2 _31989_ (.A(net316),
    .B(\tholin_riscv.regs[6][28] ),
    .Y(_25478_));
 sky130_as_sc_hs__nand3_2 _31990_ (.A(net275),
    .B(_25477_),
    .C(_25478_),
    .Y(_25479_));
 sky130_as_sc_hs__or2_2 _31991_ (.A(net191),
    .B(\tholin_riscv.regs[5][28] ),
    .Y(_25480_));
 sky130_as_sc_hs__or2_2 _31992_ (.A(net316),
    .B(\tholin_riscv.regs[4][28] ),
    .Y(_25481_));
 sky130_as_sc_hs__nand3_2 _31993_ (.A(net176),
    .B(_25480_),
    .C(_25481_),
    .Y(_25482_));
 sky130_as_sc_hs__nand3_2 _31994_ (.A(net258),
    .B(_25479_),
    .C(_25482_),
    .Y(_25483_));
 sky130_as_sc_hs__nand3_2 _31995_ (.A(net152),
    .B(_25476_),
    .C(_25483_),
    .Y(_25484_));
 sky130_as_sc_hs__nand3_2 _31996_ (.A(net249),
    .B(_25462_),
    .C(_25469_),
    .Y(_25485_));
 sky130_as_sc_hs__nand3_2 _31997_ (.A(net150),
    .B(_25484_),
    .C(_25485_),
    .Y(_25486_));
 sky130_as_sc_hs__inv_2 _31999_ (.Y(_25488_),
    .A(_25487_));
 sky130_as_sc_hs__nand3_2 _32000_ (.A(_24474_),
    .B(_25029_),
    .C(_25487_),
    .Y(_25489_));
 sky130_as_sc_hs__and2_2 _32005_ (.A(_25492_),
    .B(_25493_),
    .Y(_25494_));
 sky130_as_sc_hs__or2_2 _32008_ (.A(_25424_),
    .B(_25495_),
    .Y(_25497_));
 sky130_as_sc_hs__and2_2 _32009_ (.A(_25496_),
    .B(_25497_),
    .Y(_25498_));
 sky130_as_sc_hs__or2_2 _32011_ (.A(_25423_),
    .B(_25498_),
    .Y(_25500_));
 sky130_as_sc_hs__and2_2 _32012_ (.A(_25499_),
    .B(_25500_),
    .Y(_25501_));
 sky130_as_sc_hs__or2_2 _32014_ (.A(_25422_),
    .B(_25501_),
    .Y(_25503_));
 sky130_as_sc_hs__and2_2 _32015_ (.A(_25502_),
    .B(_25503_),
    .Y(_25504_));
 sky130_as_sc_hs__or2_2 _32017_ (.A(_25409_),
    .B(_25504_),
    .Y(_25506_));
 sky130_as_sc_hs__and2_2 _32018_ (.A(_25505_),
    .B(_25506_),
    .Y(_25507_));
 sky130_as_sc_hs__or2_2 _32020_ (.A(_25408_),
    .B(_25507_),
    .Y(_25509_));
 sky130_as_sc_hs__and2_2 _32021_ (.A(_25508_),
    .B(_25509_),
    .Y(_25510_));
 sky130_as_sc_hs__or2_2 _32023_ (.A(_25407_),
    .B(_25510_),
    .Y(_25512_));
 sky130_as_sc_hs__and2_2 _32024_ (.A(_25511_),
    .B(_25512_),
    .Y(_25513_));
 sky130_as_sc_hs__or2_2 _32026_ (.A(_25360_),
    .B(_25513_),
    .Y(_25515_));
 sky130_as_sc_hs__and2_2 _32027_ (.A(_25514_),
    .B(_25515_),
    .Y(_25516_));
 sky130_as_sc_hs__and2_2 _32031_ (.A(_24729_),
    .B(net439),
    .Y(_25520_));
 sky130_as_sc_hs__and2_2 _32032_ (.A(net480),
    .B(net444),
    .Y(_25521_));
 sky130_as_sc_hs__and2_2 _32033_ (.A(net90),
    .B(net435),
    .Y(_25522_));
 sky130_as_sc_hs__or2_2 _32035_ (.A(_25521_),
    .B(_25522_),
    .Y(_25524_));
 sky130_as_sc_hs__and2_2 _32036_ (.A(_25523_),
    .B(_25524_),
    .Y(_25525_));
 sky130_as_sc_hs__or2_2 _32038_ (.A(_25520_),
    .B(_25525_),
    .Y(_25527_));
 sky130_as_sc_hs__or2_2 _32040_ (.A(_25096_),
    .B(_25528_),
    .Y(_25529_));
 sky130_as_sc_hs__and2_2 _32042_ (.A(_25529_),
    .B(_25530_),
    .Y(_25531_));
 sky130_as_sc_hs__or2_2 _32044_ (.A(_25519_),
    .B(_25531_),
    .Y(_25533_));
 sky130_as_sc_hs__and2_2 _32045_ (.A(_25532_),
    .B(_25533_),
    .Y(_25534_));
 sky130_as_sc_hs__or2_2 _32048_ (.A(_25534_),
    .B(_25535_),
    .Y(_25537_));
 sky130_as_sc_hs__and2_2 _32049_ (.A(_25536_),
    .B(_25537_),
    .Y(_25538_));
 sky130_as_sc_hs__and2_2 _32050_ (.A(_24808_),
    .B(net430),
    .Y(_25539_));
 sky130_as_sc_hs__and2_2 _32051_ (.A(_24814_),
    .B(net432),
    .Y(_25540_));
 sky130_as_sc_hs__nand3_2 _32052_ (.A(_24216_),
    .B(_24818_),
    .C(_24819_),
    .Y(_25541_));
 sky130_as_sc_hs__nand3_2 _32053_ (.A(_24216_),
    .B(net437),
    .C(_25540_),
    .Y(_25542_));
 sky130_as_sc_hs__nand2b_2 _32054_ (.B(_25541_),
    .Y(_25543_),
    .A(_25540_));
 sky130_as_sc_hs__and2_2 _32055_ (.A(_25542_),
    .B(_25543_),
    .Y(_25544_));
 sky130_as_sc_hs__nand3_2 _32056_ (.A(_25539_),
    .B(_25542_),
    .C(_25543_),
    .Y(_25545_));
 sky130_as_sc_hs__or2_2 _32057_ (.A(_25539_),
    .B(_25544_),
    .Y(_25546_));
 sky130_as_sc_hs__and2_2 _32058_ (.A(_25545_),
    .B(_25546_),
    .Y(_25547_));
 sky130_as_sc_hs__and2_2 _32059_ (.A(_24768_),
    .B(net84),
    .Y(_25548_));
 sky130_as_sc_hs__and2_2 _32060_ (.A(net479),
    .B(_24774_),
    .Y(_25549_));
 sky130_as_sc_hs__and2_2 _32061_ (.A(_23712_),
    .B(net441),
    .Y(_25550_));
 sky130_as_sc_hs__or2_2 _32063_ (.A(_25549_),
    .B(_25550_),
    .Y(_25552_));
 sky130_as_sc_hs__and2_2 _32064_ (.A(_25551_),
    .B(_25552_),
    .Y(_25553_));
 sky130_as_sc_hs__or2_2 _32066_ (.A(_25548_),
    .B(_25553_),
    .Y(_25555_));
 sky130_as_sc_hs__and2_2 _32067_ (.A(_25554_),
    .B(_25555_),
    .Y(_25556_));
 sky130_as_sc_hs__or2_2 _32070_ (.A(_25556_),
    .B(_25557_),
    .Y(_25559_));
 sky130_as_sc_hs__and2_2 _32071_ (.A(_25558_),
    .B(_25559_),
    .Y(_25560_));
 sky130_as_sc_hs__or2_2 _32073_ (.A(_25547_),
    .B(_25560_),
    .Y(_25562_));
 sky130_as_sc_hs__and2_2 _32074_ (.A(_25561_),
    .B(_25562_),
    .Y(_25563_));
 sky130_as_sc_hs__or2_2 _32076_ (.A(_25538_),
    .B(_25563_),
    .Y(_25565_));
 sky130_as_sc_hs__and2_2 _32077_ (.A(_25564_),
    .B(_25565_),
    .Y(_25566_));
 sky130_as_sc_hs__or2_2 _32079_ (.A(_25518_),
    .B(_25566_),
    .Y(_25568_));
 sky130_as_sc_hs__and2_2 _32080_ (.A(_25567_),
    .B(_25568_),
    .Y(_25569_));
 sky130_as_sc_hs__or2_2 _32082_ (.A(_25517_),
    .B(_25569_),
    .Y(_25571_));
 sky130_as_sc_hs__and2_2 _32083_ (.A(_25570_),
    .B(_25571_),
    .Y(_25572_));
 sky130_as_sc_hs__or2_2 _32085_ (.A(_25516_),
    .B(_25572_),
    .Y(_25574_));
 sky130_as_sc_hs__and2_2 _32086_ (.A(_25573_),
    .B(_25574_),
    .Y(_25575_));
 sky130_as_sc_hs__or2_2 _32088_ (.A(_25359_),
    .B(_25575_),
    .Y(_25577_));
 sky130_as_sc_hs__and2_2 _32089_ (.A(_25576_),
    .B(_25577_),
    .Y(_25578_));
 sky130_as_sc_hs__and2_2 _32096_ (.A(net121),
    .B(_25205_),
    .Y(_25585_));
 sky130_as_sc_hs__and2_2 _32097_ (.A(_25211_),
    .B(net428),
    .Y(_25586_));
 sky130_as_sc_hs__or2_2 _32099_ (.A(_25585_),
    .B(_25586_),
    .Y(_25588_));
 sky130_as_sc_hs__and2_2 _32100_ (.A(_25587_),
    .B(_25588_),
    .Y(_25589_));
 sky130_as_sc_hs__or2_2 _32102_ (.A(_25584_),
    .B(_25589_),
    .Y(_25591_));
 sky130_as_sc_hs__or2_2 _32104_ (.A(_25320_),
    .B(_25592_),
    .Y(_25593_));
 sky130_as_sc_hs__and2_2 _32106_ (.A(_25593_),
    .B(_25594_),
    .Y(_25595_));
 sky130_as_sc_hs__or2_2 _32108_ (.A(_25583_),
    .B(_25595_),
    .Y(_25597_));
 sky130_as_sc_hs__and2_2 _32109_ (.A(_25596_),
    .B(_25597_),
    .Y(_25598_));
 sky130_as_sc_hs__or2_2 _32111_ (.A(_25582_),
    .B(_25598_),
    .Y(_25600_));
 sky130_as_sc_hs__and2_2 _32112_ (.A(_25599_),
    .B(_25600_),
    .Y(_25601_));
 sky130_as_sc_hs__or2_2 _32114_ (.A(_25581_),
    .B(_25601_),
    .Y(_25603_));
 sky130_as_sc_hs__and2_2 _32115_ (.A(_25602_),
    .B(_25603_),
    .Y(_25604_));
 sky130_as_sc_hs__or2_2 _32116_ (.A(_23703_),
    .B(_23705_),
    .Y(_25605_));
 sky130_as_sc_hs__and2_2 _32117_ (.A(_23706_),
    .B(_25605_),
    .Y(_25606_));
 sky130_as_sc_hs__or2_2 _32119_ (.A(_25604_),
    .B(_25606_),
    .Y(_25608_));
 sky130_as_sc_hs__and2_2 _32120_ (.A(_25607_),
    .B(_25608_),
    .Y(_25609_));
 sky130_as_sc_hs__or2_2 _32122_ (.A(_25580_),
    .B(_25609_),
    .Y(_25611_));
 sky130_as_sc_hs__and2_2 _32123_ (.A(_25610_),
    .B(_25611_),
    .Y(_25612_));
 sky130_as_sc_hs__or2_2 _32125_ (.A(_25579_),
    .B(_25612_),
    .Y(_25614_));
 sky130_as_sc_hs__and2_2 _32126_ (.A(_25613_),
    .B(_25614_),
    .Y(_25615_));
 sky130_as_sc_hs__or2_2 _32128_ (.A(_25578_),
    .B(_25615_),
    .Y(_25617_));
 sky130_as_sc_hs__and2_2 _32129_ (.A(_25616_),
    .B(_25617_),
    .Y(_25618_));
 sky130_as_sc_hs__or2_2 _32132_ (.A(_25358_),
    .B(_25618_),
    .Y(_25621_));
 sky130_as_sc_hs__and2_2 _32133_ (.A(_25619_),
    .B(_25621_),
    .Y(_25622_));
 sky130_as_sc_hs__and2_2 _32142_ (.A(net90),
    .B(net433),
    .Y(_25631_));
 sky130_as_sc_hs__and2_2 _32143_ (.A(_23712_),
    .B(net456),
    .Y(_25632_));
 sky130_as_sc_hs__or2_2 _32145_ (.A(_25631_),
    .B(_25632_),
    .Y(_25634_));
 sky130_as_sc_hs__or2_2 _32147_ (.A(_25364_),
    .B(_25635_),
    .Y(_25636_));
 sky130_as_sc_hs__and2_2 _32149_ (.A(_25636_),
    .B(_25637_),
    .Y(_25638_));
 sky130_as_sc_hs__and2_2 _32150_ (.A(net470),
    .B(_24545_),
    .Y(_25639_));
 sky130_as_sc_hs__nand3_2 _32151_ (.A(_24196_),
    .B(_24197_),
    .C(_24256_),
    .Y(_25640_));
 sky130_as_sc_hs__or2_2 _32153_ (.A(_25640_),
    .B(_25641_),
    .Y(_25642_));
 sky130_as_sc_hs__and2_2 _32155_ (.A(_25642_),
    .B(_25643_),
    .Y(_25644_));
 sky130_as_sc_hs__or2_2 _32157_ (.A(_25639_),
    .B(_25644_),
    .Y(_25646_));
 sky130_as_sc_hs__and2_2 _32158_ (.A(_25645_),
    .B(_25646_),
    .Y(_25647_));
 sky130_as_sc_hs__or2_2 _32160_ (.A(_25638_),
    .B(_25647_),
    .Y(_25649_));
 sky130_as_sc_hs__and2_2 _32161_ (.A(_25648_),
    .B(_25649_),
    .Y(_25650_));
 sky130_as_sc_hs__or2_2 _32163_ (.A(_25630_),
    .B(_25650_),
    .Y(_25652_));
 sky130_as_sc_hs__and2_2 _32164_ (.A(_25651_),
    .B(_25652_),
    .Y(_25653_));
 sky130_as_sc_hs__and2_2 _32167_ (.A(net461),
    .B(net453),
    .Y(_25656_));
 sky130_as_sc_hs__and2_2 _32168_ (.A(net464),
    .B(net455),
    .Y(_25657_));
 sky130_as_sc_hs__and2_2 _32169_ (.A(net462),
    .B(net86),
    .Y(_25658_));
 sky130_as_sc_hs__or2_2 _32170_ (.A(_25657_),
    .B(_25658_),
    .Y(_25659_));
 sky130_as_sc_hs__and2_2 _32172_ (.A(_25659_),
    .B(_25660_),
    .Y(_25661_));
 sky130_as_sc_hs__or2_2 _32174_ (.A(_25656_),
    .B(_25661_),
    .Y(_25663_));
 sky130_as_sc_hs__and2_2 _32175_ (.A(_25662_),
    .B(_25663_),
    .Y(_25664_));
 sky130_as_sc_hs__or2_2 _32177_ (.A(_25655_),
    .B(_25664_),
    .Y(_25666_));
 sky130_as_sc_hs__and2_2 _32178_ (.A(_25665_),
    .B(_25666_),
    .Y(_25667_));
 sky130_as_sc_hs__or2_2 _32180_ (.A(_25654_),
    .B(_25667_),
    .Y(_25669_));
 sky130_as_sc_hs__and2_2 _32181_ (.A(_25668_),
    .B(_25669_),
    .Y(_25670_));
 sky130_as_sc_hs__or2_2 _32183_ (.A(_25653_),
    .B(_25670_),
    .Y(_25672_));
 sky130_as_sc_hs__and2_2 _32184_ (.A(_25671_),
    .B(_25672_),
    .Y(_25673_));
 sky130_as_sc_hs__or2_2 _32186_ (.A(_25629_),
    .B(_25673_),
    .Y(_25675_));
 sky130_as_sc_hs__and2_2 _32187_ (.A(_25674_),
    .B(_25675_),
    .Y(_25676_));
 sky130_as_sc_hs__and2_2 _32190_ (.A(net88),
    .B(net443),
    .Y(_25679_));
 sky130_as_sc_hs__nand3_2 _32192_ (.A(_24535_),
    .B(_24536_),
    .C(net79),
    .Y(_25681_));
 sky130_as_sc_hs__or2_2 _32194_ (.A(_25680_),
    .B(_25681_),
    .Y(_25683_));
 sky130_as_sc_hs__and2_2 _32195_ (.A(_25682_),
    .B(_25683_),
    .Y(_25684_));
 sky130_as_sc_hs__or2_2 _32197_ (.A(_25679_),
    .B(_25684_),
    .Y(_25686_));
 sky130_as_sc_hs__and2_2 _32198_ (.A(_25685_),
    .B(_25686_),
    .Y(_25687_));
 sky130_as_sc_hs__or2_2 _32201_ (.A(_25687_),
    .B(_25688_),
    .Y(_25690_));
 sky130_as_sc_hs__and2_2 _32202_ (.A(_25689_),
    .B(_25690_),
    .Y(_25691_));
 sky130_as_sc_hs__and2_2 _32203_ (.A(net481),
    .B(net450),
    .Y(_25692_));
 sky130_as_sc_hs__and2_2 _32204_ (.A(_23674_),
    .B(net448),
    .Y(_25693_));
 sky130_as_sc_hs__and2_2 _32205_ (.A(net458),
    .B(net426),
    .Y(_25694_));
 sky130_as_sc_hs__or2_2 _32206_ (.A(_25693_),
    .B(_25694_),
    .Y(_25695_));
 sky130_as_sc_hs__and2_2 _32208_ (.A(_25695_),
    .B(_25696_),
    .Y(_25697_));
 sky130_as_sc_hs__or2_2 _32210_ (.A(_25692_),
    .B(_25697_),
    .Y(_25699_));
 sky130_as_sc_hs__and2_2 _32211_ (.A(_25698_),
    .B(_25699_),
    .Y(_25700_));
 sky130_as_sc_hs__or2_2 _32213_ (.A(_25691_),
    .B(_25700_),
    .Y(_25702_));
 sky130_as_sc_hs__and2_2 _32214_ (.A(_25701_),
    .B(_25702_),
    .Y(_25703_));
 sky130_as_sc_hs__or2_2 _32216_ (.A(_25678_),
    .B(_25703_),
    .Y(_25705_));
 sky130_as_sc_hs__and2_2 _32217_ (.A(_25704_),
    .B(_25705_),
    .Y(_25706_));
 sky130_as_sc_hs__or2_2 _32219_ (.A(_25677_),
    .B(_25706_),
    .Y(_25708_));
 sky130_as_sc_hs__and2_2 _32220_ (.A(_25707_),
    .B(_25708_),
    .Y(_25709_));
 sky130_as_sc_hs__or2_2 _32222_ (.A(_25676_),
    .B(_25709_),
    .Y(_25711_));
 sky130_as_sc_hs__and2_2 _32223_ (.A(_25710_),
    .B(_25711_),
    .Y(_25712_));
 sky130_as_sc_hs__or2_2 _32225_ (.A(_25628_),
    .B(_25712_),
    .Y(_25714_));
 sky130_as_sc_hs__and2_2 _32226_ (.A(_25713_),
    .B(_25714_),
    .Y(_25715_));
 sky130_as_sc_hs__and2_2 _32231_ (.A(net473),
    .B(_24729_),
    .Y(_25720_));
 sky130_as_sc_hs__and2_2 _32232_ (.A(net477),
    .B(net445),
    .Y(_25721_));
 sky130_as_sc_hs__and2_2 _32233_ (.A(_24053_),
    .B(net435),
    .Y(_25722_));
 sky130_as_sc_hs__or2_2 _32235_ (.A(_25721_),
    .B(_25722_),
    .Y(_25724_));
 sky130_as_sc_hs__and2_2 _32236_ (.A(_25723_),
    .B(_25724_),
    .Y(_25725_));
 sky130_as_sc_hs__or2_2 _32238_ (.A(_25720_),
    .B(_25725_),
    .Y(_25727_));
 sky130_as_sc_hs__and2_2 _32239_ (.A(_25726_),
    .B(_25727_),
    .Y(_25728_));
 sky130_as_sc_hs__or2_2 _32241_ (.A(_25719_),
    .B(_25728_),
    .Y(_25730_));
 sky130_as_sc_hs__and2_2 _32242_ (.A(_25729_),
    .B(_25730_),
    .Y(_25731_));
 sky130_as_sc_hs__or2_2 _32244_ (.A(_25718_),
    .B(_25731_),
    .Y(_25733_));
 sky130_as_sc_hs__and2_2 _32245_ (.A(_25732_),
    .B(_25733_),
    .Y(_25734_));
 sky130_as_sc_hs__or2_2 _32248_ (.A(_25734_),
    .B(_25735_),
    .Y(_25737_));
 sky130_as_sc_hs__and2_2 _32249_ (.A(_25736_),
    .B(_25737_),
    .Y(_25738_));
 sky130_as_sc_hs__and2_2 _32250_ (.A(_24808_),
    .B(net428),
    .Y(_25739_));
 sky130_as_sc_hs__nand3_2 _32252_ (.A(_24229_),
    .B(_24818_),
    .C(_24819_),
    .Y(_25741_));
 sky130_as_sc_hs__or2_2 _32254_ (.A(_25740_),
    .B(_25741_),
    .Y(_25743_));
 sky130_as_sc_hs__and2_2 _32255_ (.A(_25742_),
    .B(_25743_),
    .Y(_25744_));
 sky130_as_sc_hs__or2_2 _32257_ (.A(_25739_),
    .B(_25744_),
    .Y(_25746_));
 sky130_as_sc_hs__and2_2 _32258_ (.A(_25745_),
    .B(_25746_),
    .Y(_25747_));
 sky130_as_sc_hs__and2_2 _32259_ (.A(_24768_),
    .B(net432),
    .Y(_25748_));
 sky130_as_sc_hs__and2_2 _32260_ (.A(net475),
    .B(_24774_),
    .Y(_25749_));
 sky130_as_sc_hs__and2_2 _32261_ (.A(_24216_),
    .B(net441),
    .Y(_25750_));
 sky130_as_sc_hs__or2_2 _32263_ (.A(_25749_),
    .B(_25750_),
    .Y(_25752_));
 sky130_as_sc_hs__and2_2 _32264_ (.A(_25751_),
    .B(_25752_),
    .Y(_25753_));
 sky130_as_sc_hs__or2_2 _32266_ (.A(_25748_),
    .B(_25753_),
    .Y(_25755_));
 sky130_as_sc_hs__and2_2 _32267_ (.A(_25754_),
    .B(_25755_),
    .Y(_25756_));
 sky130_as_sc_hs__or2_2 _32270_ (.A(_25756_),
    .B(_25757_),
    .Y(_25759_));
 sky130_as_sc_hs__and2_2 _32271_ (.A(_25758_),
    .B(_25759_),
    .Y(_25760_));
 sky130_as_sc_hs__or2_2 _32273_ (.A(_25747_),
    .B(_25760_),
    .Y(_25762_));
 sky130_as_sc_hs__and2_2 _32274_ (.A(_25761_),
    .B(_25762_),
    .Y(_25763_));
 sky130_as_sc_hs__or2_2 _32276_ (.A(_25738_),
    .B(_25763_),
    .Y(_25765_));
 sky130_as_sc_hs__and2_2 _32277_ (.A(_25764_),
    .B(_25765_),
    .Y(_25766_));
 sky130_as_sc_hs__or2_2 _32279_ (.A(_25717_),
    .B(_25766_),
    .Y(_25768_));
 sky130_as_sc_hs__and2_2 _32280_ (.A(_25767_),
    .B(_25768_),
    .Y(_25769_));
 sky130_as_sc_hs__or2_2 _32282_ (.A(_25716_),
    .B(_25769_),
    .Y(_25771_));
 sky130_as_sc_hs__and2_2 _32283_ (.A(_25770_),
    .B(_25771_),
    .Y(_25772_));
 sky130_as_sc_hs__or2_2 _32285_ (.A(_25715_),
    .B(_25772_),
    .Y(_25774_));
 sky130_as_sc_hs__and2_2 _32286_ (.A(_25773_),
    .B(_25774_),
    .Y(_25775_));
 sky130_as_sc_hs__or2_2 _32288_ (.A(_25627_),
    .B(_25775_),
    .Y(_25777_));
 sky130_as_sc_hs__and2_2 _32289_ (.A(_25776_),
    .B(_25777_),
    .Y(_25778_));
 sky130_as_sc_hs__and2_2 _32295_ (.A(net121),
    .B(_25211_),
    .Y(_25784_));
 sky130_as_sc_hs__and2_2 _32296_ (.A(net123),
    .B(_25205_),
    .Y(_25785_));
 sky130_as_sc_hs__or2_2 _32298_ (.A(_25784_),
    .B(_25785_),
    .Y(_25787_));
 sky130_as_sc_hs__and2_2 _32299_ (.A(_25786_),
    .B(_25787_),
    .Y(_25788_));
 sky130_as_sc_hs__or2_2 _32301_ (.A(_25783_),
    .B(_25788_),
    .Y(_25790_));
 sky130_as_sc_hs__or2_2 _32303_ (.A(_25587_),
    .B(_25791_),
    .Y(_25792_));
 sky130_as_sc_hs__and2_2 _32305_ (.A(_25792_),
    .B(_25793_),
    .Y(_25794_));
 sky130_as_sc_hs__or2_2 _32307_ (.A(_25782_),
    .B(_25794_),
    .Y(_25796_));
 sky130_as_sc_hs__and2_2 _32308_ (.A(_25795_),
    .B(_25796_),
    .Y(_25797_));
 sky130_as_sc_hs__or2_2 _32310_ (.A(_25781_),
    .B(_25797_),
    .Y(_25799_));
 sky130_as_sc_hs__and2_2 _32311_ (.A(_25798_),
    .B(_25799_),
    .Y(_25800_));
 sky130_as_sc_hs__or2_2 _32314_ (.A(_25800_),
    .B(_25801_),
    .Y(_25803_));
 sky130_as_sc_hs__and2_2 _32315_ (.A(_25802_),
    .B(_25803_),
    .Y(_25804_));
 sky130_as_sc_hs__and2_2 _32316_ (.A(net479),
    .B(_23702_),
    .Y(_25805_));
 sky130_as_sc_hs__nand3_2 _32319_ (.A(net212),
    .B(_25806_),
    .C(_25807_),
    .Y(_25808_));
 sky130_as_sc_hs__nand3_2 _32322_ (.A(net352),
    .B(_25809_),
    .C(_25810_),
    .Y(_25811_));
 sky130_as_sc_hs__nand3_2 _32323_ (.A(net231),
    .B(_25808_),
    .C(_25811_),
    .Y(_25812_));
 sky130_as_sc_hs__nand3_2 _32326_ (.A(net212),
    .B(_25813_),
    .C(_25814_),
    .Y(_25815_));
 sky130_as_sc_hs__nand3_2 _32329_ (.A(net352),
    .B(_25816_),
    .C(_25817_),
    .Y(_25818_));
 sky130_as_sc_hs__nand3_2 _32330_ (.A(net342),
    .B(_25815_),
    .C(_25818_),
    .Y(_25819_));
 sky130_as_sc_hs__nand3_2 _32333_ (.A(net213),
    .B(_25820_),
    .C(_25821_),
    .Y(_25822_));
 sky130_as_sc_hs__nand3_2 _32336_ (.A(net359),
    .B(_25823_),
    .C(_25824_),
    .Y(_25825_));
 sky130_as_sc_hs__nand3_2 _32337_ (.A(net231),
    .B(_25822_),
    .C(_25825_),
    .Y(_25826_));
 sky130_as_sc_hs__nand3_2 _32340_ (.A(net359),
    .B(_25827_),
    .C(_25828_),
    .Y(_25829_));
 sky130_as_sc_hs__nand3_2 _32343_ (.A(net213),
    .B(_25830_),
    .C(_25831_),
    .Y(_25832_));
 sky130_as_sc_hs__nand3_2 _32344_ (.A(net342),
    .B(_25829_),
    .C(_25832_),
    .Y(_25833_));
 sky130_as_sc_hs__nand3_2 _32345_ (.A(net240),
    .B(_25826_),
    .C(_25833_),
    .Y(_25834_));
 sky130_as_sc_hs__nand3_2 _32346_ (.A(net337),
    .B(_25812_),
    .C(_25819_),
    .Y(_25835_));
 sky130_as_sc_hs__nand3_2 _32347_ (.A(net336),
    .B(_25834_),
    .C(_25835_),
    .Y(_25836_));
 sky130_as_sc_hs__nand3_2 _32350_ (.A(net211),
    .B(_25837_),
    .C(_25838_),
    .Y(_25839_));
 sky130_as_sc_hs__nand3_2 _32353_ (.A(net351),
    .B(_25840_),
    .C(_25841_),
    .Y(_25842_));
 sky130_as_sc_hs__nand3_2 _32354_ (.A(net232),
    .B(_25839_),
    .C(_25842_),
    .Y(_25843_));
 sky130_as_sc_hs__nand3_2 _32357_ (.A(net213),
    .B(_25844_),
    .C(_25845_),
    .Y(_25846_));
 sky130_as_sc_hs__nand3_2 _32360_ (.A(net359),
    .B(_25847_),
    .C(_25848_),
    .Y(_25849_));
 sky130_as_sc_hs__nand3_2 _32361_ (.A(net343),
    .B(_25846_),
    .C(_25849_),
    .Y(_25850_));
 sky130_as_sc_hs__nand3_2 _32364_ (.A(net212),
    .B(_25851_),
    .C(_25852_),
    .Y(_25853_));
 sky130_as_sc_hs__nand3_2 _32367_ (.A(net351),
    .B(_25854_),
    .C(_25855_),
    .Y(_25856_));
 sky130_as_sc_hs__nand3_2 _32368_ (.A(net232),
    .B(_25853_),
    .C(_25856_),
    .Y(_25857_));
 sky130_as_sc_hs__nand3_2 _32371_ (.A(net351),
    .B(_25858_),
    .C(_25859_),
    .Y(_25860_));
 sky130_as_sc_hs__nand3_2 _32374_ (.A(net212),
    .B(_25861_),
    .C(_25862_),
    .Y(_25863_));
 sky130_as_sc_hs__nand3_2 _32375_ (.A(net343),
    .B(_25860_),
    .C(_25863_),
    .Y(_25864_));
 sky130_as_sc_hs__nand3_2 _32376_ (.A(net240),
    .B(_25857_),
    .C(_25864_),
    .Y(_25865_));
 sky130_as_sc_hs__nand3_2 _32377_ (.A(net337),
    .B(_25843_),
    .C(_25850_),
    .Y(_25866_));
 sky130_as_sc_hs__nand3_2 _32378_ (.A(net246),
    .B(_25865_),
    .C(_25866_),
    .Y(_25867_));
 sky130_as_sc_hs__and2_2 _32379_ (.A(_25836_),
    .B(_25867_),
    .Y(_25868_));
 sky130_as_sc_hs__or2_2 _32381_ (.A(_23529_),
    .B(_25868_),
    .Y(_25870_));
 sky130_as_sc_hs__and2_2 _32385_ (.A(_25872_),
    .B(_25873_),
    .Y(_25874_));
 sky130_as_sc_hs__and2_2 _32386_ (.A(net115),
    .B(net424),
    .Y(_25875_));
 sky130_as_sc_hs__and2_2 _32387_ (.A(net482),
    .B(net438),
    .Y(_25876_));
 sky130_as_sc_hs__and2_2 _32388_ (.A(_23636_),
    .B(net84),
    .Y(_25877_));
 sky130_as_sc_hs__or2_2 _32389_ (.A(net197),
    .B(\tholin_riscv.regs[25][29] ),
    .Y(_25878_));
 sky130_as_sc_hs__or2_2 _32390_ (.A(net328),
    .B(\tholin_riscv.regs[24][29] ),
    .Y(_25879_));
 sky130_as_sc_hs__nand3_2 _32391_ (.A(net184),
    .B(_25878_),
    .C(_25879_),
    .Y(_25880_));
 sky130_as_sc_hs__or2_2 _32392_ (.A(net197),
    .B(\tholin_riscv.regs[27][29] ),
    .Y(_25881_));
 sky130_as_sc_hs__or2_2 _32393_ (.A(net328),
    .B(\tholin_riscv.regs[26][29] ),
    .Y(_25882_));
 sky130_as_sc_hs__nand3_2 _32394_ (.A(net279),
    .B(_25881_),
    .C(_25882_),
    .Y(_25883_));
 sky130_as_sc_hs__nand3_2 _32395_ (.A(net165),
    .B(_25880_),
    .C(_25883_),
    .Y(_25884_));
 sky130_as_sc_hs__or2_2 _32396_ (.A(net197),
    .B(\tholin_riscv.regs[29][29] ),
    .Y(_25885_));
 sky130_as_sc_hs__or2_2 _32397_ (.A(net328),
    .B(\tholin_riscv.regs[28][29] ),
    .Y(_25886_));
 sky130_as_sc_hs__nand3_2 _32398_ (.A(net184),
    .B(_25885_),
    .C(_25886_),
    .Y(_25887_));
 sky130_as_sc_hs__or2_2 _32399_ (.A(net197),
    .B(\tholin_riscv.regs[31][29] ),
    .Y(_25888_));
 sky130_as_sc_hs__or2_2 _32400_ (.A(net328),
    .B(\tholin_riscv.regs[30][29] ),
    .Y(_25889_));
 sky130_as_sc_hs__nand3_2 _32401_ (.A(net279),
    .B(_25888_),
    .C(_25889_),
    .Y(_25890_));
 sky130_as_sc_hs__nand3_2 _32402_ (.A(net261),
    .B(_25887_),
    .C(_25890_),
    .Y(_25891_));
 sky130_as_sc_hs__or2_2 _32403_ (.A(net198),
    .B(\tholin_riscv.regs[17][29] ),
    .Y(_25892_));
 sky130_as_sc_hs__or2_2 _32404_ (.A(net329),
    .B(\tholin_riscv.regs[16][29] ),
    .Y(_25893_));
 sky130_as_sc_hs__nand3_2 _32405_ (.A(net184),
    .B(_25892_),
    .C(_25893_),
    .Y(_25894_));
 sky130_as_sc_hs__or2_2 _32406_ (.A(net198),
    .B(\tholin_riscv.regs[19][29] ),
    .Y(_25895_));
 sky130_as_sc_hs__or2_2 _32407_ (.A(net328),
    .B(\tholin_riscv.regs[18][29] ),
    .Y(_25896_));
 sky130_as_sc_hs__nand3_2 _32408_ (.A(net279),
    .B(_25895_),
    .C(_25896_),
    .Y(_25897_));
 sky130_as_sc_hs__nand3_2 _32409_ (.A(net165),
    .B(_25894_),
    .C(_25897_),
    .Y(_25898_));
 sky130_as_sc_hs__or2_2 _32410_ (.A(net197),
    .B(\tholin_riscv.regs[23][29] ),
    .Y(_25899_));
 sky130_as_sc_hs__or2_2 _32411_ (.A(net328),
    .B(\tholin_riscv.regs[22][29] ),
    .Y(_25900_));
 sky130_as_sc_hs__nand3_2 _32412_ (.A(net278),
    .B(_25899_),
    .C(_25900_),
    .Y(_25901_));
 sky130_as_sc_hs__or2_2 _32413_ (.A(net198),
    .B(\tholin_riscv.regs[21][29] ),
    .Y(_25902_));
 sky130_as_sc_hs__or2_2 _32414_ (.A(net328),
    .B(\tholin_riscv.regs[20][29] ),
    .Y(_25903_));
 sky130_as_sc_hs__nand3_2 _32415_ (.A(net184),
    .B(_25902_),
    .C(_25903_),
    .Y(_25904_));
 sky130_as_sc_hs__nand3_2 _32416_ (.A(net261),
    .B(_25901_),
    .C(_25904_),
    .Y(_25905_));
 sky130_as_sc_hs__nand3_2 _32417_ (.A(net155),
    .B(_25898_),
    .C(_25905_),
    .Y(_25906_));
 sky130_as_sc_hs__nand3_2 _32418_ (.A(net252),
    .B(_25884_),
    .C(_25891_),
    .Y(_25907_));
 sky130_as_sc_hs__nand3_2 _32419_ (.A(net248),
    .B(_25906_),
    .C(_25907_),
    .Y(_25908_));
 sky130_as_sc_hs__or2_2 _32420_ (.A(net193),
    .B(\tholin_riscv.regs[9][29] ),
    .Y(_25909_));
 sky130_as_sc_hs__or2_2 _32421_ (.A(net319),
    .B(\tholin_riscv.regs[8][29] ),
    .Y(_25910_));
 sky130_as_sc_hs__nand3_2 _32422_ (.A(net177),
    .B(_25909_),
    .C(_25910_),
    .Y(_25911_));
 sky130_as_sc_hs__or2_2 _32423_ (.A(net194),
    .B(\tholin_riscv.regs[11][29] ),
    .Y(_25912_));
 sky130_as_sc_hs__or2_2 _32424_ (.A(net319),
    .B(\tholin_riscv.regs[10][29] ),
    .Y(_25913_));
 sky130_as_sc_hs__nand3_2 _32425_ (.A(net274),
    .B(_25912_),
    .C(_25913_),
    .Y(_25914_));
 sky130_as_sc_hs__nand3_2 _32426_ (.A(net159),
    .B(_25911_),
    .C(_25914_),
    .Y(_25915_));
 sky130_as_sc_hs__or2_2 _32427_ (.A(net194),
    .B(\tholin_riscv.regs[13][29] ),
    .Y(_25916_));
 sky130_as_sc_hs__or2_2 _32428_ (.A(net319),
    .B(\tholin_riscv.regs[12][29] ),
    .Y(_25917_));
 sky130_as_sc_hs__nand3_2 _32429_ (.A(net177),
    .B(_25916_),
    .C(_25917_),
    .Y(_25918_));
 sky130_as_sc_hs__or2_2 _32430_ (.A(net194),
    .B(\tholin_riscv.regs[15][29] ),
    .Y(_25919_));
 sky130_as_sc_hs__or2_2 _32431_ (.A(net319),
    .B(\tholin_riscv.regs[14][29] ),
    .Y(_25920_));
 sky130_as_sc_hs__nand3_2 _32432_ (.A(net273),
    .B(_25919_),
    .C(_25920_),
    .Y(_25921_));
 sky130_as_sc_hs__nand3_2 _32433_ (.A(net259),
    .B(_25918_),
    .C(_25921_),
    .Y(_25922_));
 sky130_as_sc_hs__or2_2 _32434_ (.A(net194),
    .B(\tholin_riscv.regs[1][29] ),
    .Y(_25923_));
 sky130_as_sc_hs__or2_2 _32435_ (.A(net319),
    .B(\tholin_riscv.regs[0][29] ),
    .Y(_25924_));
 sky130_as_sc_hs__nand3_2 _32436_ (.A(net177),
    .B(_25923_),
    .C(_25924_),
    .Y(_25925_));
 sky130_as_sc_hs__or2_2 _32437_ (.A(net194),
    .B(\tholin_riscv.regs[3][29] ),
    .Y(_25926_));
 sky130_as_sc_hs__or2_2 _32438_ (.A(net319),
    .B(\tholin_riscv.regs[2][29] ),
    .Y(_25927_));
 sky130_as_sc_hs__nand3_2 _32439_ (.A(net273),
    .B(_25926_),
    .C(_25927_),
    .Y(_25928_));
 sky130_as_sc_hs__nand3_2 _32440_ (.A(net159),
    .B(_25925_),
    .C(_25928_),
    .Y(_25929_));
 sky130_as_sc_hs__or2_2 _32441_ (.A(net193),
    .B(\tholin_riscv.regs[7][29] ),
    .Y(_25930_));
 sky130_as_sc_hs__or2_2 _32442_ (.A(net319),
    .B(\tholin_riscv.regs[6][29] ),
    .Y(_25931_));
 sky130_as_sc_hs__nand3_2 _32443_ (.A(net273),
    .B(_25930_),
    .C(_25931_),
    .Y(_25932_));
 sky130_as_sc_hs__or2_2 _32444_ (.A(net194),
    .B(\tholin_riscv.regs[5][29] ),
    .Y(_25933_));
 sky130_as_sc_hs__or2_2 _32445_ (.A(net319),
    .B(\tholin_riscv.regs[4][29] ),
    .Y(_25934_));
 sky130_as_sc_hs__nand3_2 _32446_ (.A(net177),
    .B(_25933_),
    .C(_25934_),
    .Y(_25935_));
 sky130_as_sc_hs__nand3_2 _32447_ (.A(net259),
    .B(_25932_),
    .C(_25935_),
    .Y(_25936_));
 sky130_as_sc_hs__nand3_2 _32448_ (.A(net152),
    .B(_25929_),
    .C(_25936_),
    .Y(_25937_));
 sky130_as_sc_hs__nand3_2 _32449_ (.A(net249),
    .B(_25915_),
    .C(_25922_),
    .Y(_01721_));
 sky130_as_sc_hs__nand3_2 _32450_ (.A(net150),
    .B(_25937_),
    .C(_01721_),
    .Y(_01722_));
 sky130_as_sc_hs__inv_2 _32452_ (.Y(_01724_),
    .A(_01723_));
 sky130_as_sc_hs__or2_2 _32453_ (.A(_25489_),
    .B(_01724_),
    .Y(_01725_));
 sky130_as_sc_hs__and2_2 _32458_ (.A(_01728_),
    .B(_01729_),
    .Y(_01730_));
 sky130_as_sc_hs__and2_2 _32459_ (.A(net112),
    .B(net422),
    .Y(_01731_));
 sky130_as_sc_hs__or2_2 _32461_ (.A(_25877_),
    .B(_01731_),
    .Y(_01733_));
 sky130_as_sc_hs__and2_2 _32462_ (.A(_01732_),
    .B(_01733_),
    .Y(_01734_));
 sky130_as_sc_hs__or2_2 _32464_ (.A(_25876_),
    .B(_01734_),
    .Y(_01736_));
 sky130_as_sc_hs__or2_2 _32466_ (.A(_23659_),
    .B(_01737_),
    .Y(_01738_));
 sky130_as_sc_hs__and2_2 _32468_ (.A(_01738_),
    .B(_01739_),
    .Y(_01740_));
 sky130_as_sc_hs__or2_2 _32470_ (.A(_25875_),
    .B(_01740_),
    .Y(_01742_));
 sky130_as_sc_hs__and2_2 _32471_ (.A(_01741_),
    .B(_01742_),
    .Y(_01743_));
 sky130_as_sc_hs__or2_2 _32474_ (.A(_01743_),
    .B(_01744_),
    .Y(_01746_));
 sky130_as_sc_hs__and2_2 _32475_ (.A(_01745_),
    .B(_01746_),
    .Y(_01747_));
 sky130_as_sc_hs__or2_2 _32477_ (.A(_25805_),
    .B(_01747_),
    .Y(_01749_));
 sky130_as_sc_hs__and2_2 _32478_ (.A(_01748_),
    .B(_01749_),
    .Y(_01750_));
 sky130_as_sc_hs__or2_2 _32480_ (.A(_25804_),
    .B(_01750_),
    .Y(_01752_));
 sky130_as_sc_hs__and2_2 _32481_ (.A(_01751_),
    .B(_01752_),
    .Y(_01753_));
 sky130_as_sc_hs__or2_2 _32483_ (.A(_25780_),
    .B(_01753_),
    .Y(_01755_));
 sky130_as_sc_hs__and2_2 _32484_ (.A(_01754_),
    .B(_01755_),
    .Y(_01756_));
 sky130_as_sc_hs__or2_2 _32486_ (.A(_25779_),
    .B(_01756_),
    .Y(_01758_));
 sky130_as_sc_hs__and2_2 _32487_ (.A(_01757_),
    .B(_01758_),
    .Y(_01759_));
 sky130_as_sc_hs__or2_2 _32489_ (.A(_25778_),
    .B(_01759_),
    .Y(_01761_));
 sky130_as_sc_hs__and2_2 _32490_ (.A(_01760_),
    .B(_01761_),
    .Y(_01762_));
 sky130_as_sc_hs__or2_2 _32492_ (.A(_25626_),
    .B(_01762_),
    .Y(_01764_));
 sky130_as_sc_hs__and2_2 _32493_ (.A(_01763_),
    .B(_01764_),
    .Y(_01765_));
 sky130_as_sc_hs__or2_2 _32495_ (.A(_25625_),
    .B(_01765_),
    .Y(_01767_));
 sky130_as_sc_hs__and2_2 _32496_ (.A(_01766_),
    .B(_01767_),
    .Y(_01768_));
 sky130_as_sc_hs__or2_2 _32498_ (.A(_25624_),
    .B(_01768_),
    .Y(_01770_));
 sky130_as_sc_hs__and2_2 _32499_ (.A(_01769_),
    .B(_01770_),
    .Y(_01771_));
 sky130_as_sc_hs__or2_2 _32501_ (.A(_23707_),
    .B(_01771_),
    .Y(_01773_));
 sky130_as_sc_hs__or2_2 _32503_ (.A(_24248_),
    .B(_24250_),
    .Y(_01775_));
 sky130_as_sc_hs__and2_2 _32504_ (.A(_24251_),
    .B(_01775_),
    .Y(_01776_));
 sky130_as_sc_hs__and2_2 _32505_ (.A(_24053_),
    .B(net464),
    .Y(_01777_));
 sky130_as_sc_hs__and2_2 _32506_ (.A(_23712_),
    .B(net462),
    .Y(_01778_));
 sky130_as_sc_hs__and2_2 _32508_ (.A(_24216_),
    .B(net461),
    .Y(_01780_));
 sky130_as_sc_hs__or2_2 _32509_ (.A(_01777_),
    .B(_01778_),
    .Y(_01781_));
 sky130_as_sc_hs__and2_2 _32510_ (.A(_01779_),
    .B(_01781_),
    .Y(_01782_));
 sky130_as_sc_hs__and2_2 _32513_ (.A(net468),
    .B(net458),
    .Y(_01785_));
 sky130_as_sc_hs__nand3_2 _32514_ (.A(net113),
    .B(_24196_),
    .C(_24197_),
    .Y(_01786_));
 sky130_as_sc_hs__nand3_2 _32515_ (.A(net113),
    .B(net467),
    .C(_01785_),
    .Y(_01787_));
 sky130_as_sc_hs__and2_2 _32516_ (.A(_24047_),
    .B(net90),
    .Y(_01788_));
 sky130_as_sc_hs__nand2b_2 _32517_ (.B(_01786_),
    .Y(_01789_),
    .A(_01785_));
 sky130_as_sc_hs__and2_2 _32518_ (.A(_01787_),
    .B(_01789_),
    .Y(_01790_));
 sky130_as_sc_hs__or2_2 _32521_ (.A(_24235_),
    .B(_24237_),
    .Y(_01793_));
 sky130_as_sc_hs__and2_2 _32522_ (.A(_24238_),
    .B(_01793_),
    .Y(_01794_));
 sky130_as_sc_hs__or2_2 _32524_ (.A(_01792_),
    .B(_01794_),
    .Y(_01796_));
 sky130_as_sc_hs__and2_2 _32525_ (.A(_01795_),
    .B(_01796_),
    .Y(_01797_));
 sky130_as_sc_hs__or2_2 _32527_ (.A(_01784_),
    .B(_01797_),
    .Y(_01799_));
 sky130_as_sc_hs__and2_2 _32528_ (.A(_01798_),
    .B(_01799_),
    .Y(_01800_));
 sky130_as_sc_hs__or2_2 _32530_ (.A(_24205_),
    .B(_24271_),
    .Y(_01802_));
 sky130_as_sc_hs__or2_2 _32532_ (.A(_01801_),
    .B(_01803_),
    .Y(_01804_));
 sky130_as_sc_hs__and2_2 _32534_ (.A(_01804_),
    .B(_01805_),
    .Y(_01806_));
 sky130_as_sc_hs__and2_2 _32535_ (.A(_24229_),
    .B(_24527_),
    .Y(_01807_));
 sky130_as_sc_hs__nand3_2 _32536_ (.A(_24256_),
    .B(_24535_),
    .C(_24536_),
    .Y(_01808_));
 sky130_as_sc_hs__nand3_2 _32537_ (.A(_24256_),
    .B(net89),
    .C(_01807_),
    .Y(_01809_));
 sky130_as_sc_hs__and2_2 _32538_ (.A(_24501_),
    .B(net87),
    .Y(_01810_));
 sky130_as_sc_hs__nand2b_2 _32539_ (.B(_01808_),
    .Y(_01811_),
    .A(_01807_));
 sky130_as_sc_hs__and2_2 _32540_ (.A(_01809_),
    .B(_01811_),
    .Y(_01812_));
 sky130_as_sc_hs__or2_2 _32543_ (.A(_24551_),
    .B(_24553_),
    .Y(_01815_));
 sky130_as_sc_hs__and2_2 _32544_ (.A(_24554_),
    .B(_01815_),
    .Y(_01816_));
 sky130_as_sc_hs__or2_2 _32546_ (.A(_01814_),
    .B(_01816_),
    .Y(_01818_));
 sky130_as_sc_hs__and2_2 _32547_ (.A(_01817_),
    .B(_01818_),
    .Y(_01819_));
 sky130_as_sc_hs__or2_2 _32548_ (.A(_24748_),
    .B(_24749_),
    .Y(_01820_));
 sky130_as_sc_hs__and2_2 _32549_ (.A(_24750_),
    .B(_01820_),
    .Y(_01821_));
 sky130_as_sc_hs__or2_2 _32553_ (.A(_24573_),
    .B(_24600_),
    .Y(_01825_));
 sky130_as_sc_hs__and2_2 _32554_ (.A(_24601_),
    .B(_01825_),
    .Y(_01826_));
 sky130_as_sc_hs__or2_2 _32556_ (.A(_01824_),
    .B(_01826_),
    .Y(_01828_));
 sky130_as_sc_hs__and2_2 _32557_ (.A(_01827_),
    .B(_01828_),
    .Y(_01829_));
 sky130_as_sc_hs__or2_2 _32559_ (.A(_01823_),
    .B(_01829_),
    .Y(_01831_));
 sky130_as_sc_hs__and2_2 _32560_ (.A(_01830_),
    .B(_01831_),
    .Y(_01832_));
 sky130_as_sc_hs__or2_2 _32563_ (.A(_24522_),
    .B(_24636_),
    .Y(_01835_));
 sky130_as_sc_hs__and2_2 _32564_ (.A(_24637_),
    .B(_01835_),
    .Y(_01836_));
 sky130_as_sc_hs__or2_2 _32566_ (.A(_01834_),
    .B(_01836_),
    .Y(_01838_));
 sky130_as_sc_hs__and2_2 _32567_ (.A(_01837_),
    .B(_01838_),
    .Y(_01839_));
 sky130_as_sc_hs__and2_2 _32569_ (.A(_24759_),
    .B(_01840_),
    .Y(_01841_));
 sky130_as_sc_hs__and2_2 _32570_ (.A(_24545_),
    .B(net448),
    .Y(_01842_));
 sky130_as_sc_hs__and2_2 _32571_ (.A(net455),
    .B(net451),
    .Y(_01843_));
 sky130_as_sc_hs__or2_2 _32573_ (.A(_24754_),
    .B(_24755_),
    .Y(_01845_));
 sky130_as_sc_hs__or2_2 _32575_ (.A(_01844_),
    .B(_01846_),
    .Y(_01847_));
 sky130_as_sc_hs__and2_2 _32576_ (.A(net85),
    .B(net444),
    .Y(_01848_));
 sky130_as_sc_hs__and2_2 _32577_ (.A(net446),
    .B(_24729_),
    .Y(_01849_));
 sky130_as_sc_hs__or2_2 _32581_ (.A(_01850_),
    .B(_01852_),
    .Y(_01853_));
 sky130_as_sc_hs__or2_2 _32584_ (.A(_01841_),
    .B(_01854_),
    .Y(_01856_));
 sky130_as_sc_hs__and2_2 _32585_ (.A(_01855_),
    .B(_01856_),
    .Y(_01857_));
 sky130_as_sc_hs__or2_2 _32586_ (.A(_25188_),
    .B(_25197_),
    .Y(_01858_));
 sky130_as_sc_hs__and2_2 _32587_ (.A(_25198_),
    .B(_01858_),
    .Y(_01859_));
 sky130_as_sc_hs__or2_2 _32591_ (.A(_24763_),
    .B(_24830_),
    .Y(_01863_));
 sky130_as_sc_hs__and2_2 _32592_ (.A(_24831_),
    .B(_01863_),
    .Y(_01864_));
 sky130_as_sc_hs__or2_2 _32594_ (.A(_01862_),
    .B(_01864_),
    .Y(_01866_));
 sky130_as_sc_hs__and2_2 _32595_ (.A(_01865_),
    .B(_01866_),
    .Y(_01867_));
 sky130_as_sc_hs__or2_2 _32597_ (.A(_01861_),
    .B(_01867_),
    .Y(_01869_));
 sky130_as_sc_hs__and2_2 _32598_ (.A(_01868_),
    .B(_01869_),
    .Y(_01870_));
 sky130_as_sc_hs__or2_2 _32601_ (.A(_24718_),
    .B(_24960_),
    .Y(_01873_));
 sky130_as_sc_hs__and2_2 _32602_ (.A(_24961_),
    .B(_01873_),
    .Y(_01874_));
 sky130_as_sc_hs__or2_2 _32604_ (.A(_01872_),
    .B(_01874_),
    .Y(_01876_));
 sky130_as_sc_hs__and2_2 _32605_ (.A(_01875_),
    .B(_01876_),
    .Y(_01877_));
 sky130_as_sc_hs__and2_2 _32606_ (.A(net443),
    .B(_24774_),
    .Y(_01878_));
 sky130_as_sc_hs__and2_2 _32607_ (.A(net481),
    .B(_24768_),
    .Y(_01879_));
 sky130_as_sc_hs__or2_2 _32609_ (.A(_25181_),
    .B(_25182_),
    .Y(_01881_));
 sky130_as_sc_hs__or2_2 _32611_ (.A(_01880_),
    .B(_01882_),
    .Y(_01883_));
 sky130_as_sc_hs__and2_2 _32613_ (.A(_01883_),
    .B(_01884_),
    .Y(_01885_));
 sky130_as_sc_hs__or2_2 _32614_ (.A(_25229_),
    .B(_25231_),
    .Y(_01886_));
 sky130_as_sc_hs__and2_2 _32615_ (.A(_25232_),
    .B(_01886_),
    .Y(_01887_));
 sky130_as_sc_hs__and2_2 _32619_ (.A(_25242_),
    .B(_01890_),
    .Y(_01891_));
 sky130_as_sc_hs__and2_2 _32621_ (.A(net477),
    .B(_24814_),
    .Y(_01893_));
 sky130_as_sc_hs__and2_2 _32622_ (.A(net439),
    .B(_24808_),
    .Y(_01894_));
 sky130_as_sc_hs__or2_2 _32624_ (.A(_25237_),
    .B(_25238_),
    .Y(_01896_));
 sky130_as_sc_hs__or2_2 _32626_ (.A(_01895_),
    .B(_01897_),
    .Y(_01898_));
 sky130_as_sc_hs__and2_2 _32627_ (.A(net473),
    .B(_25211_),
    .Y(_01899_));
 sky130_as_sc_hs__and2_2 _32628_ (.A(net479),
    .B(_25205_),
    .Y(_01900_));
 sky130_as_sc_hs__or2_2 _32632_ (.A(_01901_),
    .B(_01903_),
    .Y(_01904_));
 sky130_as_sc_hs__or2_2 _32634_ (.A(_01889_),
    .B(_01891_),
    .Y(_01906_));
 sky130_as_sc_hs__and2_2 _32635_ (.A(_01892_),
    .B(_01906_),
    .Y(_01907_));
 sky130_as_sc_hs__or2_2 _32638_ (.A(_25243_),
    .B(_25245_),
    .Y(_01910_));
 sky130_as_sc_hs__and2_2 _32639_ (.A(_25246_),
    .B(_01910_),
    .Y(_01911_));
 sky130_as_sc_hs__or2_2 _32641_ (.A(_01909_),
    .B(_01911_),
    .Y(_01913_));
 sky130_as_sc_hs__and2_2 _32642_ (.A(_01912_),
    .B(_01913_),
    .Y(_01914_));
 sky130_as_sc_hs__and2_2 _32643_ (.A(net481),
    .B(_23702_),
    .Y(_01915_));
 sky130_as_sc_hs__or2_2 _32644_ (.A(_25300_),
    .B(_25302_),
    .Y(_01916_));
 sky130_as_sc_hs__and2_2 _32645_ (.A(_25303_),
    .B(_01916_),
    .Y(_01917_));
 sky130_as_sc_hs__and2_2 _32646_ (.A(net480),
    .B(_23636_),
    .Y(_01918_));
 sky130_as_sc_hs__and2_2 _32647_ (.A(net482),
    .B(net446),
    .Y(_01919_));
 sky130_as_sc_hs__or2_2 _32649_ (.A(_25296_),
    .B(_25297_),
    .Y(_01921_));
 sky130_as_sc_hs__or2_2 _32651_ (.A(_01920_),
    .B(_01922_),
    .Y(_01923_));
 sky130_as_sc_hs__and2_2 _32652_ (.A(net115),
    .B(net432),
    .Y(_01924_));
 sky130_as_sc_hs__and2_2 _32654_ (.A(_01923_),
    .B(_01925_),
    .Y(_01926_));
 sky130_as_sc_hs__or2_2 _32658_ (.A(_01917_),
    .B(_01928_),
    .Y(_01930_));
 sky130_as_sc_hs__and2_2 _32659_ (.A(_01929_),
    .B(_01930_),
    .Y(_01931_));
 sky130_as_sc_hs__or2_2 _32661_ (.A(_01915_),
    .B(_01931_),
    .Y(_01933_));
 sky130_as_sc_hs__and2_2 _32662_ (.A(_01932_),
    .B(_01933_),
    .Y(_01934_));
 sky130_as_sc_hs__or2_2 _32666_ (.A(_25275_),
    .B(_25310_),
    .Y(_01938_));
 sky130_as_sc_hs__and2_2 _32667_ (.A(_25311_),
    .B(_01938_),
    .Y(_01939_));
 sky130_as_sc_hs__or2_2 _32669_ (.A(_01937_),
    .B(_01939_),
    .Y(_01941_));
 sky130_as_sc_hs__and2_2 _32670_ (.A(_01940_),
    .B(_01941_),
    .Y(_01942_));
 sky130_as_sc_hs__or2_2 _32672_ (.A(_01936_),
    .B(_01942_),
    .Y(_01944_));
 sky130_as_sc_hs__and2_2 _32673_ (.A(_01943_),
    .B(_01944_),
    .Y(_01945_));
 sky130_as_sc_hs__or2_2 _32676_ (.A(_25180_),
    .B(_25356_),
    .Y(_01948_));
 sky130_as_sc_hs__and2_2 _32677_ (.A(_25357_),
    .B(_01948_),
    .Y(_01949_));
 sky130_as_sc_hs__or2_2 _32680_ (.A(_01947_),
    .B(_01949_),
    .Y(_01952_));
 sky130_as_sc_hs__and2_2 _32681_ (.A(_01950_),
    .B(_01952_),
    .Y(_01953_));
 sky130_as_sc_hs__or2_2 _32684_ (.A(_25620_),
    .B(_25622_),
    .Y(_01956_));
 sky130_as_sc_hs__and2_2 _32685_ (.A(_25623_),
    .B(_01956_),
    .Y(_01957_));
 sky130_as_sc_hs__or2_2 _32688_ (.A(_01955_),
    .B(_01957_),
    .Y(_01960_));
 sky130_as_sc_hs__and2_2 _32689_ (.A(_01958_),
    .B(_01960_),
    .Y(_01961_));
 sky130_as_sc_hs__and2_2 _32691_ (.A(_01958_),
    .B(_01962_),
    .Y(_01963_));
 sky130_as_sc_hs__or2_2 _32693_ (.A(_01774_),
    .B(_01963_),
    .Y(_01965_));
 sky130_as_sc_hs__and2_2 _32694_ (.A(_01964_),
    .B(_01965_),
    .Y(_01966_));
 sky130_as_sc_hs__or2_2 _32695_ (.A(_01959_),
    .B(_01961_),
    .Y(_01967_));
 sky130_as_sc_hs__and2_2 _32696_ (.A(_01962_),
    .B(_01967_),
    .Y(_01968_));
 sky130_as_sc_hs__or2_2 _32697_ (.A(_01788_),
    .B(_01790_),
    .Y(_01969_));
 sky130_as_sc_hs__and2_2 _32698_ (.A(_01791_),
    .B(_01969_),
    .Y(_01970_));
 sky130_as_sc_hs__and2_2 _32699_ (.A(net90),
    .B(net464),
    .Y(_01971_));
 sky130_as_sc_hs__and2_2 _32700_ (.A(_24053_),
    .B(net463),
    .Y(_01972_));
 sky130_as_sc_hs__and2_2 _32702_ (.A(_23712_),
    .B(net461),
    .Y(_01974_));
 sky130_as_sc_hs__or2_2 _32703_ (.A(_01971_),
    .B(_01972_),
    .Y(_01975_));
 sky130_as_sc_hs__and2_2 _32704_ (.A(_01973_),
    .B(_01975_),
    .Y(_01976_));
 sky130_as_sc_hs__and2_2 _32707_ (.A(net112),
    .B(net469),
    .Y(_01979_));
 sky130_as_sc_hs__and2_2 _32708_ (.A(net470),
    .B(net458),
    .Y(_01980_));
 sky130_as_sc_hs__or2_2 _32710_ (.A(_01780_),
    .B(_01782_),
    .Y(_01982_));
 sky130_as_sc_hs__or2_2 _32712_ (.A(_01981_),
    .B(_01983_),
    .Y(_01984_));
 sky130_as_sc_hs__and2_2 _32714_ (.A(_01984_),
    .B(_01985_),
    .Y(_01986_));
 sky130_as_sc_hs__or2_2 _32716_ (.A(_01978_),
    .B(_01986_),
    .Y(_01988_));
 sky130_as_sc_hs__and2_2 _32717_ (.A(_01987_),
    .B(_01988_),
    .Y(_01989_));
 sky130_as_sc_hs__or2_2 _32719_ (.A(_01776_),
    .B(_01800_),
    .Y(_01991_));
 sky130_as_sc_hs__or2_2 _32721_ (.A(_01990_),
    .B(_01992_),
    .Y(_01993_));
 sky130_as_sc_hs__and2_2 _32723_ (.A(_01993_),
    .B(_01994_),
    .Y(_01995_));
 sky130_as_sc_hs__and2_2 _32724_ (.A(_24216_),
    .B(_24527_),
    .Y(_01996_));
 sky130_as_sc_hs__nand3_2 _32725_ (.A(_24229_),
    .B(_24535_),
    .C(_24536_),
    .Y(_01997_));
 sky130_as_sc_hs__nand3_2 _32726_ (.A(_24229_),
    .B(net89),
    .C(_01996_),
    .Y(_01998_));
 sky130_as_sc_hs__and2_2 _32727_ (.A(_24256_),
    .B(net87),
    .Y(_01999_));
 sky130_as_sc_hs__nand2b_2 _32728_ (.B(_01997_),
    .Y(_02000_),
    .A(_01996_));
 sky130_as_sc_hs__and2_2 _32729_ (.A(_01998_),
    .B(_02000_),
    .Y(_02001_));
 sky130_as_sc_hs__or2_2 _32732_ (.A(_01810_),
    .B(_01812_),
    .Y(_02004_));
 sky130_as_sc_hs__and2_2 _32733_ (.A(_01813_),
    .B(_02004_),
    .Y(_02005_));
 sky130_as_sc_hs__or2_2 _32735_ (.A(_02003_),
    .B(_02005_),
    .Y(_02007_));
 sky130_as_sc_hs__and2_2 _32736_ (.A(_02006_),
    .B(_02007_),
    .Y(_02008_));
 sky130_as_sc_hs__or2_2 _32737_ (.A(_01842_),
    .B(_01843_),
    .Y(_02009_));
 sky130_as_sc_hs__and2_2 _32738_ (.A(_01844_),
    .B(_02009_),
    .Y(_02010_));
 sky130_as_sc_hs__or2_2 _32742_ (.A(_01819_),
    .B(_01821_),
    .Y(_02014_));
 sky130_as_sc_hs__and2_2 _32743_ (.A(_01822_),
    .B(_02014_),
    .Y(_02015_));
 sky130_as_sc_hs__or2_2 _32745_ (.A(_02013_),
    .B(_02015_),
    .Y(_02017_));
 sky130_as_sc_hs__and2_2 _32746_ (.A(_02016_),
    .B(_02017_),
    .Y(_02018_));
 sky130_as_sc_hs__or2_2 _32748_ (.A(_02012_),
    .B(_02018_),
    .Y(_02020_));
 sky130_as_sc_hs__and2_2 _32749_ (.A(_02019_),
    .B(_02020_),
    .Y(_02021_));
 sky130_as_sc_hs__or2_2 _32752_ (.A(_01806_),
    .B(_01832_),
    .Y(_02024_));
 sky130_as_sc_hs__and2_2 _32753_ (.A(_01833_),
    .B(_02024_),
    .Y(_02025_));
 sky130_as_sc_hs__or2_2 _32755_ (.A(_02023_),
    .B(_02025_),
    .Y(_02027_));
 sky130_as_sc_hs__and2_2 _32756_ (.A(_02026_),
    .B(_02027_),
    .Y(_02028_));
 sky130_as_sc_hs__and2_2 _32758_ (.A(_01853_),
    .B(_02029_),
    .Y(_02030_));
 sky130_as_sc_hs__and2_2 _32759_ (.A(_24501_),
    .B(net448),
    .Y(_02031_));
 sky130_as_sc_hs__and2_2 _32760_ (.A(_24545_),
    .B(net450),
    .Y(_02032_));
 sky130_as_sc_hs__or2_2 _32762_ (.A(_01848_),
    .B(_01849_),
    .Y(_02034_));
 sky130_as_sc_hs__or2_2 _32764_ (.A(_02033_),
    .B(_02035_),
    .Y(_02036_));
 sky130_as_sc_hs__and2_2 _32765_ (.A(net454),
    .B(net444),
    .Y(_02037_));
 sky130_as_sc_hs__and2_2 _32766_ (.A(net452),
    .B(_24729_),
    .Y(_02038_));
 sky130_as_sc_hs__or2_2 _32770_ (.A(_02039_),
    .B(_02041_),
    .Y(_02042_));
 sky130_as_sc_hs__or2_2 _32773_ (.A(_02030_),
    .B(_02043_),
    .Y(_02045_));
 sky130_as_sc_hs__and2_2 _32774_ (.A(_02044_),
    .B(_02045_),
    .Y(_02046_));
 sky130_as_sc_hs__or2_2 _32775_ (.A(_01885_),
    .B(_01887_),
    .Y(_02047_));
 sky130_as_sc_hs__and2_2 _32776_ (.A(_01888_),
    .B(_02047_),
    .Y(_02048_));
 sky130_as_sc_hs__or2_2 _32780_ (.A(_01857_),
    .B(_01859_),
    .Y(_02052_));
 sky130_as_sc_hs__and2_2 _32781_ (.A(_01860_),
    .B(_02052_),
    .Y(_02053_));
 sky130_as_sc_hs__or2_2 _32783_ (.A(_02051_),
    .B(_02053_),
    .Y(_02055_));
 sky130_as_sc_hs__and2_2 _32784_ (.A(_02054_),
    .B(_02055_),
    .Y(_02056_));
 sky130_as_sc_hs__or2_2 _32786_ (.A(_02050_),
    .B(_02056_),
    .Y(_02058_));
 sky130_as_sc_hs__and2_2 _32787_ (.A(_02057_),
    .B(_02058_),
    .Y(_02059_));
 sky130_as_sc_hs__or2_2 _32790_ (.A(_01839_),
    .B(_01870_),
    .Y(_02062_));
 sky130_as_sc_hs__and2_2 _32791_ (.A(_01871_),
    .B(_02062_),
    .Y(_02063_));
 sky130_as_sc_hs__or2_2 _32793_ (.A(_02061_),
    .B(_02063_),
    .Y(_02065_));
 sky130_as_sc_hs__and2_2 _32794_ (.A(_02064_),
    .B(_02065_),
    .Y(_02066_));
 sky130_as_sc_hs__and2_2 _32795_ (.A(net78),
    .B(_24774_),
    .Y(_02067_));
 sky130_as_sc_hs__and2_2 _32796_ (.A(_23674_),
    .B(_24768_),
    .Y(_02068_));
 sky130_as_sc_hs__or2_2 _32798_ (.A(_01878_),
    .B(_01879_),
    .Y(_02070_));
 sky130_as_sc_hs__or2_2 _32800_ (.A(_02069_),
    .B(_02071_),
    .Y(_02072_));
 sky130_as_sc_hs__or2_2 _32801_ (.A(_01893_),
    .B(_01894_),
    .Y(_02073_));
 sky130_as_sc_hs__and2_2 _32802_ (.A(_01895_),
    .B(_02073_),
    .Y(_02074_));
 sky130_as_sc_hs__and2_2 _32804_ (.A(_02072_),
    .B(_02075_),
    .Y(_02076_));
 sky130_as_sc_hs__and2_2 _32808_ (.A(_01904_),
    .B(_02079_),
    .Y(_02080_));
 sky130_as_sc_hs__and2_2 _32810_ (.A(net481),
    .B(_24814_),
    .Y(_02082_));
 sky130_as_sc_hs__and2_2 _32811_ (.A(net477),
    .B(_24808_),
    .Y(_02083_));
 sky130_as_sc_hs__or2_2 _32813_ (.A(_01899_),
    .B(_01900_),
    .Y(_02085_));
 sky130_as_sc_hs__or2_2 _32815_ (.A(_02084_),
    .B(_02086_),
    .Y(_02087_));
 sky130_as_sc_hs__and2_2 _32816_ (.A(net439),
    .B(_25211_),
    .Y(_02088_));
 sky130_as_sc_hs__and2_2 _32817_ (.A(net473),
    .B(_25205_),
    .Y(_02089_));
 sky130_as_sc_hs__or2_2 _32821_ (.A(_02090_),
    .B(_02092_),
    .Y(_02093_));
 sky130_as_sc_hs__or2_2 _32823_ (.A(_02078_),
    .B(_02080_),
    .Y(_02095_));
 sky130_as_sc_hs__and2_2 _32824_ (.A(_02081_),
    .B(_02095_),
    .Y(_02096_));
 sky130_as_sc_hs__or2_2 _32827_ (.A(_01905_),
    .B(_01907_),
    .Y(_02099_));
 sky130_as_sc_hs__and2_2 _32828_ (.A(_01908_),
    .B(_02099_),
    .Y(_02100_));
 sky130_as_sc_hs__or2_2 _32830_ (.A(_02098_),
    .B(_02100_),
    .Y(_02102_));
 sky130_as_sc_hs__and2_2 _32831_ (.A(_02101_),
    .B(_02102_),
    .Y(_02103_));
 sky130_as_sc_hs__and2_2 _32832_ (.A(_23674_),
    .B(_23702_),
    .Y(_02104_));
 sky130_as_sc_hs__or2_2 _32833_ (.A(_01924_),
    .B(_01926_),
    .Y(_02105_));
 sky130_as_sc_hs__and2_2 _32834_ (.A(_01927_),
    .B(_02105_),
    .Y(_02106_));
 sky130_as_sc_hs__and2_2 _32835_ (.A(_23636_),
    .B(_23674_),
    .Y(_02107_));
 sky130_as_sc_hs__and2_2 _32836_ (.A(net482),
    .B(net452),
    .Y(_02108_));
 sky130_as_sc_hs__or2_2 _32838_ (.A(_01918_),
    .B(_01919_),
    .Y(_02110_));
 sky130_as_sc_hs__or2_2 _32840_ (.A(_02109_),
    .B(_02111_),
    .Y(_02112_));
 sky130_as_sc_hs__and2_2 _32841_ (.A(net115),
    .B(net84),
    .Y(_02113_));
 sky130_as_sc_hs__and2_2 _32843_ (.A(_02112_),
    .B(_02114_),
    .Y(_02115_));
 sky130_as_sc_hs__or2_2 _32847_ (.A(_02106_),
    .B(_02117_),
    .Y(_02119_));
 sky130_as_sc_hs__and2_2 _32848_ (.A(_02118_),
    .B(_02119_),
    .Y(_02120_));
 sky130_as_sc_hs__or2_2 _32850_ (.A(_02104_),
    .B(_02120_),
    .Y(_02122_));
 sky130_as_sc_hs__and2_2 _32851_ (.A(_02121_),
    .B(_02122_),
    .Y(_02123_));
 sky130_as_sc_hs__or2_2 _32855_ (.A(_01914_),
    .B(_01934_),
    .Y(_02127_));
 sky130_as_sc_hs__and2_2 _32856_ (.A(_01935_),
    .B(_02127_),
    .Y(_02128_));
 sky130_as_sc_hs__or2_2 _32858_ (.A(_02126_),
    .B(_02128_),
    .Y(_02130_));
 sky130_as_sc_hs__and2_2 _32859_ (.A(_02129_),
    .B(_02130_),
    .Y(_02131_));
 sky130_as_sc_hs__or2_2 _32861_ (.A(_02125_),
    .B(_02131_),
    .Y(_02133_));
 sky130_as_sc_hs__and2_2 _32862_ (.A(_02132_),
    .B(_02133_),
    .Y(_02134_));
 sky130_as_sc_hs__nand3_2 _32863_ (.A(_02066_),
    .B(_02132_),
    .C(_02133_),
    .Y(_02135_));
 sky130_as_sc_hs__or2_2 _32865_ (.A(_01877_),
    .B(_01945_),
    .Y(_02137_));
 sky130_as_sc_hs__and2_2 _32866_ (.A(_01946_),
    .B(_02137_),
    .Y(_02138_));
 sky130_as_sc_hs__or2_2 _32869_ (.A(_02136_),
    .B(_02138_),
    .Y(_02141_));
 sky130_as_sc_hs__and2_2 _32870_ (.A(_02139_),
    .B(_02141_),
    .Y(_02142_));
 sky130_as_sc_hs__or2_2 _32873_ (.A(_01951_),
    .B(_01953_),
    .Y(_02145_));
 sky130_as_sc_hs__and2_2 _32874_ (.A(_01954_),
    .B(_02145_),
    .Y(_02146_));
 sky130_as_sc_hs__or2_2 _32877_ (.A(_02144_),
    .B(_02146_),
    .Y(_02149_));
 sky130_as_sc_hs__and2_2 _32878_ (.A(_02147_),
    .B(_02149_),
    .Y(_02150_));
 sky130_as_sc_hs__or2_2 _32882_ (.A(_01968_),
    .B(_02152_),
    .Y(_02154_));
 sky130_as_sc_hs__and2_2 _32883_ (.A(_02153_),
    .B(_02154_),
    .Y(_02155_));
 sky130_as_sc_hs__and2_2 _32884_ (.A(_01966_),
    .B(_02155_),
    .Y(_02156_));
 sky130_as_sc_hs__and2_2 _32892_ (.A(_24053_),
    .B(_25035_),
    .Y(_02164_));
 sky130_as_sc_hs__and2_2 _32893_ (.A(_24216_),
    .B(net456),
    .Y(_02165_));
 sky130_as_sc_hs__or2_2 _32895_ (.A(_02164_),
    .B(_02165_),
    .Y(_02167_));
 sky130_as_sc_hs__or2_2 _32897_ (.A(_25633_),
    .B(_02168_),
    .Y(_02169_));
 sky130_as_sc_hs__and2_2 _32899_ (.A(_02169_),
    .B(_02170_),
    .Y(_02171_));
 sky130_as_sc_hs__and2_2 _32900_ (.A(net470),
    .B(net454),
    .Y(_02172_));
 sky130_as_sc_hs__and2_2 _32901_ (.A(net467),
    .B(_24501_),
    .Y(_02173_));
 sky130_as_sc_hs__and2_2 _32902_ (.A(net469),
    .B(_24545_),
    .Y(_02174_));
 sky130_as_sc_hs__or2_2 _32904_ (.A(_02173_),
    .B(_02174_),
    .Y(_02176_));
 sky130_as_sc_hs__and2_2 _32905_ (.A(_02175_),
    .B(_02176_),
    .Y(_02177_));
 sky130_as_sc_hs__or2_2 _32907_ (.A(_02172_),
    .B(_02177_),
    .Y(_02179_));
 sky130_as_sc_hs__and2_2 _32908_ (.A(_02178_),
    .B(_02179_),
    .Y(_02180_));
 sky130_as_sc_hs__or2_2 _32910_ (.A(_02171_),
    .B(_02180_),
    .Y(_02182_));
 sky130_as_sc_hs__and2_2 _32911_ (.A(_02181_),
    .B(_02182_),
    .Y(_02183_));
 sky130_as_sc_hs__or2_2 _32913_ (.A(_02163_),
    .B(_02183_),
    .Y(_02185_));
 sky130_as_sc_hs__and2_2 _32914_ (.A(_02184_),
    .B(_02185_),
    .Y(_02186_));
 sky130_as_sc_hs__and2_2 _32917_ (.A(net461),
    .B(net447),
    .Y(_02189_));
 sky130_as_sc_hs__and2_2 _32918_ (.A(net464),
    .B(net85),
    .Y(_02190_));
 sky130_as_sc_hs__and2_2 _32919_ (.A(net462),
    .B(net453),
    .Y(_02191_));
 sky130_as_sc_hs__or2_2 _32920_ (.A(_02190_),
    .B(_02191_),
    .Y(_02192_));
 sky130_as_sc_hs__and2_2 _32922_ (.A(_02192_),
    .B(_02193_),
    .Y(_02194_));
 sky130_as_sc_hs__or2_2 _32924_ (.A(_02189_),
    .B(_02194_),
    .Y(_02196_));
 sky130_as_sc_hs__and2_2 _32925_ (.A(_02195_),
    .B(_02196_),
    .Y(_02197_));
 sky130_as_sc_hs__or2_2 _32927_ (.A(_02188_),
    .B(_02197_),
    .Y(_02199_));
 sky130_as_sc_hs__and2_2 _32928_ (.A(_02198_),
    .B(_02199_),
    .Y(_02200_));
 sky130_as_sc_hs__or2_2 _32930_ (.A(_02187_),
    .B(_02200_),
    .Y(_02202_));
 sky130_as_sc_hs__and2_2 _32931_ (.A(_02201_),
    .B(_02202_),
    .Y(_02203_));
 sky130_as_sc_hs__or2_2 _32933_ (.A(_02186_),
    .B(_02203_),
    .Y(_02205_));
 sky130_as_sc_hs__and2_2 _32934_ (.A(_02204_),
    .B(_02205_),
    .Y(_02206_));
 sky130_as_sc_hs__or2_2 _32936_ (.A(_02162_),
    .B(_02206_),
    .Y(_02208_));
 sky130_as_sc_hs__and2_2 _32937_ (.A(_02207_),
    .B(_02208_),
    .Y(_02209_));
 sky130_as_sc_hs__and2_2 _32940_ (.A(_23674_),
    .B(net87),
    .Y(_02212_));
 sky130_as_sc_hs__and2_2 _32941_ (.A(_24527_),
    .B(net79),
    .Y(_02213_));
 sky130_as_sc_hs__and2_2 _32942_ (.A(net89),
    .B(net443),
    .Y(_02214_));
 sky130_as_sc_hs__or2_2 _32943_ (.A(_02213_),
    .B(_02214_),
    .Y(_02215_));
 sky130_as_sc_hs__and2_2 _32945_ (.A(_02215_),
    .B(_02216_),
    .Y(_02217_));
 sky130_as_sc_hs__or2_2 _32947_ (.A(_02212_),
    .B(_02217_),
    .Y(_02219_));
 sky130_as_sc_hs__and2_2 _32948_ (.A(_02218_),
    .B(_02219_),
    .Y(_02220_));
 sky130_as_sc_hs__or2_2 _32951_ (.A(_02220_),
    .B(_02221_),
    .Y(_02223_));
 sky130_as_sc_hs__and2_2 _32952_ (.A(_02222_),
    .B(_02223_),
    .Y(_02224_));
 sky130_as_sc_hs__and2_2 _32953_ (.A(net477),
    .B(net450),
    .Y(_02225_));
 sky130_as_sc_hs__and2_2 _32954_ (.A(net481),
    .B(net448),
    .Y(_02226_));
 sky130_as_sc_hs__and2_2 _32955_ (.A(net90),
    .B(net426),
    .Y(_02227_));
 sky130_as_sc_hs__or2_2 _32956_ (.A(_02226_),
    .B(_02227_),
    .Y(_02228_));
 sky130_as_sc_hs__and2_2 _32958_ (.A(_02228_),
    .B(_02229_),
    .Y(_02230_));
 sky130_as_sc_hs__or2_2 _32960_ (.A(_02225_),
    .B(_02230_),
    .Y(_02232_));
 sky130_as_sc_hs__and2_2 _32961_ (.A(_02231_),
    .B(_02232_),
    .Y(_02233_));
 sky130_as_sc_hs__or2_2 _32963_ (.A(_02224_),
    .B(_02233_),
    .Y(_02235_));
 sky130_as_sc_hs__and2_2 _32964_ (.A(_02234_),
    .B(_02235_),
    .Y(_02236_));
 sky130_as_sc_hs__or2_2 _32966_ (.A(_02211_),
    .B(_02236_),
    .Y(_02238_));
 sky130_as_sc_hs__and2_2 _32967_ (.A(_02237_),
    .B(_02238_),
    .Y(_02239_));
 sky130_as_sc_hs__or2_2 _32969_ (.A(_02210_),
    .B(_02239_),
    .Y(_02241_));
 sky130_as_sc_hs__and2_2 _32970_ (.A(_02240_),
    .B(_02241_),
    .Y(_02242_));
 sky130_as_sc_hs__or2_2 _32972_ (.A(_02209_),
    .B(_02242_),
    .Y(_02244_));
 sky130_as_sc_hs__and2_2 _32973_ (.A(_02243_),
    .B(_02244_),
    .Y(_02245_));
 sky130_as_sc_hs__or2_2 _32975_ (.A(_02161_),
    .B(_02245_),
    .Y(_02247_));
 sky130_as_sc_hs__and2_2 _32976_ (.A(_02246_),
    .B(_02247_),
    .Y(_02248_));
 sky130_as_sc_hs__and2_2 _32981_ (.A(net479),
    .B(_24729_),
    .Y(_02253_));
 sky130_as_sc_hs__and2_2 _32982_ (.A(net445),
    .B(net439),
    .Y(_02254_));
 sky130_as_sc_hs__and2_2 _32983_ (.A(_23712_),
    .B(net435),
    .Y(_02255_));
 sky130_as_sc_hs__or2_2 _32984_ (.A(_02254_),
    .B(_02255_),
    .Y(_02256_));
 sky130_as_sc_hs__and2_2 _32986_ (.A(_02256_),
    .B(_02257_),
    .Y(_02258_));
 sky130_as_sc_hs__or2_2 _32988_ (.A(_02253_),
    .B(_02258_),
    .Y(_02260_));
 sky130_as_sc_hs__and2_2 _32989_ (.A(_02259_),
    .B(_02260_),
    .Y(_02261_));
 sky130_as_sc_hs__or2_2 _32991_ (.A(_02252_),
    .B(_02261_),
    .Y(_02263_));
 sky130_as_sc_hs__and2_2 _32992_ (.A(_02262_),
    .B(_02263_),
    .Y(_02264_));
 sky130_as_sc_hs__or2_2 _32994_ (.A(_02251_),
    .B(_02264_),
    .Y(_02266_));
 sky130_as_sc_hs__and2_2 _32995_ (.A(_02265_),
    .B(_02266_),
    .Y(_02267_));
 sky130_as_sc_hs__or2_2 _32998_ (.A(_02267_),
    .B(_02268_),
    .Y(_02270_));
 sky130_as_sc_hs__and2_2 _32999_ (.A(_02269_),
    .B(_02270_),
    .Y(_02271_));
 sky130_as_sc_hs__and2_2 _33000_ (.A(_24768_),
    .B(net430),
    .Y(_02272_));
 sky130_as_sc_hs__and2_2 _33001_ (.A(_24774_),
    .B(net84),
    .Y(_02273_));
 sky130_as_sc_hs__and2_2 _33002_ (.A(_24229_),
    .B(net441),
    .Y(_02274_));
 sky130_as_sc_hs__or2_2 _33003_ (.A(_02273_),
    .B(_02274_),
    .Y(_02275_));
 sky130_as_sc_hs__and2_2 _33005_ (.A(_02275_),
    .B(_02276_),
    .Y(_02277_));
 sky130_as_sc_hs__or2_2 _33007_ (.A(_02272_),
    .B(_02277_),
    .Y(_02279_));
 sky130_as_sc_hs__and2_2 _33008_ (.A(_02278_),
    .B(_02279_),
    .Y(_02280_));
 sky130_as_sc_hs__or2_2 _33011_ (.A(_02280_),
    .B(_02281_),
    .Y(_02283_));
 sky130_as_sc_hs__and2_2 _33012_ (.A(_02282_),
    .B(_02283_),
    .Y(_02284_));
 sky130_as_sc_hs__nand3_2 _33014_ (.A(_24256_),
    .B(_24818_),
    .C(_24819_),
    .Y(_02286_));
 sky130_as_sc_hs__or2_2 _33016_ (.A(_02285_),
    .B(_02286_),
    .Y(_02288_));
 sky130_as_sc_hs__and2_2 _33017_ (.A(_02287_),
    .B(_02288_),
    .Y(_02289_));
 sky130_as_sc_hs__and2_2 _33018_ (.A(net121),
    .B(_24808_),
    .Y(_02290_));
 sky130_as_sc_hs__or2_2 _33020_ (.A(_02289_),
    .B(_02290_),
    .Y(_02292_));
 sky130_as_sc_hs__and2_2 _33021_ (.A(_02291_),
    .B(_02292_),
    .Y(_02293_));
 sky130_as_sc_hs__or2_2 _33023_ (.A(_02284_),
    .B(_02293_),
    .Y(_02295_));
 sky130_as_sc_hs__and2_2 _33024_ (.A(_02294_),
    .B(_02295_),
    .Y(_02296_));
 sky130_as_sc_hs__or2_2 _33026_ (.A(_02271_),
    .B(_02296_),
    .Y(_02298_));
 sky130_as_sc_hs__and2_2 _33027_ (.A(_02297_),
    .B(_02298_),
    .Y(_02299_));
 sky130_as_sc_hs__or2_2 _33029_ (.A(_02250_),
    .B(_02299_),
    .Y(_02301_));
 sky130_as_sc_hs__and2_2 _33030_ (.A(_02300_),
    .B(_02301_),
    .Y(_02302_));
 sky130_as_sc_hs__or2_2 _33032_ (.A(_02249_),
    .B(_02302_),
    .Y(_02304_));
 sky130_as_sc_hs__and2_2 _33033_ (.A(_02303_),
    .B(_02304_),
    .Y(_02305_));
 sky130_as_sc_hs__or2_2 _33035_ (.A(_02248_),
    .B(_02305_),
    .Y(_02307_));
 sky130_as_sc_hs__and2_2 _33036_ (.A(_02306_),
    .B(_02307_),
    .Y(_02308_));
 sky130_as_sc_hs__or2_2 _33038_ (.A(_02160_),
    .B(_02308_),
    .Y(_02310_));
 sky130_as_sc_hs__and2_2 _33039_ (.A(_02309_),
    .B(_02310_),
    .Y(_02311_));
 sky130_as_sc_hs__and2_2 _33045_ (.A(_25205_),
    .B(net424),
    .Y(_02317_));
 sky130_as_sc_hs__and2_2 _33046_ (.A(net123),
    .B(_25211_),
    .Y(_02318_));
 sky130_as_sc_hs__nand3_2 _33049_ (.A(net183),
    .B(_02319_),
    .C(_02320_),
    .Y(_02321_));
 sky130_as_sc_hs__nand3_2 _33052_ (.A(net278),
    .B(_02322_),
    .C(_02323_),
    .Y(_02324_));
 sky130_as_sc_hs__nand3_2 _33053_ (.A(net163),
    .B(_02321_),
    .C(_02324_),
    .Y(_02325_));
 sky130_as_sc_hs__nand3_2 _33056_ (.A(net183),
    .B(_02326_),
    .C(_02327_),
    .Y(_02328_));
 sky130_as_sc_hs__nand3_2 _33059_ (.A(net278),
    .B(_02329_),
    .C(_02330_),
    .Y(_02331_));
 sky130_as_sc_hs__nand3_2 _33060_ (.A(net261),
    .B(_02328_),
    .C(_02331_),
    .Y(_02332_));
 sky130_as_sc_hs__nand3_2 _33063_ (.A(net183),
    .B(_02333_),
    .C(_02334_),
    .Y(_02335_));
 sky130_as_sc_hs__nand3_2 _33066_ (.A(net278),
    .B(_02336_),
    .C(_02337_),
    .Y(_02338_));
 sky130_as_sc_hs__nand3_2 _33067_ (.A(net163),
    .B(_02335_),
    .C(_02338_),
    .Y(_02339_));
 sky130_as_sc_hs__nand3_2 _33070_ (.A(net278),
    .B(_02340_),
    .C(_02341_),
    .Y(_02342_));
 sky130_as_sc_hs__nand3_2 _33073_ (.A(net183),
    .B(_02343_),
    .C(_02344_),
    .Y(_02345_));
 sky130_as_sc_hs__nand3_2 _33074_ (.A(net261),
    .B(_02342_),
    .C(_02345_),
    .Y(_02346_));
 sky130_as_sc_hs__nand3_2 _33075_ (.A(net155),
    .B(_02339_),
    .C(_02346_),
    .Y(_02347_));
 sky130_as_sc_hs__nand3_2 _33076_ (.A(net252),
    .B(_02325_),
    .C(_02332_),
    .Y(_02348_));
 sky130_as_sc_hs__nand3_2 _33077_ (.A(net248),
    .B(_02347_),
    .C(_02348_),
    .Y(_02349_));
 sky130_as_sc_hs__nand3_2 _33080_ (.A(net177),
    .B(_02350_),
    .C(_02351_),
    .Y(_02352_));
 sky130_as_sc_hs__nand3_2 _33083_ (.A(net273),
    .B(_02353_),
    .C(_02354_),
    .Y(_02355_));
 sky130_as_sc_hs__nand3_2 _33084_ (.A(net159),
    .B(_02352_),
    .C(_02355_),
    .Y(_02356_));
 sky130_as_sc_hs__nand3_2 _33087_ (.A(net177),
    .B(_02357_),
    .C(_02358_),
    .Y(_02359_));
 sky130_as_sc_hs__nand3_2 _33090_ (.A(net273),
    .B(_02360_),
    .C(_02361_),
    .Y(_02362_));
 sky130_as_sc_hs__nand3_2 _33091_ (.A(net258),
    .B(_02359_),
    .C(_02362_),
    .Y(_02363_));
 sky130_as_sc_hs__nand3_2 _33094_ (.A(net177),
    .B(_02364_),
    .C(_02365_),
    .Y(_02366_));
 sky130_as_sc_hs__nand3_2 _33097_ (.A(net273),
    .B(_02367_),
    .C(_02368_),
    .Y(_02369_));
 sky130_as_sc_hs__nand3_2 _33098_ (.A(net159),
    .B(_02366_),
    .C(_02369_),
    .Y(_02370_));
 sky130_as_sc_hs__nand3_2 _33101_ (.A(net273),
    .B(_02371_),
    .C(_02372_),
    .Y(_02373_));
 sky130_as_sc_hs__nand3_2 _33104_ (.A(net177),
    .B(_02374_),
    .C(_02375_),
    .Y(_02376_));
 sky130_as_sc_hs__nand3_2 _33105_ (.A(net258),
    .B(_02373_),
    .C(_02376_),
    .Y(_02377_));
 sky130_as_sc_hs__nand3_2 _33106_ (.A(net152),
    .B(_02370_),
    .C(_02377_),
    .Y(_02378_));
 sky130_as_sc_hs__nand3_2 _33107_ (.A(net249),
    .B(_02356_),
    .C(_02363_),
    .Y(_02379_));
 sky130_as_sc_hs__nand3_2 _33108_ (.A(_19538_),
    .B(_02378_),
    .C(_02379_),
    .Y(_02380_));
 sky130_as_sc_hs__or2_2 _33110_ (.A(_01725_),
    .B(_02381_),
    .Y(_02382_));
 sky130_as_sc_hs__or2_2 _33114_ (.A(_23607_),
    .B(_02381_),
    .Y(_02386_));
 sky130_as_sc_hs__and2_2 _33115_ (.A(_02385_),
    .B(_02386_),
    .Y(_02387_));
 sky130_as_sc_hs__and2_2 _33116_ (.A(net112),
    .B(net129),
    .Y(_02388_));
 sky130_as_sc_hs__or2_2 _33117_ (.A(_02318_),
    .B(_02388_),
    .Y(_02389_));
 sky130_as_sc_hs__and2_2 _33119_ (.A(_02389_),
    .B(_02390_),
    .Y(_02391_));
 sky130_as_sc_hs__or2_2 _33121_ (.A(_02317_),
    .B(_02391_),
    .Y(_02393_));
 sky130_as_sc_hs__and2_2 _33122_ (.A(_02392_),
    .B(_02393_),
    .Y(_02394_));
 sky130_as_sc_hs__or2_2 _33124_ (.A(_02316_),
    .B(_02394_),
    .Y(_02396_));
 sky130_as_sc_hs__or2_2 _33126_ (.A(_25786_),
    .B(_02397_),
    .Y(_02398_));
 sky130_as_sc_hs__and2_2 _33128_ (.A(_02398_),
    .B(_02399_),
    .Y(_02400_));
 sky130_as_sc_hs__or2_2 _33130_ (.A(_02315_),
    .B(_02400_),
    .Y(_02402_));
 sky130_as_sc_hs__and2_2 _33131_ (.A(_02401_),
    .B(_02402_),
    .Y(_02403_));
 sky130_as_sc_hs__or2_2 _33133_ (.A(_02314_),
    .B(_02403_),
    .Y(_02405_));
 sky130_as_sc_hs__and2_2 _33134_ (.A(_02404_),
    .B(_02405_),
    .Y(_02406_));
 sky130_as_sc_hs__or2_2 _33137_ (.A(_02406_),
    .B(_02407_),
    .Y(_02409_));
 sky130_as_sc_hs__and2_2 _33138_ (.A(_02408_),
    .B(_02409_),
    .Y(_02410_));
 sky130_as_sc_hs__and2_2 _33139_ (.A(net475),
    .B(_23702_),
    .Y(_02411_));
 sky130_as_sc_hs__nand3_2 _33142_ (.A(net212),
    .B(_02412_),
    .C(_02413_),
    .Y(_02414_));
 sky130_as_sc_hs__nand3_2 _33145_ (.A(net352),
    .B(_02415_),
    .C(_02416_),
    .Y(_02417_));
 sky130_as_sc_hs__nand3_2 _33146_ (.A(net231),
    .B(_02414_),
    .C(_02417_),
    .Y(_02418_));
 sky130_as_sc_hs__nand3_2 _33149_ (.A(net212),
    .B(_02419_),
    .C(_02420_),
    .Y(_02421_));
 sky130_as_sc_hs__nand3_2 _33152_ (.A(net352),
    .B(_02422_),
    .C(_02423_),
    .Y(_02424_));
 sky130_as_sc_hs__nand3_2 _33153_ (.A(net342),
    .B(_02421_),
    .C(_02424_),
    .Y(_02425_));
 sky130_as_sc_hs__nand3_2 _33156_ (.A(net211),
    .B(_02426_),
    .C(_02427_),
    .Y(_02428_));
 sky130_as_sc_hs__nand3_2 _33159_ (.A(net351),
    .B(_02429_),
    .C(_02430_),
    .Y(_02431_));
 sky130_as_sc_hs__nand3_2 _33160_ (.A(net232),
    .B(_02428_),
    .C(_02431_),
    .Y(_02432_));
 sky130_as_sc_hs__nand3_2 _33163_ (.A(net351),
    .B(_02433_),
    .C(_02434_),
    .Y(_02435_));
 sky130_as_sc_hs__nand3_2 _33166_ (.A(net212),
    .B(_02436_),
    .C(_02437_),
    .Y(_02438_));
 sky130_as_sc_hs__nand3_2 _33167_ (.A(net343),
    .B(_02435_),
    .C(_02438_),
    .Y(_02439_));
 sky130_as_sc_hs__nand3_2 _33168_ (.A(net240),
    .B(_02432_),
    .C(_02439_),
    .Y(_02440_));
 sky130_as_sc_hs__nand3_2 _33169_ (.A(net337),
    .B(_02418_),
    .C(_02425_),
    .Y(_02441_));
 sky130_as_sc_hs__nand3_2 _33170_ (.A(net336),
    .B(_02440_),
    .C(_02441_),
    .Y(_02442_));
 sky130_as_sc_hs__nand3_2 _33173_ (.A(net211),
    .B(_02443_),
    .C(_02444_),
    .Y(_02445_));
 sky130_as_sc_hs__nand3_2 _33176_ (.A(net351),
    .B(_02446_),
    .C(_02447_),
    .Y(_02448_));
 sky130_as_sc_hs__nand3_2 _33177_ (.A(net232),
    .B(_02445_),
    .C(_02448_),
    .Y(_02449_));
 sky130_as_sc_hs__nand3_2 _33180_ (.A(net211),
    .B(_02450_),
    .C(_02451_),
    .Y(_02452_));
 sky130_as_sc_hs__nand3_2 _33183_ (.A(net351),
    .B(_02453_),
    .C(_02454_),
    .Y(_02455_));
 sky130_as_sc_hs__nand3_2 _33184_ (.A(net343),
    .B(_02452_),
    .C(_02455_),
    .Y(_02456_));
 sky130_as_sc_hs__nand3_2 _33187_ (.A(net212),
    .B(_02457_),
    .C(_02458_),
    .Y(_02459_));
 sky130_as_sc_hs__nand3_2 _33190_ (.A(net352),
    .B(_02460_),
    .C(_02461_),
    .Y(_02462_));
 sky130_as_sc_hs__nand3_2 _33191_ (.A(net231),
    .B(_02459_),
    .C(_02462_),
    .Y(_02463_));
 sky130_as_sc_hs__nand3_2 _33194_ (.A(net352),
    .B(_02464_),
    .C(_02465_),
    .Y(_02466_));
 sky130_as_sc_hs__nand3_2 _33197_ (.A(net212),
    .B(_02467_),
    .C(_02468_),
    .Y(_02469_));
 sky130_as_sc_hs__nand3_2 _33198_ (.A(net342),
    .B(_02466_),
    .C(_02469_),
    .Y(_02470_));
 sky130_as_sc_hs__nand3_2 _33199_ (.A(net240),
    .B(_02463_),
    .C(_02470_),
    .Y(_02471_));
 sky130_as_sc_hs__nand3_2 _33200_ (.A(net337),
    .B(_02449_),
    .C(_02456_),
    .Y(_02472_));
 sky130_as_sc_hs__nand3_2 _33201_ (.A(net246),
    .B(_02471_),
    .C(_02472_),
    .Y(_02473_));
 sky130_as_sc_hs__and2_2 _33202_ (.A(_02442_),
    .B(_02473_),
    .Y(_02474_));
 sky130_as_sc_hs__inv_2 _33203_ (.Y(_02475_),
    .A(_02474_));
 sky130_as_sc_hs__nor2_2 _33204_ (.A(_25869_),
    .B(_02475_),
    .Y(_02476_));
 sky130_as_sc_hs__and2_2 _33205_ (.A(_25869_),
    .B(_02475_),
    .Y(_02477_));
 sky130_as_sc_hs__or2_2 _33206_ (.A(_02476_),
    .B(_02477_),
    .Y(_02478_));
 sky130_as_sc_hs__and2_2 _33209_ (.A(_02479_),
    .B(_02480_),
    .Y(_02481_));
 sky130_as_sc_hs__and2_2 _33210_ (.A(net114),
    .B(net420),
    .Y(_02482_));
 sky130_as_sc_hs__and2_2 _33211_ (.A(net483),
    .B(net473),
    .Y(_02483_));
 sky130_as_sc_hs__and2_2 _33212_ (.A(_23636_),
    .B(net432),
    .Y(_02484_));
 sky130_as_sc_hs__and2_2 _33213_ (.A(net459),
    .B(net422),
    .Y(_02485_));
 sky130_as_sc_hs__or2_2 _33215_ (.A(_02484_),
    .B(_02485_),
    .Y(_02487_));
 sky130_as_sc_hs__and2_2 _33216_ (.A(_02486_),
    .B(_02487_),
    .Y(_02488_));
 sky130_as_sc_hs__or2_2 _33218_ (.A(_02483_),
    .B(_02488_),
    .Y(_02490_));
 sky130_as_sc_hs__and2_2 _33219_ (.A(_02489_),
    .B(_02490_),
    .Y(_02491_));
 sky130_as_sc_hs__or2_2 _33222_ (.A(_02491_),
    .B(_02492_),
    .Y(_02494_));
 sky130_as_sc_hs__and2_2 _33223_ (.A(_02493_),
    .B(_02494_),
    .Y(_02495_));
 sky130_as_sc_hs__or2_2 _33225_ (.A(_02482_),
    .B(_02495_),
    .Y(_02497_));
 sky130_as_sc_hs__and2_2 _33226_ (.A(_02496_),
    .B(_02497_),
    .Y(_02498_));
 sky130_as_sc_hs__or2_2 _33229_ (.A(_02498_),
    .B(_02499_),
    .Y(_02501_));
 sky130_as_sc_hs__and2_2 _33230_ (.A(_02500_),
    .B(_02501_),
    .Y(_02502_));
 sky130_as_sc_hs__or2_2 _33232_ (.A(_02411_),
    .B(_02502_),
    .Y(_02504_));
 sky130_as_sc_hs__and2_2 _33233_ (.A(_02503_),
    .B(_02504_),
    .Y(_02505_));
 sky130_as_sc_hs__or2_2 _33235_ (.A(_02410_),
    .B(_02505_),
    .Y(_02507_));
 sky130_as_sc_hs__and2_2 _33236_ (.A(_02506_),
    .B(_02507_),
    .Y(_02508_));
 sky130_as_sc_hs__or2_2 _33238_ (.A(_02313_),
    .B(_02508_),
    .Y(_02510_));
 sky130_as_sc_hs__and2_2 _33239_ (.A(_02509_),
    .B(_02510_),
    .Y(_02511_));
 sky130_as_sc_hs__or2_2 _33241_ (.A(_02312_),
    .B(_02511_),
    .Y(_02513_));
 sky130_as_sc_hs__and2_2 _33242_ (.A(_02512_),
    .B(_02513_),
    .Y(_02514_));
 sky130_as_sc_hs__or2_2 _33244_ (.A(_02311_),
    .B(_02514_),
    .Y(_02516_));
 sky130_as_sc_hs__and2_2 _33245_ (.A(_02515_),
    .B(_02516_),
    .Y(_02517_));
 sky130_as_sc_hs__or2_2 _33247_ (.A(_02159_),
    .B(_02517_),
    .Y(_02519_));
 sky130_as_sc_hs__and2_2 _33248_ (.A(_02518_),
    .B(_02519_),
    .Y(_02520_));
 sky130_as_sc_hs__or2_2 _33250_ (.A(_02158_),
    .B(_02520_),
    .Y(_02522_));
 sky130_as_sc_hs__and2_2 _33251_ (.A(_02521_),
    .B(_02522_),
    .Y(_02523_));
 sky130_as_sc_hs__or2_2 _33254_ (.A(_02157_),
    .B(_02523_),
    .Y(_02526_));
 sky130_as_sc_hs__and2_2 _33255_ (.A(_02524_),
    .B(_02526_),
    .Y(_02527_));
 sky130_as_sc_hs__and2_2 _33257_ (.A(_02524_),
    .B(_02528_),
    .Y(_02529_));
 sky130_as_sc_hs__and2_2 _33266_ (.A(net467),
    .B(_24545_),
    .Y(_02538_));
 sky130_as_sc_hs__and2_2 _33267_ (.A(net469),
    .B(net455),
    .Y(_02539_));
 sky130_as_sc_hs__or2_2 _33269_ (.A(_02538_),
    .B(_02539_),
    .Y(_02541_));
 sky130_as_sc_hs__and2_2 _33270_ (.A(_02540_),
    .B(_02541_),
    .Y(_02542_));
 sky130_as_sc_hs__and2_2 _33271_ (.A(net470),
    .B(net86),
    .Y(_02543_));
 sky130_as_sc_hs__or2_2 _33273_ (.A(_02542_),
    .B(_02543_),
    .Y(_02545_));
 sky130_as_sc_hs__and2_2 _33274_ (.A(_02544_),
    .B(_02545_),
    .Y(_02546_));
 sky130_as_sc_hs__and2_2 _33275_ (.A(_24229_),
    .B(net456),
    .Y(_02547_));
 sky130_as_sc_hs__nand3_2 _33276_ (.A(_23712_),
    .B(_25033_),
    .C(_25034_),
    .Y(_02548_));
 sky130_as_sc_hs__and2_2 _33278_ (.A(_23598_),
    .B(_02549_),
    .Y(_02550_));
 sky130_as_sc_hs__nand3_2 _33279_ (.A(net112),
    .B(_23598_),
    .C(_02549_),
    .Y(_02551_));
 sky130_as_sc_hs__or2_2 _33280_ (.A(_02548_),
    .B(_02551_),
    .Y(_02552_));
 sky130_as_sc_hs__and2_2 _33282_ (.A(_02552_),
    .B(_02553_),
    .Y(_02554_));
 sky130_as_sc_hs__or2_2 _33284_ (.A(_02547_),
    .B(_02554_),
    .Y(_02556_));
 sky130_as_sc_hs__or2_2 _33286_ (.A(_02166_),
    .B(_02557_),
    .Y(_02558_));
 sky130_as_sc_hs__and2_2 _33288_ (.A(_02558_),
    .B(_02559_),
    .Y(_02560_));
 sky130_as_sc_hs__or2_2 _33290_ (.A(_02546_),
    .B(_02560_),
    .Y(_02562_));
 sky130_as_sc_hs__and2_2 _33291_ (.A(_02561_),
    .B(_02562_),
    .Y(_02563_));
 sky130_as_sc_hs__or2_2 _33293_ (.A(_02537_),
    .B(_02563_),
    .Y(_02565_));
 sky130_as_sc_hs__and2_2 _33294_ (.A(_02564_),
    .B(_02565_),
    .Y(_02566_));
 sky130_as_sc_hs__and2_2 _33297_ (.A(net461),
    .B(net79),
    .Y(_02569_));
 sky130_as_sc_hs__and2_2 _33298_ (.A(net464),
    .B(net453),
    .Y(_02570_));
 sky130_as_sc_hs__and2_2 _33299_ (.A(net462),
    .B(net447),
    .Y(_02571_));
 sky130_as_sc_hs__or2_2 _33300_ (.A(_02570_),
    .B(_02571_),
    .Y(_02572_));
 sky130_as_sc_hs__and2_2 _33302_ (.A(_02572_),
    .B(_02573_),
    .Y(_02574_));
 sky130_as_sc_hs__or2_2 _33304_ (.A(_02569_),
    .B(_02574_),
    .Y(_02576_));
 sky130_as_sc_hs__and2_2 _33305_ (.A(_02575_),
    .B(_02576_),
    .Y(_02577_));
 sky130_as_sc_hs__or2_2 _33307_ (.A(_02568_),
    .B(_02577_),
    .Y(_02579_));
 sky130_as_sc_hs__and2_2 _33308_ (.A(_02578_),
    .B(_02579_),
    .Y(_02580_));
 sky130_as_sc_hs__or2_2 _33310_ (.A(_02567_),
    .B(_02580_),
    .Y(_02582_));
 sky130_as_sc_hs__and2_2 _33311_ (.A(_02581_),
    .B(_02582_),
    .Y(_02583_));
 sky130_as_sc_hs__or2_2 _33313_ (.A(_02566_),
    .B(_02583_),
    .Y(_02585_));
 sky130_as_sc_hs__and2_2 _33314_ (.A(_02584_),
    .B(_02585_),
    .Y(_02586_));
 sky130_as_sc_hs__or2_2 _33316_ (.A(_02536_),
    .B(_02586_),
    .Y(_02588_));
 sky130_as_sc_hs__and2_2 _33317_ (.A(_02587_),
    .B(_02588_),
    .Y(_02589_));
 sky130_as_sc_hs__and2_2 _33320_ (.A(net481),
    .B(net87),
    .Y(_02592_));
 sky130_as_sc_hs__and2_2 _33321_ (.A(_24527_),
    .B(net443),
    .Y(_02593_));
 sky130_as_sc_hs__and2_2 _33322_ (.A(_23674_),
    .B(_24537_),
    .Y(_02594_));
 sky130_as_sc_hs__or2_2 _33323_ (.A(_02593_),
    .B(_02594_),
    .Y(_02595_));
 sky130_as_sc_hs__and2_2 _33325_ (.A(_02595_),
    .B(_02596_),
    .Y(_02597_));
 sky130_as_sc_hs__or2_2 _33327_ (.A(_02592_),
    .B(_02597_),
    .Y(_02599_));
 sky130_as_sc_hs__and2_2 _33328_ (.A(_02598_),
    .B(_02599_),
    .Y(_02600_));
 sky130_as_sc_hs__or2_2 _33331_ (.A(_02600_),
    .B(_02601_),
    .Y(_02603_));
 sky130_as_sc_hs__and2_2 _33332_ (.A(_02602_),
    .B(_02603_),
    .Y(_02604_));
 sky130_as_sc_hs__and2_2 _33333_ (.A(net450),
    .B(net439),
    .Y(_02605_));
 sky130_as_sc_hs__and2_2 _33334_ (.A(net477),
    .B(net449),
    .Y(_02606_));
 sky130_as_sc_hs__and2_2 _33335_ (.A(_24053_),
    .B(net426),
    .Y(_02607_));
 sky130_as_sc_hs__or2_2 _33336_ (.A(_02606_),
    .B(_02607_),
    .Y(_02608_));
 sky130_as_sc_hs__and2_2 _33338_ (.A(_02608_),
    .B(_02609_),
    .Y(_02610_));
 sky130_as_sc_hs__or2_2 _33340_ (.A(_02605_),
    .B(_02610_),
    .Y(_02612_));
 sky130_as_sc_hs__and2_2 _33341_ (.A(_02611_),
    .B(_02612_),
    .Y(_02613_));
 sky130_as_sc_hs__or2_2 _33343_ (.A(_02604_),
    .B(_02613_),
    .Y(_02615_));
 sky130_as_sc_hs__and2_2 _33344_ (.A(_02614_),
    .B(_02615_),
    .Y(_02616_));
 sky130_as_sc_hs__or2_2 _33346_ (.A(_02591_),
    .B(_02616_),
    .Y(_02618_));
 sky130_as_sc_hs__and2_2 _33347_ (.A(_02617_),
    .B(_02618_),
    .Y(_02619_));
 sky130_as_sc_hs__or2_2 _33349_ (.A(_02590_),
    .B(_02619_),
    .Y(_02621_));
 sky130_as_sc_hs__and2_2 _33350_ (.A(_02620_),
    .B(_02621_),
    .Y(_02622_));
 sky130_as_sc_hs__or2_2 _33352_ (.A(_02589_),
    .B(_02622_),
    .Y(_02624_));
 sky130_as_sc_hs__and2_2 _33353_ (.A(_02623_),
    .B(_02624_),
    .Y(_02625_));
 sky130_as_sc_hs__or2_2 _33355_ (.A(_02535_),
    .B(_02625_),
    .Y(_02627_));
 sky130_as_sc_hs__and2_2 _33356_ (.A(_02626_),
    .B(_02627_),
    .Y(_02628_));
 sky130_as_sc_hs__and2_2 _33361_ (.A(net475),
    .B(_24729_),
    .Y(_02633_));
 sky130_as_sc_hs__and2_2 _33362_ (.A(net473),
    .B(net445),
    .Y(_02634_));
 sky130_as_sc_hs__and2_2 _33363_ (.A(_24216_),
    .B(net435),
    .Y(_02635_));
 sky130_as_sc_hs__or2_2 _33364_ (.A(_02634_),
    .B(_02635_),
    .Y(_02636_));
 sky130_as_sc_hs__and2_2 _33366_ (.A(_02636_),
    .B(_02637_),
    .Y(_02638_));
 sky130_as_sc_hs__or2_2 _33368_ (.A(_02633_),
    .B(_02638_),
    .Y(_02640_));
 sky130_as_sc_hs__and2_2 _33369_ (.A(_02639_),
    .B(_02640_),
    .Y(_02641_));
 sky130_as_sc_hs__or2_2 _33371_ (.A(_02632_),
    .B(_02641_),
    .Y(_02643_));
 sky130_as_sc_hs__and2_2 _33372_ (.A(_02642_),
    .B(_02643_),
    .Y(_02644_));
 sky130_as_sc_hs__or2_2 _33374_ (.A(_02631_),
    .B(_02644_),
    .Y(_02646_));
 sky130_as_sc_hs__and2_2 _33375_ (.A(_02645_),
    .B(_02646_),
    .Y(_02647_));
 sky130_as_sc_hs__or2_2 _33378_ (.A(_02647_),
    .B(_02648_),
    .Y(_02650_));
 sky130_as_sc_hs__and2_2 _33379_ (.A(_02649_),
    .B(_02650_),
    .Y(_02651_));
 sky130_as_sc_hs__or2_2 _33383_ (.A(_02652_),
    .B(_02653_),
    .Y(_02655_));
 sky130_as_sc_hs__and2_2 _33384_ (.A(_02654_),
    .B(_02655_),
    .Y(_02656_));
 sky130_as_sc_hs__and2_2 _33385_ (.A(net123),
    .B(_24808_),
    .Y(_02657_));
 sky130_as_sc_hs__or2_2 _33387_ (.A(_02656_),
    .B(_02657_),
    .Y(_02659_));
 sky130_as_sc_hs__and2_2 _33388_ (.A(_02658_),
    .B(_02659_),
    .Y(_02660_));
 sky130_as_sc_hs__and2_2 _33389_ (.A(_24768_),
    .B(net428),
    .Y(_02661_));
 sky130_as_sc_hs__and2_2 _33390_ (.A(_24774_),
    .B(net432),
    .Y(_02662_));
 sky130_as_sc_hs__and2_2 _33391_ (.A(_24256_),
    .B(net441),
    .Y(_02663_));
 sky130_as_sc_hs__or2_2 _33392_ (.A(_02662_),
    .B(_02663_),
    .Y(_02664_));
 sky130_as_sc_hs__and2_2 _33394_ (.A(_02664_),
    .B(_02665_),
    .Y(_02666_));
 sky130_as_sc_hs__or2_2 _33396_ (.A(_02661_),
    .B(_02666_),
    .Y(_02668_));
 sky130_as_sc_hs__and2_2 _33397_ (.A(_02667_),
    .B(_02668_),
    .Y(_02669_));
 sky130_as_sc_hs__or2_2 _33400_ (.A(_02669_),
    .B(_02670_),
    .Y(_02672_));
 sky130_as_sc_hs__and2_2 _33401_ (.A(_02671_),
    .B(_02672_),
    .Y(_02673_));
 sky130_as_sc_hs__or2_2 _33403_ (.A(_02660_),
    .B(_02673_),
    .Y(_02675_));
 sky130_as_sc_hs__and2_2 _33404_ (.A(_02674_),
    .B(_02675_),
    .Y(_02676_));
 sky130_as_sc_hs__or2_2 _33406_ (.A(_02651_),
    .B(_02676_),
    .Y(_02678_));
 sky130_as_sc_hs__and2_2 _33407_ (.A(_02677_),
    .B(_02678_),
    .Y(_02679_));
 sky130_as_sc_hs__or2_2 _33409_ (.A(_02630_),
    .B(_02679_),
    .Y(_02681_));
 sky130_as_sc_hs__and2_2 _33410_ (.A(_02680_),
    .B(_02681_),
    .Y(_02682_));
 sky130_as_sc_hs__or2_2 _33412_ (.A(_02629_),
    .B(_02682_),
    .Y(_02684_));
 sky130_as_sc_hs__and2_2 _33413_ (.A(_02683_),
    .B(_02684_),
    .Y(_02685_));
 sky130_as_sc_hs__or2_2 _33415_ (.A(_02628_),
    .B(_02685_),
    .Y(_02687_));
 sky130_as_sc_hs__and2_2 _33416_ (.A(_02686_),
    .B(_02687_),
    .Y(_02688_));
 sky130_as_sc_hs__or2_2 _33418_ (.A(_02534_),
    .B(_02688_),
    .Y(_02690_));
 sky130_as_sc_hs__and2_2 _33419_ (.A(_02689_),
    .B(_02690_),
    .Y(_02691_));
 sky130_as_sc_hs__and2_2 _33426_ (.A(_25205_),
    .B(net420),
    .Y(_02698_));
 sky130_as_sc_hs__and2_2 _33427_ (.A(_25211_),
    .B(net424),
    .Y(_02699_));
 sky130_as_sc_hs__and2_2 _33428_ (.A(net459),
    .B(net129),
    .Y(_02700_));
 sky130_as_sc_hs__or2_2 _33429_ (.A(_02699_),
    .B(_02700_),
    .Y(_02701_));
 sky130_as_sc_hs__and2_2 _33431_ (.A(_02701_),
    .B(_02702_),
    .Y(_02703_));
 sky130_as_sc_hs__or2_2 _33433_ (.A(_02698_),
    .B(_02703_),
    .Y(_02705_));
 sky130_as_sc_hs__and2_2 _33434_ (.A(_02704_),
    .B(_02705_),
    .Y(_02706_));
 sky130_as_sc_hs__or2_2 _33436_ (.A(_02697_),
    .B(_02706_),
    .Y(_02708_));
 sky130_as_sc_hs__and2_2 _33437_ (.A(_02707_),
    .B(_02708_),
    .Y(_02709_));
 sky130_as_sc_hs__or2_2 _33439_ (.A(_02696_),
    .B(_02709_),
    .Y(_02711_));
 sky130_as_sc_hs__and2_2 _33440_ (.A(_02710_),
    .B(_02711_),
    .Y(_02712_));
 sky130_as_sc_hs__or2_2 _33442_ (.A(_02695_),
    .B(_02712_),
    .Y(_02714_));
 sky130_as_sc_hs__and2_2 _33443_ (.A(_02713_),
    .B(_02714_),
    .Y(_02715_));
 sky130_as_sc_hs__or2_2 _33445_ (.A(_02694_),
    .B(_02715_),
    .Y(_02717_));
 sky130_as_sc_hs__and2_2 _33446_ (.A(_02716_),
    .B(_02717_),
    .Y(_02718_));
 sky130_as_sc_hs__or2_2 _33449_ (.A(_02718_),
    .B(_02719_),
    .Y(_02721_));
 sky130_as_sc_hs__and2_2 _33450_ (.A(_02720_),
    .B(_02721_),
    .Y(_02722_));
 sky130_as_sc_hs__and2_2 _33451_ (.A(_23702_),
    .B(net84),
    .Y(_02723_));
 sky130_as_sc_hs__nand2b_2 _33452_ (.B(_21658_),
    .Y(_02724_),
    .A(_02476_));
 sky130_as_sc_hs__and2_2 _33453_ (.A(_21655_),
    .B(_02724_),
    .Y(_02725_));
 sky130_as_sc_hs__and2_2 _33454_ (.A(net114),
    .B(net75),
    .Y(_02726_));
 sky130_as_sc_hs__and2_2 _33455_ (.A(net482),
    .B(_23643_),
    .Y(_02727_));
 sky130_as_sc_hs__and2_2 _33456_ (.A(_23636_),
    .B(net430),
    .Y(_02728_));
 sky130_as_sc_hs__and2_2 _33457_ (.A(net91),
    .B(net422),
    .Y(_02729_));
 sky130_as_sc_hs__or2_2 _33458_ (.A(_02728_),
    .B(_02729_),
    .Y(_02730_));
 sky130_as_sc_hs__and2_2 _33460_ (.A(_02730_),
    .B(_02731_),
    .Y(_02732_));
 sky130_as_sc_hs__or2_2 _33462_ (.A(_02727_),
    .B(_02732_),
    .Y(_02734_));
 sky130_as_sc_hs__and2_2 _33463_ (.A(_02733_),
    .B(_02734_),
    .Y(_02735_));
 sky130_as_sc_hs__or2_2 _33466_ (.A(_02735_),
    .B(_02736_),
    .Y(_02738_));
 sky130_as_sc_hs__and2_2 _33467_ (.A(_02737_),
    .B(_02738_),
    .Y(_02739_));
 sky130_as_sc_hs__or2_2 _33469_ (.A(_02726_),
    .B(_02739_),
    .Y(_02741_));
 sky130_as_sc_hs__and2_2 _33470_ (.A(_02740_),
    .B(_02741_),
    .Y(_02742_));
 sky130_as_sc_hs__or2_2 _33473_ (.A(_02742_),
    .B(_02743_),
    .Y(_02745_));
 sky130_as_sc_hs__and2_2 _33474_ (.A(_02744_),
    .B(_02745_),
    .Y(_02746_));
 sky130_as_sc_hs__or2_2 _33476_ (.A(_02723_),
    .B(_02746_),
    .Y(_02748_));
 sky130_as_sc_hs__and2_2 _33477_ (.A(_02747_),
    .B(_02748_),
    .Y(_02749_));
 sky130_as_sc_hs__or2_2 _33479_ (.A(_02722_),
    .B(_02749_),
    .Y(_02751_));
 sky130_as_sc_hs__and2_2 _33480_ (.A(_02750_),
    .B(_02751_),
    .Y(_02752_));
 sky130_as_sc_hs__or2_2 _33482_ (.A(_02693_),
    .B(_02752_),
    .Y(_02754_));
 sky130_as_sc_hs__and2_2 _33483_ (.A(_02753_),
    .B(_02754_),
    .Y(_02755_));
 sky130_as_sc_hs__or2_2 _33485_ (.A(_02692_),
    .B(_02755_),
    .Y(_02757_));
 sky130_as_sc_hs__and2_2 _33486_ (.A(_02756_),
    .B(_02757_),
    .Y(_02758_));
 sky130_as_sc_hs__or2_2 _33488_ (.A(_02691_),
    .B(_02758_),
    .Y(_02760_));
 sky130_as_sc_hs__and2_2 _33489_ (.A(_02759_),
    .B(_02760_),
    .Y(_02761_));
 sky130_as_sc_hs__or2_2 _33491_ (.A(_02533_),
    .B(_02761_),
    .Y(_02763_));
 sky130_as_sc_hs__and2_2 _33492_ (.A(_02762_),
    .B(_02763_),
    .Y(_02764_));
 sky130_as_sc_hs__or2_2 _33494_ (.A(_02532_),
    .B(_02764_),
    .Y(_02766_));
 sky130_as_sc_hs__and2_2 _33495_ (.A(_02765_),
    .B(_02766_),
    .Y(_02767_));
 sky130_as_sc_hs__or2_2 _33497_ (.A(_02531_),
    .B(_02767_),
    .Y(_02769_));
 sky130_as_sc_hs__and2_2 _33498_ (.A(_02768_),
    .B(_02769_),
    .Y(_02770_));
 sky130_as_sc_hs__or2_2 _33500_ (.A(_02530_),
    .B(_02770_),
    .Y(_02772_));
 sky130_as_sc_hs__or2_2 _33502_ (.A(_02529_),
    .B(_02773_),
    .Y(_02774_));
 sky130_as_sc_hs__and2_2 _33504_ (.A(_02774_),
    .B(_02775_),
    .Y(_02776_));
 sky130_as_sc_hs__or2_2 _33505_ (.A(_02525_),
    .B(_02527_),
    .Y(_02777_));
 sky130_as_sc_hs__and2_2 _33506_ (.A(_02528_),
    .B(_02777_),
    .Y(_02778_));
 sky130_as_sc_hs__or2_2 _33509_ (.A(_02778_),
    .B(_02779_),
    .Y(_02781_));
 sky130_as_sc_hs__and2_2 _33510_ (.A(_02780_),
    .B(_02781_),
    .Y(_02782_));
 sky130_as_sc_hs__nand3_2 _33512_ (.A(_02156_),
    .B(_02776_),
    .C(_02782_),
    .Y(_02784_));
 sky130_as_sc_hs__or2_2 _33513_ (.A(_02148_),
    .B(_02150_),
    .Y(_02785_));
 sky130_as_sc_hs__or2_2 _33515_ (.A(_01979_),
    .B(_01980_),
    .Y(_02787_));
 sky130_as_sc_hs__and2_2 _33516_ (.A(_01981_),
    .B(_02787_),
    .Y(_02788_));
 sky130_as_sc_hs__or2_2 _33517_ (.A(_01974_),
    .B(_01976_),
    .Y(_02789_));
 sky130_as_sc_hs__and2_2 _33518_ (.A(_01977_),
    .B(_02789_),
    .Y(_02790_));
 sky130_as_sc_hs__and2_2 _33519_ (.A(net464),
    .B(net458),
    .Y(_02791_));
 sky130_as_sc_hs__and2_2 _33520_ (.A(net90),
    .B(net462),
    .Y(_02792_));
 sky130_as_sc_hs__and2_2 _33522_ (.A(_24053_),
    .B(net461),
    .Y(_02794_));
 sky130_as_sc_hs__or2_2 _33523_ (.A(_02791_),
    .B(_02792_),
    .Y(_02795_));
 sky130_as_sc_hs__and2_2 _33524_ (.A(_02793_),
    .B(_02795_),
    .Y(_02796_));
 sky130_as_sc_hs__or2_2 _33528_ (.A(_02790_),
    .B(_02798_),
    .Y(_02800_));
 sky130_as_sc_hs__and2_2 _33529_ (.A(_02799_),
    .B(_02800_),
    .Y(_02801_));
 sky130_as_sc_hs__or2_2 _33531_ (.A(_01970_),
    .B(_01989_),
    .Y(_02803_));
 sky130_as_sc_hs__or2_2 _33533_ (.A(_02802_),
    .B(_02804_),
    .Y(_02805_));
 sky130_as_sc_hs__and2_2 _33535_ (.A(_02805_),
    .B(_02806_),
    .Y(_02807_));
 sky130_as_sc_hs__and2_2 _33536_ (.A(_23712_),
    .B(_24527_),
    .Y(_02808_));
 sky130_as_sc_hs__nand3_2 _33537_ (.A(_24216_),
    .B(_24535_),
    .C(_24536_),
    .Y(_02809_));
 sky130_as_sc_hs__nand3_2 _33538_ (.A(_24216_),
    .B(_24537_),
    .C(_02808_),
    .Y(_02810_));
 sky130_as_sc_hs__and2_2 _33539_ (.A(_24229_),
    .B(net87),
    .Y(_02811_));
 sky130_as_sc_hs__nand2b_2 _33540_ (.B(_02809_),
    .Y(_02812_),
    .A(_02808_));
 sky130_as_sc_hs__and2_2 _33541_ (.A(_02810_),
    .B(_02812_),
    .Y(_02813_));
 sky130_as_sc_hs__or2_2 _33544_ (.A(_01999_),
    .B(_02001_),
    .Y(_02816_));
 sky130_as_sc_hs__and2_2 _33545_ (.A(_02002_),
    .B(_02816_),
    .Y(_02817_));
 sky130_as_sc_hs__or2_2 _33547_ (.A(_02815_),
    .B(_02817_),
    .Y(_02819_));
 sky130_as_sc_hs__and2_2 _33548_ (.A(_02818_),
    .B(_02819_),
    .Y(_02820_));
 sky130_as_sc_hs__or2_2 _33549_ (.A(_02031_),
    .B(_02032_),
    .Y(_02821_));
 sky130_as_sc_hs__and2_2 _33550_ (.A(_02033_),
    .B(_02821_),
    .Y(_02822_));
 sky130_as_sc_hs__or2_2 _33553_ (.A(_02008_),
    .B(_02010_),
    .Y(_02825_));
 sky130_as_sc_hs__or2_2 _33555_ (.A(_02799_),
    .B(_02826_),
    .Y(_02827_));
 sky130_as_sc_hs__and2_2 _33557_ (.A(_02827_),
    .B(_02828_),
    .Y(_02829_));
 sky130_as_sc_hs__or2_2 _33559_ (.A(_02824_),
    .B(_02829_),
    .Y(_02831_));
 sky130_as_sc_hs__and2_2 _33560_ (.A(_02830_),
    .B(_02831_),
    .Y(_02832_));
 sky130_as_sc_hs__or2_2 _33563_ (.A(_01995_),
    .B(_02021_),
    .Y(_02835_));
 sky130_as_sc_hs__and2_2 _33564_ (.A(_02022_),
    .B(_02835_),
    .Y(_02836_));
 sky130_as_sc_hs__or2_2 _33566_ (.A(_02834_),
    .B(_02836_),
    .Y(_02838_));
 sky130_as_sc_hs__and2_2 _33567_ (.A(_02837_),
    .B(_02838_),
    .Y(_02839_));
 sky130_as_sc_hs__and2_2 _33569_ (.A(_02042_),
    .B(_02840_),
    .Y(_02841_));
 sky130_as_sc_hs__and2_2 _33570_ (.A(_24256_),
    .B(net448),
    .Y(_02842_));
 sky130_as_sc_hs__and2_2 _33571_ (.A(_24501_),
    .B(net450),
    .Y(_02843_));
 sky130_as_sc_hs__or2_2 _33573_ (.A(_02037_),
    .B(_02038_),
    .Y(_02845_));
 sky130_as_sc_hs__or2_2 _33575_ (.A(_02844_),
    .B(_02846_),
    .Y(_02847_));
 sky130_as_sc_hs__and2_2 _33576_ (.A(_24545_),
    .B(net445),
    .Y(_02848_));
 sky130_as_sc_hs__and2_2 _33577_ (.A(net85),
    .B(_24729_),
    .Y(_02849_));
 sky130_as_sc_hs__or2_2 _33581_ (.A(_02850_),
    .B(_02852_),
    .Y(_02853_));
 sky130_as_sc_hs__or2_2 _33584_ (.A(_02841_),
    .B(_02854_),
    .Y(_02856_));
 sky130_as_sc_hs__and2_2 _33585_ (.A(_02855_),
    .B(_02856_),
    .Y(_02857_));
 sky130_as_sc_hs__or2_2 _33586_ (.A(_02074_),
    .B(_02076_),
    .Y(_02858_));
 sky130_as_sc_hs__and2_2 _33587_ (.A(_02077_),
    .B(_02858_),
    .Y(_02859_));
 sky130_as_sc_hs__or2_2 _33591_ (.A(_02046_),
    .B(_02048_),
    .Y(_02863_));
 sky130_as_sc_hs__and2_2 _33592_ (.A(_02049_),
    .B(_02863_),
    .Y(_02864_));
 sky130_as_sc_hs__or2_2 _33594_ (.A(_02862_),
    .B(_02864_),
    .Y(_02866_));
 sky130_as_sc_hs__and2_2 _33595_ (.A(_02865_),
    .B(_02866_),
    .Y(_02867_));
 sky130_as_sc_hs__or2_2 _33597_ (.A(_02861_),
    .B(_02867_),
    .Y(_02869_));
 sky130_as_sc_hs__and2_2 _33598_ (.A(_02868_),
    .B(_02869_),
    .Y(_02870_));
 sky130_as_sc_hs__or2_2 _33601_ (.A(_02028_),
    .B(_02059_),
    .Y(_02873_));
 sky130_as_sc_hs__and2_2 _33602_ (.A(_02060_),
    .B(_02873_),
    .Y(_02874_));
 sky130_as_sc_hs__or2_2 _33604_ (.A(_02872_),
    .B(_02874_),
    .Y(_02876_));
 sky130_as_sc_hs__and2_2 _33605_ (.A(_02875_),
    .B(_02876_),
    .Y(_02877_));
 sky130_as_sc_hs__or2_2 _33606_ (.A(_02094_),
    .B(_02096_),
    .Y(_02878_));
 sky130_as_sc_hs__and2_2 _33607_ (.A(_02097_),
    .B(_02878_),
    .Y(_02879_));
 sky130_as_sc_hs__and2_2 _33608_ (.A(net446),
    .B(_24774_),
    .Y(_02880_));
 sky130_as_sc_hs__and2_2 _33609_ (.A(net442),
    .B(_24768_),
    .Y(_02881_));
 sky130_as_sc_hs__or2_2 _33611_ (.A(_02067_),
    .B(_02068_),
    .Y(_02883_));
 sky130_as_sc_hs__or2_2 _33613_ (.A(_02882_),
    .B(_02884_),
    .Y(_02885_));
 sky130_as_sc_hs__or2_2 _33614_ (.A(_02082_),
    .B(_02083_),
    .Y(_02886_));
 sky130_as_sc_hs__and2_2 _33615_ (.A(_02084_),
    .B(_02886_),
    .Y(_02887_));
 sky130_as_sc_hs__and2_2 _33617_ (.A(_02885_),
    .B(_02888_),
    .Y(_02889_));
 sky130_as_sc_hs__and2_2 _33621_ (.A(_02093_),
    .B(_02892_),
    .Y(_02893_));
 sky130_as_sc_hs__and2_2 _33623_ (.A(_23674_),
    .B(_24814_),
    .Y(_02895_));
 sky130_as_sc_hs__and2_2 _33624_ (.A(net481),
    .B(_24808_),
    .Y(_02896_));
 sky130_as_sc_hs__or2_2 _33626_ (.A(_02088_),
    .B(_02089_),
    .Y(_02898_));
 sky130_as_sc_hs__or2_2 _33628_ (.A(_02897_),
    .B(_02899_),
    .Y(_02900_));
 sky130_as_sc_hs__and2_2 _33629_ (.A(net477),
    .B(_25211_),
    .Y(_02901_));
 sky130_as_sc_hs__and2_2 _33630_ (.A(net439),
    .B(_25205_),
    .Y(_02902_));
 sky130_as_sc_hs__or2_2 _33634_ (.A(_02903_),
    .B(_02905_),
    .Y(_02906_));
 sky130_as_sc_hs__or2_2 _33636_ (.A(_02891_),
    .B(_02893_),
    .Y(_02908_));
 sky130_as_sc_hs__and2_2 _33637_ (.A(_02894_),
    .B(_02908_),
    .Y(_02909_));
 sky130_as_sc_hs__or2_2 _33641_ (.A(_02879_),
    .B(_02911_),
    .Y(_02913_));
 sky130_as_sc_hs__and2_2 _33642_ (.A(_02912_),
    .B(_02913_),
    .Y(_02914_));
 sky130_as_sc_hs__and2_2 _33643_ (.A(_23702_),
    .B(net443),
    .Y(_02915_));
 sky130_as_sc_hs__or2_2 _33644_ (.A(_02113_),
    .B(_02115_),
    .Y(_02916_));
 sky130_as_sc_hs__and2_2 _33645_ (.A(_02116_),
    .B(_02916_),
    .Y(_02917_));
 sky130_as_sc_hs__or2_2 _33646_ (.A(_02107_),
    .B(_02108_),
    .Y(_02918_));
 sky130_as_sc_hs__and2_2 _33648_ (.A(_23636_),
    .B(net442),
    .Y(_02920_));
 sky130_as_sc_hs__and2_2 _33649_ (.A(net482),
    .B(net85),
    .Y(_02921_));
 sky130_as_sc_hs__or2_2 _33651_ (.A(_02919_),
    .B(_02922_),
    .Y(_02923_));
 sky130_as_sc_hs__and2_2 _33652_ (.A(net114),
    .B(net475),
    .Y(_02924_));
 sky130_as_sc_hs__and2_2 _33654_ (.A(_02923_),
    .B(_02925_),
    .Y(_02926_));
 sky130_as_sc_hs__or2_2 _33658_ (.A(_02917_),
    .B(_02928_),
    .Y(_02930_));
 sky130_as_sc_hs__and2_2 _33659_ (.A(_02929_),
    .B(_02930_),
    .Y(_02931_));
 sky130_as_sc_hs__or2_2 _33661_ (.A(_02915_),
    .B(_02931_),
    .Y(_02933_));
 sky130_as_sc_hs__and2_2 _33662_ (.A(_02932_),
    .B(_02933_),
    .Y(_02934_));
 sky130_as_sc_hs__or2_2 _33666_ (.A(_02103_),
    .B(_02123_),
    .Y(_02938_));
 sky130_as_sc_hs__and2_2 _33667_ (.A(_02124_),
    .B(_02938_),
    .Y(_02939_));
 sky130_as_sc_hs__or2_2 _33669_ (.A(_02937_),
    .B(_02939_),
    .Y(_02941_));
 sky130_as_sc_hs__and2_2 _33670_ (.A(_02940_),
    .B(_02941_),
    .Y(_02942_));
 sky130_as_sc_hs__or2_2 _33672_ (.A(_02936_),
    .B(_02942_),
    .Y(_02944_));
 sky130_as_sc_hs__and2_2 _33673_ (.A(_02943_),
    .B(_02944_),
    .Y(_02945_));
 sky130_as_sc_hs__or2_2 _33676_ (.A(_02066_),
    .B(_02134_),
    .Y(_02948_));
 sky130_as_sc_hs__and2_2 _33677_ (.A(_02135_),
    .B(_02948_),
    .Y(_02949_));
 sky130_as_sc_hs__or2_2 _33680_ (.A(_02947_),
    .B(_02949_),
    .Y(_02952_));
 sky130_as_sc_hs__and2_2 _33681_ (.A(_02950_),
    .B(_02952_),
    .Y(_02953_));
 sky130_as_sc_hs__nand3_2 _33682_ (.A(_02950_),
    .B(_02951_),
    .C(_02952_),
    .Y(_02954_));
 sky130_as_sc_hs__or2_2 _33684_ (.A(_02140_),
    .B(_02142_),
    .Y(_02956_));
 sky130_as_sc_hs__and2_2 _33685_ (.A(_02143_),
    .B(_02956_),
    .Y(_02957_));
 sky130_as_sc_hs__or2_2 _33688_ (.A(_02955_),
    .B(_02957_),
    .Y(_02960_));
 sky130_as_sc_hs__and2_2 _33689_ (.A(_02958_),
    .B(_02960_),
    .Y(_02961_));
 sky130_as_sc_hs__and2_2 _33691_ (.A(_02958_),
    .B(_02962_),
    .Y(_02963_));
 sky130_as_sc_hs__or2_2 _33692_ (.A(_02786_),
    .B(_02963_),
    .Y(_02964_));
 sky130_as_sc_hs__and2_2 _33694_ (.A(_02964_),
    .B(_02965_),
    .Y(_02966_));
 sky130_as_sc_hs__or2_2 _33695_ (.A(_02959_),
    .B(_02961_),
    .Y(_02967_));
 sky130_as_sc_hs__and2_2 _33696_ (.A(_02962_),
    .B(_02967_),
    .Y(_02968_));
 sky130_as_sc_hs__and2_2 _33697_ (.A(net113),
    .B(net470),
    .Y(_02969_));
 sky130_as_sc_hs__and2_2 _33698_ (.A(net462),
    .B(net458),
    .Y(_02970_));
 sky130_as_sc_hs__and2_2 _33699_ (.A(net113),
    .B(_24210_),
    .Y(_02971_));
 sky130_as_sc_hs__and2_2 _33701_ (.A(net90),
    .B(net461),
    .Y(_02973_));
 sky130_as_sc_hs__or2_2 _33702_ (.A(_02970_),
    .B(_02971_),
    .Y(_02974_));
 sky130_as_sc_hs__and2_2 _33703_ (.A(_02972_),
    .B(_02974_),
    .Y(_02975_));
 sky130_as_sc_hs__or2_2 _33706_ (.A(_02794_),
    .B(_02796_),
    .Y(_02978_));
 sky130_as_sc_hs__and2_2 _33707_ (.A(_02797_),
    .B(_02978_),
    .Y(_02979_));
 sky130_as_sc_hs__or2_2 _33709_ (.A(_02977_),
    .B(_02979_),
    .Y(_02981_));
 sky130_as_sc_hs__and2_2 _33710_ (.A(_02980_),
    .B(_02981_),
    .Y(_02982_));
 sky130_as_sc_hs__or2_2 _33712_ (.A(_02788_),
    .B(_02801_),
    .Y(_02984_));
 sky130_as_sc_hs__or2_2 _33714_ (.A(_02983_),
    .B(_02985_),
    .Y(_02986_));
 sky130_as_sc_hs__and2_2 _33716_ (.A(_02986_),
    .B(_02987_),
    .Y(_02988_));
 sky130_as_sc_hs__and2_2 _33717_ (.A(_24053_),
    .B(_24527_),
    .Y(_02989_));
 sky130_as_sc_hs__nand3_2 _33718_ (.A(_23712_),
    .B(_24535_),
    .C(_24536_),
    .Y(_02990_));
 sky130_as_sc_hs__nand3_2 _33719_ (.A(_23712_),
    .B(_24537_),
    .C(_02989_),
    .Y(_02991_));
 sky130_as_sc_hs__and2_2 _33720_ (.A(_24216_),
    .B(net87),
    .Y(_02992_));
 sky130_as_sc_hs__nand2b_2 _33721_ (.B(_02990_),
    .Y(_02993_),
    .A(_02989_));
 sky130_as_sc_hs__and2_2 _33722_ (.A(_02991_),
    .B(_02993_),
    .Y(_02994_));
 sky130_as_sc_hs__or2_2 _33725_ (.A(_02811_),
    .B(_02813_),
    .Y(_02997_));
 sky130_as_sc_hs__and2_2 _33726_ (.A(_02814_),
    .B(_02997_),
    .Y(_02998_));
 sky130_as_sc_hs__or2_2 _33728_ (.A(_02996_),
    .B(_02998_),
    .Y(_03000_));
 sky130_as_sc_hs__and2_2 _33729_ (.A(_02999_),
    .B(_03000_),
    .Y(_03001_));
 sky130_as_sc_hs__or2_2 _33730_ (.A(_02842_),
    .B(_02843_),
    .Y(_03002_));
 sky130_as_sc_hs__and2_2 _33731_ (.A(_02844_),
    .B(_03002_),
    .Y(_03003_));
 sky130_as_sc_hs__or2_2 _33734_ (.A(_02820_),
    .B(_02822_),
    .Y(_03006_));
 sky130_as_sc_hs__or2_2 _33736_ (.A(_02980_),
    .B(_03007_),
    .Y(_03008_));
 sky130_as_sc_hs__and2_2 _33738_ (.A(_03008_),
    .B(_03009_),
    .Y(_03010_));
 sky130_as_sc_hs__or2_2 _33740_ (.A(_03005_),
    .B(_03010_),
    .Y(_03012_));
 sky130_as_sc_hs__and2_2 _33741_ (.A(_03011_),
    .B(_03012_),
    .Y(_03013_));
 sky130_as_sc_hs__or2_2 _33744_ (.A(_02807_),
    .B(_02832_),
    .Y(_03016_));
 sky130_as_sc_hs__and2_2 _33745_ (.A(_02833_),
    .B(_03016_),
    .Y(_03017_));
 sky130_as_sc_hs__or2_2 _33747_ (.A(_03015_),
    .B(_03017_),
    .Y(_03019_));
 sky130_as_sc_hs__and2_2 _33748_ (.A(_03018_),
    .B(_03019_),
    .Y(_03020_));
 sky130_as_sc_hs__and2_2 _33750_ (.A(_02853_),
    .B(_03021_),
    .Y(_03022_));
 sky130_as_sc_hs__and2_2 _33751_ (.A(_24256_),
    .B(net450),
    .Y(_03023_));
 sky130_as_sc_hs__and2_2 _33752_ (.A(_24229_),
    .B(net448),
    .Y(_03024_));
 sky130_as_sc_hs__or2_2 _33754_ (.A(_02848_),
    .B(_02849_),
    .Y(_03026_));
 sky130_as_sc_hs__or2_2 _33756_ (.A(_03025_),
    .B(_03027_),
    .Y(_03028_));
 sky130_as_sc_hs__and2_2 _33757_ (.A(net454),
    .B(_24729_),
    .Y(_03029_));
 sky130_as_sc_hs__and2_2 _33758_ (.A(_24501_),
    .B(net444),
    .Y(_03030_));
 sky130_as_sc_hs__or2_2 _33762_ (.A(_03031_),
    .B(_03033_),
    .Y(_03034_));
 sky130_as_sc_hs__or2_2 _33765_ (.A(_03022_),
    .B(_03035_),
    .Y(_03037_));
 sky130_as_sc_hs__and2_2 _33766_ (.A(_03036_),
    .B(_03037_),
    .Y(_03038_));
 sky130_as_sc_hs__or2_2 _33767_ (.A(_02887_),
    .B(_02889_),
    .Y(_03039_));
 sky130_as_sc_hs__and2_2 _33768_ (.A(_02890_),
    .B(_03039_),
    .Y(_03040_));
 sky130_as_sc_hs__or2_2 _33772_ (.A(_02857_),
    .B(_02859_),
    .Y(_03044_));
 sky130_as_sc_hs__and2_2 _33773_ (.A(_02860_),
    .B(_03044_),
    .Y(_03045_));
 sky130_as_sc_hs__or2_2 _33775_ (.A(_03043_),
    .B(_03045_),
    .Y(_03047_));
 sky130_as_sc_hs__and2_2 _33776_ (.A(_03046_),
    .B(_03047_),
    .Y(_03048_));
 sky130_as_sc_hs__or2_2 _33778_ (.A(_03042_),
    .B(_03048_),
    .Y(_03050_));
 sky130_as_sc_hs__and2_2 _33779_ (.A(_03049_),
    .B(_03050_),
    .Y(_03051_));
 sky130_as_sc_hs__or2_2 _33782_ (.A(_02839_),
    .B(_02870_),
    .Y(_03054_));
 sky130_as_sc_hs__and2_2 _33783_ (.A(_02871_),
    .B(_03054_),
    .Y(_03055_));
 sky130_as_sc_hs__or2_2 _33785_ (.A(_03053_),
    .B(_03055_),
    .Y(_03057_));
 sky130_as_sc_hs__and2_2 _33786_ (.A(_03056_),
    .B(_03057_),
    .Y(_03058_));
 sky130_as_sc_hs__and2_2 _33787_ (.A(net79),
    .B(_24768_),
    .Y(_03059_));
 sky130_as_sc_hs__and2_2 _33788_ (.A(net453),
    .B(_24774_),
    .Y(_03060_));
 sky130_as_sc_hs__or2_2 _33790_ (.A(_02880_),
    .B(_02881_),
    .Y(_03062_));
 sky130_as_sc_hs__or2_2 _33792_ (.A(_03061_),
    .B(_03063_),
    .Y(_03064_));
 sky130_as_sc_hs__or2_2 _33793_ (.A(_02895_),
    .B(_02896_),
    .Y(_03065_));
 sky130_as_sc_hs__and2_2 _33794_ (.A(_02897_),
    .B(_03065_),
    .Y(_03066_));
 sky130_as_sc_hs__and2_2 _33796_ (.A(_03064_),
    .B(_03067_),
    .Y(_03068_));
 sky130_as_sc_hs__and2_2 _33800_ (.A(_02906_),
    .B(_03071_),
    .Y(_03072_));
 sky130_as_sc_hs__and2_2 _33802_ (.A(_23674_),
    .B(_24808_),
    .Y(_03074_));
 sky130_as_sc_hs__and2_2 _33803_ (.A(net443),
    .B(_24814_),
    .Y(_03075_));
 sky130_as_sc_hs__or2_2 _33805_ (.A(_02901_),
    .B(_02902_),
    .Y(_03077_));
 sky130_as_sc_hs__or2_2 _33807_ (.A(_03076_),
    .B(_03078_),
    .Y(_03079_));
 sky130_as_sc_hs__and2_2 _33808_ (.A(net477),
    .B(_25205_),
    .Y(_03080_));
 sky130_as_sc_hs__and2_2 _33809_ (.A(net481),
    .B(_25211_),
    .Y(_03081_));
 sky130_as_sc_hs__or2_2 _33813_ (.A(_03082_),
    .B(_03084_),
    .Y(_03085_));
 sky130_as_sc_hs__or2_2 _33815_ (.A(_03070_),
    .B(_03072_),
    .Y(_03087_));
 sky130_as_sc_hs__and2_2 _33816_ (.A(_03073_),
    .B(_03087_),
    .Y(_03088_));
 sky130_as_sc_hs__or2_2 _33819_ (.A(_02907_),
    .B(_02909_),
    .Y(_03091_));
 sky130_as_sc_hs__and2_2 _33820_ (.A(_02910_),
    .B(_03091_),
    .Y(_03092_));
 sky130_as_sc_hs__or2_2 _33822_ (.A(_03090_),
    .B(_03092_),
    .Y(_03094_));
 sky130_as_sc_hs__and2_2 _33823_ (.A(_03093_),
    .B(_03094_),
    .Y(_03095_));
 sky130_as_sc_hs__and2_2 _33824_ (.A(_23702_),
    .B(net79),
    .Y(_03096_));
 sky130_as_sc_hs__or2_2 _33825_ (.A(_02924_),
    .B(_02926_),
    .Y(_03097_));
 sky130_as_sc_hs__and2_2 _33826_ (.A(_02927_),
    .B(_03097_),
    .Y(_03098_));
 sky130_as_sc_hs__or2_2 _33827_ (.A(_02920_),
    .B(_02921_),
    .Y(_03099_));
 sky130_as_sc_hs__and2_2 _33829_ (.A(_23636_),
    .B(net78),
    .Y(_03101_));
 sky130_as_sc_hs__and2_2 _33830_ (.A(net483),
    .B(net454),
    .Y(_03102_));
 sky130_as_sc_hs__or2_2 _33832_ (.A(_03100_),
    .B(_03103_),
    .Y(_03104_));
 sky130_as_sc_hs__and2_2 _33833_ (.A(net115),
    .B(net479),
    .Y(_03105_));
 sky130_as_sc_hs__and2_2 _33835_ (.A(_03104_),
    .B(_03106_),
    .Y(_03107_));
 sky130_as_sc_hs__or2_2 _33839_ (.A(_03098_),
    .B(_03109_),
    .Y(_03111_));
 sky130_as_sc_hs__and2_2 _33840_ (.A(_03110_),
    .B(_03111_),
    .Y(_03112_));
 sky130_as_sc_hs__or2_2 _33842_ (.A(_03096_),
    .B(_03112_),
    .Y(_03114_));
 sky130_as_sc_hs__and2_2 _33843_ (.A(_03113_),
    .B(_03114_),
    .Y(_03115_));
 sky130_as_sc_hs__or2_2 _33847_ (.A(_02914_),
    .B(_02934_),
    .Y(_03119_));
 sky130_as_sc_hs__and2_2 _33848_ (.A(_02935_),
    .B(_03119_),
    .Y(_03120_));
 sky130_as_sc_hs__or2_2 _33850_ (.A(_03118_),
    .B(_03120_),
    .Y(_03122_));
 sky130_as_sc_hs__and2_2 _33851_ (.A(_03121_),
    .B(_03122_),
    .Y(_03123_));
 sky130_as_sc_hs__or2_2 _33853_ (.A(_03117_),
    .B(_03123_),
    .Y(_03125_));
 sky130_as_sc_hs__and2_2 _33854_ (.A(_03124_),
    .B(_03125_),
    .Y(_03126_));
 sky130_as_sc_hs__or2_2 _33857_ (.A(_02877_),
    .B(_02945_),
    .Y(_03129_));
 sky130_as_sc_hs__and2_2 _33858_ (.A(_02946_),
    .B(_03129_),
    .Y(_03130_));
 sky130_as_sc_hs__or2_2 _33861_ (.A(_03128_),
    .B(_03130_),
    .Y(_03133_));
 sky130_as_sc_hs__and2_2 _33862_ (.A(_03131_),
    .B(_03133_),
    .Y(_03134_));
 sky130_as_sc_hs__or2_2 _33865_ (.A(_02951_),
    .B(_02953_),
    .Y(_03137_));
 sky130_as_sc_hs__and2_2 _33866_ (.A(_02954_),
    .B(_03137_),
    .Y(_03138_));
 sky130_as_sc_hs__or2_2 _33869_ (.A(_03136_),
    .B(_03138_),
    .Y(_03141_));
 sky130_as_sc_hs__and2_2 _33870_ (.A(_03139_),
    .B(_03141_),
    .Y(_03142_));
 sky130_as_sc_hs__nand3_2 _33871_ (.A(_03139_),
    .B(_03140_),
    .C(_03141_),
    .Y(_03143_));
 sky130_as_sc_hs__or2_2 _33874_ (.A(_02968_),
    .B(_03144_),
    .Y(_03146_));
 sky130_as_sc_hs__and2_2 _33875_ (.A(_03145_),
    .B(_03146_),
    .Y(_03147_));
 sky130_as_sc_hs__and2_2 _33876_ (.A(_02966_),
    .B(_03147_),
    .Y(_03148_));
 sky130_as_sc_hs__or2_2 _33878_ (.A(_02969_),
    .B(_02982_),
    .Y(_03150_));
 sky130_as_sc_hs__and2_2 _33879_ (.A(_02983_),
    .B(_03150_),
    .Y(_03151_));
 sky130_as_sc_hs__nand3_2 _33880_ (.A(_24053_),
    .B(_24535_),
    .C(_24536_),
    .Y(_03152_));
 sky130_as_sc_hs__or2_2 _33882_ (.A(_03152_),
    .B(_03153_),
    .Y(_03154_));
 sky130_as_sc_hs__and2_2 _33883_ (.A(_23712_),
    .B(net87),
    .Y(_03155_));
 sky130_as_sc_hs__and2_2 _33885_ (.A(_03154_),
    .B(_03156_),
    .Y(_03157_));
 sky130_as_sc_hs__or2_2 _33888_ (.A(_02992_),
    .B(_02994_),
    .Y(_03160_));
 sky130_as_sc_hs__and2_2 _33889_ (.A(_02995_),
    .B(_03160_),
    .Y(_03161_));
 sky130_as_sc_hs__or2_2 _33891_ (.A(_03023_),
    .B(_03024_),
    .Y(_03163_));
 sky130_as_sc_hs__and2_2 _33892_ (.A(_03025_),
    .B(_03163_),
    .Y(_03164_));
 sky130_as_sc_hs__or2_2 _33893_ (.A(_03159_),
    .B(_03161_),
    .Y(_03165_));
 sky130_as_sc_hs__and2_2 _33894_ (.A(_03162_),
    .B(_03165_),
    .Y(_03166_));
 sky130_as_sc_hs__or2_2 _33897_ (.A(_02973_),
    .B(_02975_),
    .Y(_03169_));
 sky130_as_sc_hs__and2_2 _33898_ (.A(_02976_),
    .B(_03169_),
    .Y(_03170_));
 sky130_as_sc_hs__and2_2 _33899_ (.A(net113),
    .B(net462),
    .Y(_03171_));
 sky130_as_sc_hs__and2_2 _33900_ (.A(net461),
    .B(net458),
    .Y(_03172_));
 sky130_as_sc_hs__inv_2 _33902_ (.Y(_03174_),
    .A(_03173_));
 sky130_as_sc_hs__or2_2 _33904_ (.A(_03001_),
    .B(_03003_),
    .Y(_03176_));
 sky130_as_sc_hs__or2_2 _33906_ (.A(_03175_),
    .B(_03177_),
    .Y(_03178_));
 sky130_as_sc_hs__and2_2 _33908_ (.A(_03178_),
    .B(_03179_),
    .Y(_03180_));
 sky130_as_sc_hs__or2_2 _33910_ (.A(_03168_),
    .B(_03180_),
    .Y(_03182_));
 sky130_as_sc_hs__and2_2 _33911_ (.A(_03181_),
    .B(_03182_),
    .Y(_03183_));
 sky130_as_sc_hs__or2_2 _33913_ (.A(_02988_),
    .B(_03013_),
    .Y(_03185_));
 sky130_as_sc_hs__or2_2 _33915_ (.A(_03184_),
    .B(_03186_),
    .Y(_03187_));
 sky130_as_sc_hs__and2_2 _33917_ (.A(_03187_),
    .B(_03188_),
    .Y(_03189_));
 sky130_as_sc_hs__and2_2 _33919_ (.A(_03034_),
    .B(_03190_),
    .Y(_03191_));
 sky130_as_sc_hs__and2_2 _33920_ (.A(_24229_),
    .B(net451),
    .Y(_03192_));
 sky130_as_sc_hs__and2_2 _33921_ (.A(_24216_),
    .B(net448),
    .Y(_03193_));
 sky130_as_sc_hs__or2_2 _33923_ (.A(_03029_),
    .B(_03030_),
    .Y(_03195_));
 sky130_as_sc_hs__or2_2 _33925_ (.A(_03194_),
    .B(_03196_),
    .Y(_03197_));
 sky130_as_sc_hs__and2_2 _33928_ (.A(_24545_),
    .B(_24729_),
    .Y(_03200_));
 sky130_as_sc_hs__and2_2 _33929_ (.A(_24256_),
    .B(net444),
    .Y(_03201_));
 sky130_as_sc_hs__or2_2 _33931_ (.A(_03199_),
    .B(_03202_),
    .Y(_03203_));
 sky130_as_sc_hs__or2_2 _33934_ (.A(_03191_),
    .B(_03204_),
    .Y(_03206_));
 sky130_as_sc_hs__and2_2 _33935_ (.A(_03205_),
    .B(_03206_),
    .Y(_03207_));
 sky130_as_sc_hs__or2_2 _33936_ (.A(_03066_),
    .B(_03068_),
    .Y(_03208_));
 sky130_as_sc_hs__and2_2 _33937_ (.A(_03069_),
    .B(_03208_),
    .Y(_03209_));
 sky130_as_sc_hs__or2_2 _33941_ (.A(_03038_),
    .B(_03040_),
    .Y(_03213_));
 sky130_as_sc_hs__and2_2 _33942_ (.A(_03041_),
    .B(_03213_),
    .Y(_03214_));
 sky130_as_sc_hs__or2_2 _33944_ (.A(_03212_),
    .B(_03214_),
    .Y(_03216_));
 sky130_as_sc_hs__and2_2 _33945_ (.A(_03215_),
    .B(_03216_),
    .Y(_03217_));
 sky130_as_sc_hs__or2_2 _33947_ (.A(_03211_),
    .B(_03217_),
    .Y(_03219_));
 sky130_as_sc_hs__and2_2 _33948_ (.A(_03218_),
    .B(_03219_),
    .Y(_03220_));
 sky130_as_sc_hs__or2_2 _33951_ (.A(_03020_),
    .B(_03051_),
    .Y(_03223_));
 sky130_as_sc_hs__and2_2 _33952_ (.A(_03052_),
    .B(_03223_),
    .Y(_03224_));
 sky130_as_sc_hs__or2_2 _33954_ (.A(_03222_),
    .B(_03224_),
    .Y(_03226_));
 sky130_as_sc_hs__and2_2 _33955_ (.A(_03225_),
    .B(_03226_),
    .Y(_03227_));
 sky130_as_sc_hs__or2_2 _33956_ (.A(_03059_),
    .B(_03060_),
    .Y(_03228_));
 sky130_as_sc_hs__and2_2 _33958_ (.A(net447),
    .B(_24768_),
    .Y(_03230_));
 sky130_as_sc_hs__and2_2 _33959_ (.A(net85),
    .B(_24774_),
    .Y(_03231_));
 sky130_as_sc_hs__or2_2 _33961_ (.A(_03229_),
    .B(_03232_),
    .Y(_03233_));
 sky130_as_sc_hs__and2_2 _33963_ (.A(_03233_),
    .B(_03234_),
    .Y(_03235_));
 sky130_as_sc_hs__or2_2 _33964_ (.A(_03074_),
    .B(_03075_),
    .Y(_03236_));
 sky130_as_sc_hs__and2_2 _33965_ (.A(_03076_),
    .B(_03236_),
    .Y(_03237_));
 sky130_as_sc_hs__and2_2 _33969_ (.A(_03085_),
    .B(_03240_),
    .Y(_03241_));
 sky130_as_sc_hs__or2_2 _33971_ (.A(_03080_),
    .B(_03081_),
    .Y(_03243_));
 sky130_as_sc_hs__and2_2 _33973_ (.A(net443),
    .B(_24808_),
    .Y(_03245_));
 sky130_as_sc_hs__and2_2 _33974_ (.A(net79),
    .B(_24814_),
    .Y(_03246_));
 sky130_as_sc_hs__or2_2 _33976_ (.A(_03244_),
    .B(_03247_),
    .Y(_03248_));
 sky130_as_sc_hs__and2_2 _33979_ (.A(net481),
    .B(_25205_),
    .Y(_03251_));
 sky130_as_sc_hs__and2_2 _33980_ (.A(_23674_),
    .B(_25211_),
    .Y(_03252_));
 sky130_as_sc_hs__or2_2 _33982_ (.A(_03250_),
    .B(_03253_),
    .Y(_03254_));
 sky130_as_sc_hs__or2_2 _33984_ (.A(_03239_),
    .B(_03241_),
    .Y(_03256_));
 sky130_as_sc_hs__and2_2 _33985_ (.A(_03242_),
    .B(_03256_),
    .Y(_03257_));
 sky130_as_sc_hs__or2_2 _33988_ (.A(_03086_),
    .B(_03088_),
    .Y(_03260_));
 sky130_as_sc_hs__and2_2 _33989_ (.A(_03089_),
    .B(_03260_),
    .Y(_03261_));
 sky130_as_sc_hs__or2_2 _33991_ (.A(_03259_),
    .B(_03261_),
    .Y(_03263_));
 sky130_as_sc_hs__and2_2 _33992_ (.A(_03262_),
    .B(_03263_),
    .Y(_03264_));
 sky130_as_sc_hs__and2_2 _33993_ (.A(_23702_),
    .B(net447),
    .Y(_03265_));
 sky130_as_sc_hs__or2_2 _33994_ (.A(_03105_),
    .B(_03107_),
    .Y(_03266_));
 sky130_as_sc_hs__and2_2 _33995_ (.A(_03108_),
    .B(_03266_),
    .Y(_03267_));
 sky130_as_sc_hs__or2_2 _33996_ (.A(_03101_),
    .B(_03102_),
    .Y(_03268_));
 sky130_as_sc_hs__and2_2 _33998_ (.A(net482),
    .B(_24545_),
    .Y(_03270_));
 sky130_as_sc_hs__and2_2 _33999_ (.A(_23636_),
    .B(net446),
    .Y(_03271_));
 sky130_as_sc_hs__or2_2 _34001_ (.A(_03269_),
    .B(_03272_),
    .Y(_03273_));
 sky130_as_sc_hs__and2_2 _34002_ (.A(net114),
    .B(net473),
    .Y(_03274_));
 sky130_as_sc_hs__and2_2 _34004_ (.A(_03273_),
    .B(_03275_),
    .Y(_03276_));
 sky130_as_sc_hs__or2_2 _34008_ (.A(_03267_),
    .B(_03278_),
    .Y(_03280_));
 sky130_as_sc_hs__and2_2 _34009_ (.A(_03279_),
    .B(_03280_),
    .Y(_03281_));
 sky130_as_sc_hs__or2_2 _34011_ (.A(_03265_),
    .B(_03281_),
    .Y(_03283_));
 sky130_as_sc_hs__and2_2 _34012_ (.A(_03282_),
    .B(_03283_),
    .Y(_03284_));
 sky130_as_sc_hs__or2_2 _34016_ (.A(_03095_),
    .B(_03115_),
    .Y(_03288_));
 sky130_as_sc_hs__and2_2 _34017_ (.A(_03116_),
    .B(_03288_),
    .Y(_03289_));
 sky130_as_sc_hs__or2_2 _34019_ (.A(_03287_),
    .B(_03289_),
    .Y(_03291_));
 sky130_as_sc_hs__and2_2 _34020_ (.A(_03290_),
    .B(_03291_),
    .Y(_03292_));
 sky130_as_sc_hs__or2_2 _34022_ (.A(_03286_),
    .B(_03292_),
    .Y(_03294_));
 sky130_as_sc_hs__and2_2 _34023_ (.A(_03293_),
    .B(_03294_),
    .Y(_03295_));
 sky130_as_sc_hs__or2_2 _34026_ (.A(_03058_),
    .B(_03126_),
    .Y(_03298_));
 sky130_as_sc_hs__and2_2 _34027_ (.A(_03127_),
    .B(_03298_),
    .Y(_03299_));
 sky130_as_sc_hs__or2_2 _34030_ (.A(_03297_),
    .B(_03299_),
    .Y(_03302_));
 sky130_as_sc_hs__and2_2 _34031_ (.A(_03300_),
    .B(_03302_),
    .Y(_03303_));
 sky130_as_sc_hs__or2_2 _34034_ (.A(_03132_),
    .B(_03134_),
    .Y(_03306_));
 sky130_as_sc_hs__and2_2 _34035_ (.A(_03135_),
    .B(_03306_),
    .Y(_03307_));
 sky130_as_sc_hs__or2_2 _34037_ (.A(_03305_),
    .B(_03307_),
    .Y(_03309_));
 sky130_as_sc_hs__and2_2 _34038_ (.A(_03308_),
    .B(_03309_),
    .Y(_03310_));
 sky130_as_sc_hs__or2_2 _34040_ (.A(_03149_),
    .B(_03310_),
    .Y(_03312_));
 sky130_as_sc_hs__and2_2 _34041_ (.A(_03311_),
    .B(_03312_),
    .Y(_03313_));
 sky130_as_sc_hs__or2_2 _34042_ (.A(_03151_),
    .B(_03183_),
    .Y(_03314_));
 sky130_as_sc_hs__or2_2 _34044_ (.A(_03170_),
    .B(_03174_),
    .Y(_03316_));
 sky130_as_sc_hs__and2_2 _34045_ (.A(_03175_),
    .B(_03316_),
    .Y(_03317_));
 sky130_as_sc_hs__or2_2 _34046_ (.A(_03164_),
    .B(_03166_),
    .Y(_03318_));
 sky130_as_sc_hs__and2_2 _34047_ (.A(_03167_),
    .B(_03318_),
    .Y(_03319_));
 sky130_as_sc_hs__nand3_2 _34048_ (.A(net90),
    .B(_24535_),
    .C(_24536_),
    .Y(_03320_));
 sky130_as_sc_hs__or2_2 _34050_ (.A(_03320_),
    .B(_03321_),
    .Y(_03322_));
 sky130_as_sc_hs__and2_2 _34051_ (.A(_24053_),
    .B(net87),
    .Y(_03323_));
 sky130_as_sc_hs__and2_2 _34053_ (.A(_03322_),
    .B(_03324_),
    .Y(_03325_));
 sky130_as_sc_hs__or2_2 _34056_ (.A(_03155_),
    .B(_03157_),
    .Y(_03328_));
 sky130_as_sc_hs__and2_2 _34057_ (.A(_03158_),
    .B(_03328_),
    .Y(_03329_));
 sky130_as_sc_hs__or2_2 _34059_ (.A(_03192_),
    .B(_03193_),
    .Y(_03331_));
 sky130_as_sc_hs__and2_2 _34060_ (.A(_03194_),
    .B(_03331_),
    .Y(_03332_));
 sky130_as_sc_hs__or2_2 _34061_ (.A(_03327_),
    .B(_03329_),
    .Y(_03333_));
 sky130_as_sc_hs__and2_2 _34062_ (.A(_03330_),
    .B(_03333_),
    .Y(_03334_));
 sky130_as_sc_hs__or2_2 _34066_ (.A(_03319_),
    .B(_03336_),
    .Y(_03338_));
 sky130_as_sc_hs__and2_2 _34067_ (.A(_03337_),
    .B(_03338_),
    .Y(_03339_));
 sky130_as_sc_hs__or2_2 _34069_ (.A(_03315_),
    .B(_03340_),
    .Y(_03341_));
 sky130_as_sc_hs__and2_2 _34071_ (.A(_03341_),
    .B(_03342_),
    .Y(_03343_));
 sky130_as_sc_hs__and2_2 _34073_ (.A(_03203_),
    .B(_03344_),
    .Y(_03345_));
 sky130_as_sc_hs__or2_2 _34074_ (.A(_03200_),
    .B(_03201_),
    .Y(_03346_));
 sky130_as_sc_hs__and2_2 _34076_ (.A(_23712_),
    .B(net449),
    .Y(_03348_));
 sky130_as_sc_hs__and2_2 _34077_ (.A(_24216_),
    .B(_24585_),
    .Y(_03349_));
 sky130_as_sc_hs__or2_2 _34079_ (.A(_03347_),
    .B(_03350_),
    .Y(_03351_));
 sky130_as_sc_hs__and2_2 _34082_ (.A(_24229_),
    .B(net445),
    .Y(_03354_));
 sky130_as_sc_hs__and2_2 _34083_ (.A(_24501_),
    .B(_24729_),
    .Y(_03355_));
 sky130_as_sc_hs__or2_2 _34085_ (.A(_03353_),
    .B(_03356_),
    .Y(_03357_));
 sky130_as_sc_hs__or2_2 _34088_ (.A(_03345_),
    .B(_03358_),
    .Y(_03360_));
 sky130_as_sc_hs__and2_2 _34089_ (.A(_03359_),
    .B(_03360_),
    .Y(_03361_));
 sky130_as_sc_hs__or2_2 _34090_ (.A(_03235_),
    .B(_03237_),
    .Y(_03362_));
 sky130_as_sc_hs__and2_2 _34091_ (.A(_03238_),
    .B(_03362_),
    .Y(_03363_));
 sky130_as_sc_hs__or2_2 _34094_ (.A(_03207_),
    .B(_03209_),
    .Y(_03366_));
 sky130_as_sc_hs__or2_2 _34096_ (.A(_03337_),
    .B(_03367_),
    .Y(_03368_));
 sky130_as_sc_hs__and2_2 _34098_ (.A(_03368_),
    .B(_03369_),
    .Y(_03370_));
 sky130_as_sc_hs__or2_2 _34100_ (.A(_03365_),
    .B(_03370_),
    .Y(_03372_));
 sky130_as_sc_hs__and2_2 _34101_ (.A(_03371_),
    .B(_03372_),
    .Y(_03373_));
 sky130_as_sc_hs__or2_2 _34104_ (.A(_03189_),
    .B(_03220_),
    .Y(_03376_));
 sky130_as_sc_hs__and2_2 _34105_ (.A(_03221_),
    .B(_03376_),
    .Y(_03377_));
 sky130_as_sc_hs__or2_2 _34107_ (.A(_03375_),
    .B(_03377_),
    .Y(_03379_));
 sky130_as_sc_hs__and2_2 _34108_ (.A(_03378_),
    .B(_03379_),
    .Y(_03380_));
 sky130_as_sc_hs__or2_2 _34109_ (.A(_03255_),
    .B(_03257_),
    .Y(_03381_));
 sky130_as_sc_hs__and2_2 _34110_ (.A(_03258_),
    .B(_03381_),
    .Y(_03382_));
 sky130_as_sc_hs__or2_2 _34111_ (.A(_03230_),
    .B(_03231_),
    .Y(_03383_));
 sky130_as_sc_hs__and2_2 _34113_ (.A(net455),
    .B(_24774_),
    .Y(_03385_));
 sky130_as_sc_hs__and2_2 _34114_ (.A(net453),
    .B(_24768_),
    .Y(_03386_));
 sky130_as_sc_hs__or2_2 _34116_ (.A(_03384_),
    .B(_03387_),
    .Y(_03388_));
 sky130_as_sc_hs__and2_2 _34118_ (.A(_03388_),
    .B(_03389_),
    .Y(_03390_));
 sky130_as_sc_hs__or2_2 _34119_ (.A(_03245_),
    .B(_03246_),
    .Y(_03391_));
 sky130_as_sc_hs__and2_2 _34120_ (.A(_03247_),
    .B(_03391_),
    .Y(_03392_));
 sky130_as_sc_hs__and2_2 _34124_ (.A(_03254_),
    .B(_03395_),
    .Y(_03396_));
 sky130_as_sc_hs__or2_2 _34126_ (.A(_03251_),
    .B(_03252_),
    .Y(_03398_));
 sky130_as_sc_hs__and2_2 _34128_ (.A(net79),
    .B(_24808_),
    .Y(_03400_));
 sky130_as_sc_hs__and2_2 _34129_ (.A(net447),
    .B(_24814_),
    .Y(_03401_));
 sky130_as_sc_hs__or2_2 _34131_ (.A(_03399_),
    .B(_03402_),
    .Y(_03403_));
 sky130_as_sc_hs__and2_2 _34134_ (.A(_23674_),
    .B(_25205_),
    .Y(_03406_));
 sky130_as_sc_hs__nand3_2 _34135_ (.A(_24740_),
    .B(_24741_),
    .C(_25211_),
    .Y(_03407_));
 sky130_as_sc_hs__nand3_2 _34136_ (.A(net443),
    .B(_25211_),
    .C(_03406_),
    .Y(_03408_));
 sky130_as_sc_hs__or2_2 _34137_ (.A(_03405_),
    .B(_03408_),
    .Y(_03409_));
 sky130_as_sc_hs__or2_2 _34139_ (.A(_03394_),
    .B(_03396_),
    .Y(_03411_));
 sky130_as_sc_hs__and2_2 _34140_ (.A(_03397_),
    .B(_03411_),
    .Y(_03412_));
 sky130_as_sc_hs__or2_2 _34144_ (.A(_03382_),
    .B(_03414_),
    .Y(_03416_));
 sky130_as_sc_hs__and2_2 _34145_ (.A(_03415_),
    .B(_03416_),
    .Y(_03417_));
 sky130_as_sc_hs__and2_2 _34146_ (.A(_23702_),
    .B(net453),
    .Y(_03418_));
 sky130_as_sc_hs__or2_2 _34147_ (.A(_03274_),
    .B(_03276_),
    .Y(_03419_));
 sky130_as_sc_hs__and2_2 _34148_ (.A(_03277_),
    .B(_03419_),
    .Y(_03420_));
 sky130_as_sc_hs__or2_2 _34149_ (.A(_03270_),
    .B(_03271_),
    .Y(_03421_));
 sky130_as_sc_hs__and2_2 _34151_ (.A(net482),
    .B(_24501_),
    .Y(_03423_));
 sky130_as_sc_hs__and2_2 _34152_ (.A(_23636_),
    .B(net452),
    .Y(_03424_));
 sky130_as_sc_hs__or2_2 _34154_ (.A(_03422_),
    .B(_03425_),
    .Y(_03426_));
 sky130_as_sc_hs__and2_2 _34155_ (.A(net115),
    .B(net439),
    .Y(_03427_));
 sky130_as_sc_hs__and2_2 _34157_ (.A(_03426_),
    .B(_03428_),
    .Y(_03429_));
 sky130_as_sc_hs__or2_2 _34161_ (.A(_03420_),
    .B(_03431_),
    .Y(_03433_));
 sky130_as_sc_hs__and2_2 _34162_ (.A(_03432_),
    .B(_03433_),
    .Y(_03434_));
 sky130_as_sc_hs__or2_2 _34164_ (.A(_03418_),
    .B(_03434_),
    .Y(_03436_));
 sky130_as_sc_hs__and2_2 _34165_ (.A(_03435_),
    .B(_03436_),
    .Y(_03437_));
 sky130_as_sc_hs__or2_2 _34169_ (.A(_03264_),
    .B(_03284_),
    .Y(_03441_));
 sky130_as_sc_hs__and2_2 _34170_ (.A(_03285_),
    .B(_03441_),
    .Y(_03442_));
 sky130_as_sc_hs__or2_2 _34172_ (.A(_03440_),
    .B(_03442_),
    .Y(_03444_));
 sky130_as_sc_hs__and2_2 _34173_ (.A(_03443_),
    .B(_03444_),
    .Y(_03445_));
 sky130_as_sc_hs__or2_2 _34175_ (.A(_03439_),
    .B(_03445_),
    .Y(_03447_));
 sky130_as_sc_hs__and2_2 _34176_ (.A(_03446_),
    .B(_03447_),
    .Y(_03448_));
 sky130_as_sc_hs__or2_2 _34179_ (.A(_03227_),
    .B(_03295_),
    .Y(_03451_));
 sky130_as_sc_hs__and2_2 _34180_ (.A(_03296_),
    .B(_03451_),
    .Y(_03452_));
 sky130_as_sc_hs__or2_2 _34183_ (.A(_03450_),
    .B(_03452_),
    .Y(_03455_));
 sky130_as_sc_hs__and2_2 _34184_ (.A(_03453_),
    .B(_03455_),
    .Y(_03456_));
 sky130_as_sc_hs__or2_2 _34187_ (.A(_03301_),
    .B(_03303_),
    .Y(_03459_));
 sky130_as_sc_hs__and2_2 _34188_ (.A(_03304_),
    .B(_03459_),
    .Y(_03460_));
 sky130_as_sc_hs__or2_2 _34191_ (.A(_03458_),
    .B(_03460_),
    .Y(_03463_));
 sky130_as_sc_hs__and2_2 _34192_ (.A(_03461_),
    .B(_03463_),
    .Y(_03464_));
 sky130_as_sc_hs__or2_2 _34196_ (.A(_03313_),
    .B(_03466_),
    .Y(_03468_));
 sky130_as_sc_hs__and2_2 _34197_ (.A(_03467_),
    .B(_03468_),
    .Y(_03469_));
 sky130_as_sc_hs__or2_2 _34198_ (.A(_03140_),
    .B(_03142_),
    .Y(_03470_));
 sky130_as_sc_hs__and2_2 _34200_ (.A(_03308_),
    .B(_03311_),
    .Y(_03472_));
 sky130_as_sc_hs__or2_2 _34202_ (.A(_03471_),
    .B(_03472_),
    .Y(_03474_));
 sky130_as_sc_hs__and2_2 _34203_ (.A(_03473_),
    .B(_03474_),
    .Y(_03475_));
 sky130_as_sc_hs__nand3_2 _34204_ (.A(_03148_),
    .B(_03469_),
    .C(_03475_),
    .Y(_03476_));
 sky130_as_sc_hs__or2_2 _34205_ (.A(_02784_),
    .B(_03476_),
    .Y(_03477_));
 sky130_as_sc_hs__and2_2 _34206_ (.A(net116),
    .B(net79),
    .Y(_03478_));
 sky130_as_sc_hs__and2_2 _34207_ (.A(_23636_),
    .B(_24256_),
    .Y(_03479_));
 sky130_as_sc_hs__and2_2 _34208_ (.A(net483),
    .B(_24053_),
    .Y(_03480_));
 sky130_as_sc_hs__and2_2 _34210_ (.A(_23636_),
    .B(_24501_),
    .Y(_03482_));
 sky130_as_sc_hs__and2_2 _34211_ (.A(net483),
    .B(_23712_),
    .Y(_03483_));
 sky130_as_sc_hs__or2_2 _34213_ (.A(_03482_),
    .B(_03483_),
    .Y(_03485_));
 sky130_as_sc_hs__or2_2 _34215_ (.A(_03481_),
    .B(_03486_),
    .Y(_03487_));
 sky130_as_sc_hs__and2_2 _34217_ (.A(_03487_),
    .B(_03488_),
    .Y(_03489_));
 sky130_as_sc_hs__or2_2 _34219_ (.A(_03478_),
    .B(_03489_),
    .Y(_03491_));
 sky130_as_sc_hs__and2_2 _34220_ (.A(_03490_),
    .B(_03491_),
    .Y(_03492_));
 sky130_as_sc_hs__and2_2 _34221_ (.A(_23636_),
    .B(_24229_),
    .Y(_03493_));
 sky130_as_sc_hs__and2_2 _34222_ (.A(net483),
    .B(net91),
    .Y(_03494_));
 sky130_as_sc_hs__or2_2 _34224_ (.A(_03479_),
    .B(_03480_),
    .Y(_03496_));
 sky130_as_sc_hs__or2_2 _34226_ (.A(_03495_),
    .B(_03497_),
    .Y(_03498_));
 sky130_as_sc_hs__and2_2 _34227_ (.A(net116),
    .B(net446),
    .Y(_03499_));
 sky130_as_sc_hs__and2_2 _34229_ (.A(_03498_),
    .B(_03500_),
    .Y(_03501_));
 sky130_as_sc_hs__inv_2 _34234_ (.Y(_03506_),
    .A(_03505_));
 sky130_as_sc_hs__or2_2 _34235_ (.A(_03492_),
    .B(_03503_),
    .Y(_03507_));
 sky130_as_sc_hs__and2_2 _34236_ (.A(_03504_),
    .B(_03507_),
    .Y(_03508_));
 sky130_as_sc_hs__and2_2 _34239_ (.A(_24545_),
    .B(_24814_),
    .Y(_03511_));
 sky130_as_sc_hs__and2_2 _34240_ (.A(net455),
    .B(_24808_),
    .Y(_03512_));
 sky130_as_sc_hs__or2_2 _34242_ (.A(_03511_),
    .B(_03512_),
    .Y(_03514_));
 sky130_as_sc_hs__and2_2 _34243_ (.A(_03513_),
    .B(_03514_),
    .Y(_03515_));
 sky130_as_sc_hs__and2_2 _34244_ (.A(_24229_),
    .B(_24774_),
    .Y(_03516_));
 sky130_as_sc_hs__and2_2 _34245_ (.A(_24501_),
    .B(_24768_),
    .Y(_03517_));
 sky130_as_sc_hs__or2_2 _34247_ (.A(_03516_),
    .B(_03517_),
    .Y(_03519_));
 sky130_as_sc_hs__and2_2 _34249_ (.A(_24216_),
    .B(_24774_),
    .Y(_03521_));
 sky130_as_sc_hs__and2_2 _34250_ (.A(_24256_),
    .B(_24768_),
    .Y(_03522_));
 sky130_as_sc_hs__or2_2 _34252_ (.A(_03520_),
    .B(_03523_),
    .Y(_03524_));
 sky130_as_sc_hs__and2_2 _34254_ (.A(_03524_),
    .B(_03525_),
    .Y(_03526_));
 sky130_as_sc_hs__or2_2 _34256_ (.A(_03515_),
    .B(_03526_),
    .Y(_03528_));
 sky130_as_sc_hs__and2_2 _34257_ (.A(_03527_),
    .B(_03528_),
    .Y(_03529_));
 sky130_as_sc_hs__and2_2 _34258_ (.A(net91),
    .B(net445),
    .Y(_03530_));
 sky130_as_sc_hs__and2_2 _34259_ (.A(_23712_),
    .B(_24729_),
    .Y(_03531_));
 sky130_as_sc_hs__and2_2 _34260_ (.A(_03530_),
    .B(_03531_),
    .Y(_03532_));
 sky130_as_sc_hs__or2_2 _34261_ (.A(_03530_),
    .B(_03531_),
    .Y(_03533_));
 sky130_as_sc_hs__nand2b_2 _34262_ (.B(_03533_),
    .Y(_03534_),
    .A(_03532_));
 sky130_as_sc_hs__and2_2 _34263_ (.A(net458),
    .B(net445),
    .Y(_03535_));
 sky130_as_sc_hs__and2_2 _34264_ (.A(_24053_),
    .B(_24729_),
    .Y(_03536_));
 sky130_as_sc_hs__and2_2 _34266_ (.A(net112),
    .B(net445),
    .Y(_03538_));
 sky130_as_sc_hs__and2_2 _34267_ (.A(net90),
    .B(_24729_),
    .Y(_03539_));
 sky130_as_sc_hs__or2_2 _34269_ (.A(_03535_),
    .B(_03536_),
    .Y(_03541_));
 sky130_as_sc_hs__or2_2 _34271_ (.A(_03540_),
    .B(_03542_),
    .Y(_03543_));
 sky130_as_sc_hs__and2_2 _34272_ (.A(_03537_),
    .B(_03543_),
    .Y(_03544_));
 sky130_as_sc_hs__or2_2 _34273_ (.A(_03534_),
    .B(_03544_),
    .Y(_03545_));
 sky130_as_sc_hs__and2_2 _34275_ (.A(_03545_),
    .B(_03546_),
    .Y(_03547_));
 sky130_as_sc_hs__or2_2 _34277_ (.A(_03529_),
    .B(_03547_),
    .Y(_03549_));
 sky130_as_sc_hs__and2_2 _34279_ (.A(_24501_),
    .B(_24814_),
    .Y(_03551_));
 sky130_as_sc_hs__and2_2 _34280_ (.A(_24545_),
    .B(_24808_),
    .Y(_03552_));
 sky130_as_sc_hs__or2_2 _34282_ (.A(_03551_),
    .B(_03552_),
    .Y(_03554_));
 sky130_as_sc_hs__and2_2 _34283_ (.A(_03553_),
    .B(_03554_),
    .Y(_03555_));
 sky130_as_sc_hs__and2_2 _34284_ (.A(_23712_),
    .B(_24774_),
    .Y(_03556_));
 sky130_as_sc_hs__and2_2 _34285_ (.A(_24229_),
    .B(_24768_),
    .Y(_03557_));
 sky130_as_sc_hs__or2_2 _34287_ (.A(_03521_),
    .B(_03522_),
    .Y(_03559_));
 sky130_as_sc_hs__or2_2 _34289_ (.A(_03558_),
    .B(_03560_),
    .Y(_03561_));
 sky130_as_sc_hs__and2_2 _34291_ (.A(_03561_),
    .B(_03562_),
    .Y(_03563_));
 sky130_as_sc_hs__or2_2 _34293_ (.A(_03555_),
    .B(_03563_),
    .Y(_03565_));
 sky130_as_sc_hs__and2_2 _34294_ (.A(_03564_),
    .B(_03565_),
    .Y(_03566_));
 sky130_as_sc_hs__and2_2 _34296_ (.A(_03543_),
    .B(_03567_),
    .Y(_03568_));
 sky130_as_sc_hs__or2_2 _34298_ (.A(_03550_),
    .B(_03569_),
    .Y(_03570_));
 sky130_as_sc_hs__and2_2 _34299_ (.A(net452),
    .B(_25205_),
    .Y(_03571_));
 sky130_as_sc_hs__and2_2 _34300_ (.A(net86),
    .B(_25211_),
    .Y(_03572_));
 sky130_as_sc_hs__or2_2 _34302_ (.A(_03571_),
    .B(_03572_),
    .Y(_03574_));
 sky130_as_sc_hs__or2_2 _34304_ (.A(_03553_),
    .B(_03575_),
    .Y(_03576_));
 sky130_as_sc_hs__and2_2 _34305_ (.A(net86),
    .B(_25205_),
    .Y(_03577_));
 sky130_as_sc_hs__and2_2 _34306_ (.A(net454),
    .B(_25211_),
    .Y(_03578_));
 sky130_as_sc_hs__or2_2 _34310_ (.A(_03579_),
    .B(_03581_),
    .Y(_03582_));
 sky130_as_sc_hs__and2_2 _34313_ (.A(net452),
    .B(_25211_),
    .Y(_03585_));
 sky130_as_sc_hs__and2_2 _34314_ (.A(net447),
    .B(_25205_),
    .Y(_03586_));
 sky130_as_sc_hs__or2_2 _34316_ (.A(_03585_),
    .B(_03586_),
    .Y(_03588_));
 sky130_as_sc_hs__or2_2 _34318_ (.A(_03513_),
    .B(_03589_),
    .Y(_03590_));
 sky130_as_sc_hs__or2_2 _34321_ (.A(_03573_),
    .B(_03592_),
    .Y(_03593_));
 sky130_as_sc_hs__and2_2 _34323_ (.A(_03593_),
    .B(_03594_),
    .Y(_03595_));
 sky130_as_sc_hs__or2_2 _34325_ (.A(_03584_),
    .B(_03595_),
    .Y(_03597_));
 sky130_as_sc_hs__and2_2 _34326_ (.A(_03596_),
    .B(_03597_),
    .Y(_03598_));
 sky130_as_sc_hs__or2_2 _34328_ (.A(_03583_),
    .B(_03598_),
    .Y(_03600_));
 sky130_as_sc_hs__and2_2 _34329_ (.A(_03599_),
    .B(_03600_),
    .Y(_03601_));
 sky130_as_sc_hs__and2_2 _34332_ (.A(_03582_),
    .B(_03603_),
    .Y(_03604_));
 sky130_as_sc_hs__and2_2 _34334_ (.A(_24256_),
    .B(_24814_),
    .Y(_03606_));
 sky130_as_sc_hs__and2_2 _34335_ (.A(_24501_),
    .B(_24808_),
    .Y(_03607_));
 sky130_as_sc_hs__or2_2 _34337_ (.A(_03577_),
    .B(_03578_),
    .Y(_03609_));
 sky130_as_sc_hs__or2_2 _34339_ (.A(_03608_),
    .B(_03610_),
    .Y(_03611_));
 sky130_as_sc_hs__and2_2 _34340_ (.A(net454),
    .B(_25205_),
    .Y(_03612_));
 sky130_as_sc_hs__and2_2 _34341_ (.A(_24545_),
    .B(_25211_),
    .Y(_03613_));
 sky130_as_sc_hs__or2_2 _34345_ (.A(_03614_),
    .B(_03616_),
    .Y(_03617_));
 sky130_as_sc_hs__or2_2 _34347_ (.A(_03602_),
    .B(_03604_),
    .Y(_03619_));
 sky130_as_sc_hs__and2_2 _34348_ (.A(_03605_),
    .B(_03619_),
    .Y(_03620_));
 sky130_as_sc_hs__or2_2 _34352_ (.A(_03601_),
    .B(_03622_),
    .Y(_03624_));
 sky130_as_sc_hs__and2_2 _34353_ (.A(_03623_),
    .B(_03624_),
    .Y(_03625_));
 sky130_as_sc_hs__or2_2 _34354_ (.A(_03506_),
    .B(_03508_),
    .Y(_03626_));
 sky130_as_sc_hs__and2_2 _34355_ (.A(_03509_),
    .B(_03626_),
    .Y(_03627_));
 sky130_as_sc_hs__or2_2 _34357_ (.A(_03625_),
    .B(_03627_),
    .Y(_03629_));
 sky130_as_sc_hs__or2_2 _34359_ (.A(_03570_),
    .B(_03630_),
    .Y(_03631_));
 sky130_as_sc_hs__and2_2 _34361_ (.A(_03631_),
    .B(_03632_),
    .Y(_03633_));
 sky130_as_sc_hs__or2_2 _34362_ (.A(_03618_),
    .B(_03620_),
    .Y(_03634_));
 sky130_as_sc_hs__and2_2 _34363_ (.A(_03621_),
    .B(_03634_),
    .Y(_03635_));
 sky130_as_sc_hs__and2_2 _34364_ (.A(_24053_),
    .B(_24774_),
    .Y(_03636_));
 sky130_as_sc_hs__and2_2 _34365_ (.A(_24216_),
    .B(_24768_),
    .Y(_03637_));
 sky130_as_sc_hs__or2_2 _34367_ (.A(_03556_),
    .B(_03557_),
    .Y(_03639_));
 sky130_as_sc_hs__or2_2 _34369_ (.A(_03638_),
    .B(_03640_),
    .Y(_03641_));
 sky130_as_sc_hs__or2_2 _34370_ (.A(_03606_),
    .B(_03607_),
    .Y(_03642_));
 sky130_as_sc_hs__and2_2 _34371_ (.A(_03608_),
    .B(_03642_),
    .Y(_03643_));
 sky130_as_sc_hs__and2_2 _34373_ (.A(_03641_),
    .B(_03644_),
    .Y(_03645_));
 sky130_as_sc_hs__and2_2 _34377_ (.A(_03617_),
    .B(_03648_),
    .Y(_03649_));
 sky130_as_sc_hs__and2_2 _34379_ (.A(_24229_),
    .B(_24814_),
    .Y(_03651_));
 sky130_as_sc_hs__and2_2 _34380_ (.A(_24256_),
    .B(_24808_),
    .Y(_03652_));
 sky130_as_sc_hs__or2_2 _34382_ (.A(_03612_),
    .B(_03613_),
    .Y(_03654_));
 sky130_as_sc_hs__or2_2 _34384_ (.A(_03653_),
    .B(_03655_),
    .Y(_03656_));
 sky130_as_sc_hs__and2_2 _34387_ (.A(_24545_),
    .B(_25205_),
    .Y(_03659_));
 sky130_as_sc_hs__and2_2 _34388_ (.A(_24501_),
    .B(_25211_),
    .Y(_03660_));
 sky130_as_sc_hs__or2_2 _34390_ (.A(_03658_),
    .B(_03661_),
    .Y(_03662_));
 sky130_as_sc_hs__or2_2 _34392_ (.A(_03647_),
    .B(_03649_),
    .Y(_03664_));
 sky130_as_sc_hs__and2_2 _34393_ (.A(_03650_),
    .B(_03664_),
    .Y(_03665_));
 sky130_as_sc_hs__or2_2 _34397_ (.A(_03635_),
    .B(_03667_),
    .Y(_03669_));
 sky130_as_sc_hs__and2_2 _34398_ (.A(_03668_),
    .B(_03669_),
    .Y(_03670_));
 sky130_as_sc_hs__inv_2 _34400_ (.Y(_03672_),
    .A(_03671_));
 sky130_as_sc_hs__or2_2 _34401_ (.A(_03499_),
    .B(_03501_),
    .Y(_03673_));
 sky130_as_sc_hs__and2_2 _34402_ (.A(_03502_),
    .B(_03673_),
    .Y(_03674_));
 sky130_as_sc_hs__or2_2 _34403_ (.A(_03493_),
    .B(_03494_),
    .Y(_03675_));
 sky130_as_sc_hs__and2_2 _34405_ (.A(_23636_),
    .B(_24216_),
    .Y(_03677_));
 sky130_as_sc_hs__and2_2 _34406_ (.A(net483),
    .B(net459),
    .Y(_03678_));
 sky130_as_sc_hs__or2_2 _34408_ (.A(_03676_),
    .B(_03679_),
    .Y(_03680_));
 sky130_as_sc_hs__and2_2 _34409_ (.A(net116),
    .B(net452),
    .Y(_03681_));
 sky130_as_sc_hs__and2_2 _34411_ (.A(_03680_),
    .B(_03682_),
    .Y(_03683_));
 sky130_as_sc_hs__or2_2 _34415_ (.A(_03674_),
    .B(_03685_),
    .Y(_03687_));
 sky130_as_sc_hs__and2_2 _34416_ (.A(_03686_),
    .B(_03687_),
    .Y(_03688_));
 sky130_as_sc_hs__or2_2 _34418_ (.A(_03672_),
    .B(_03688_),
    .Y(_03690_));
 sky130_as_sc_hs__and2_2 _34419_ (.A(_03689_),
    .B(_03690_),
    .Y(_03691_));
 sky130_as_sc_hs__and2_2 _34424_ (.A(net455),
    .B(_24814_),
    .Y(_03696_));
 sky130_as_sc_hs__and2_2 _34425_ (.A(net86),
    .B(_24808_),
    .Y(_03697_));
 sky130_as_sc_hs__or2_2 _34427_ (.A(_03696_),
    .B(_03697_),
    .Y(_03699_));
 sky130_as_sc_hs__and2_2 _34428_ (.A(_03698_),
    .B(_03699_),
    .Y(_03700_));
 sky130_as_sc_hs__and2_2 _34429_ (.A(_24256_),
    .B(_24774_),
    .Y(_03701_));
 sky130_as_sc_hs__and2_2 _34430_ (.A(_24545_),
    .B(_24768_),
    .Y(_03702_));
 sky130_as_sc_hs__or2_2 _34432_ (.A(_03701_),
    .B(_03702_),
    .Y(_03704_));
 sky130_as_sc_hs__or2_2 _34434_ (.A(_03518_),
    .B(_03705_),
    .Y(_03706_));
 sky130_as_sc_hs__and2_2 _34436_ (.A(_03706_),
    .B(_03707_),
    .Y(_03708_));
 sky130_as_sc_hs__or2_2 _34438_ (.A(_03700_),
    .B(_03708_),
    .Y(_03710_));
 sky130_as_sc_hs__and2_2 _34439_ (.A(_03709_),
    .B(_03710_),
    .Y(_03711_));
 sky130_as_sc_hs__and2_2 _34440_ (.A(net112),
    .B(net448),
    .Y(_03712_));
 sky130_as_sc_hs__and2_2 _34441_ (.A(net459),
    .B(net450),
    .Y(_03713_));
 sky130_as_sc_hs__inv_2 _34443_ (.Y(_03715_),
    .A(_03714_));
 sky130_as_sc_hs__and2_2 _34444_ (.A(_24053_),
    .B(net445),
    .Y(_03716_));
 sky130_as_sc_hs__and2_2 _34445_ (.A(_24216_),
    .B(_24729_),
    .Y(_03717_));
 sky130_as_sc_hs__or2_2 _34447_ (.A(_03716_),
    .B(_03717_),
    .Y(_03719_));
 sky130_as_sc_hs__and2_2 _34448_ (.A(_03718_),
    .B(_03719_),
    .Y(_03720_));
 sky130_as_sc_hs__or2_2 _34450_ (.A(_03715_),
    .B(_03720_),
    .Y(_03722_));
 sky130_as_sc_hs__and2_2 _34451_ (.A(_03721_),
    .B(_03722_),
    .Y(_03723_));
 sky130_as_sc_hs__nor2_2 _34452_ (.A(_03534_),
    .B(_03537_),
    .Y(_03724_));
 sky130_as_sc_hs__or2_2 _34453_ (.A(_03532_),
    .B(_03724_),
    .Y(_03725_));
 sky130_as_sc_hs__or2_2 _34455_ (.A(_03723_),
    .B(_03725_),
    .Y(_03727_));
 sky130_as_sc_hs__and2_2 _34456_ (.A(_03726_),
    .B(_03727_),
    .Y(_03728_));
 sky130_as_sc_hs__or2_2 _34458_ (.A(_03711_),
    .B(_03728_),
    .Y(_03730_));
 sky130_as_sc_hs__and2_2 _34459_ (.A(_03729_),
    .B(_03730_),
    .Y(_03731_));
 sky130_as_sc_hs__or2_2 _34460_ (.A(_03534_),
    .B(_03543_),
    .Y(_03732_));
 sky130_as_sc_hs__and2_2 _34465_ (.A(net447),
    .B(_25211_),
    .Y(_03737_));
 sky130_as_sc_hs__and2_2 _34466_ (.A(net79),
    .B(_25205_),
    .Y(_03738_));
 sky130_as_sc_hs__or2_2 _34468_ (.A(_03737_),
    .B(_03738_),
    .Y(_03740_));
 sky130_as_sc_hs__or2_2 _34470_ (.A(_03698_),
    .B(_03741_),
    .Y(_03742_));
 sky130_as_sc_hs__or2_2 _34473_ (.A(_03587_),
    .B(_03744_),
    .Y(_03745_));
 sky130_as_sc_hs__and2_2 _34475_ (.A(_03745_),
    .B(_03746_),
    .Y(_03747_));
 sky130_as_sc_hs__or2_2 _34477_ (.A(_03736_),
    .B(_03747_),
    .Y(_03749_));
 sky130_as_sc_hs__and2_2 _34478_ (.A(_03748_),
    .B(_03749_),
    .Y(_03750_));
 sky130_as_sc_hs__or2_2 _34480_ (.A(_03735_),
    .B(_03750_),
    .Y(_03752_));
 sky130_as_sc_hs__and2_2 _34481_ (.A(_03751_),
    .B(_03752_),
    .Y(_03753_));
 sky130_as_sc_hs__or2_2 _34484_ (.A(_03753_),
    .B(_03754_),
    .Y(_03756_));
 sky130_as_sc_hs__and2_2 _34485_ (.A(_03755_),
    .B(_03756_),
    .Y(_03757_));
 sky130_as_sc_hs__inv_2 _34487_ (.Y(_03759_),
    .A(_03758_));
 sky130_as_sc_hs__and2_2 _34488_ (.A(net116),
    .B(net442),
    .Y(_03760_));
 sky130_as_sc_hs__and2_2 _34489_ (.A(net482),
    .B(_24216_),
    .Y(_03761_));
 sky130_as_sc_hs__and2_2 _34490_ (.A(_23636_),
    .B(_24545_),
    .Y(_03762_));
 sky130_as_sc_hs__or2_2 _34492_ (.A(_03761_),
    .B(_03762_),
    .Y(_03764_));
 sky130_as_sc_hs__or2_2 _34494_ (.A(_03484_),
    .B(_03765_),
    .Y(_03766_));
 sky130_as_sc_hs__and2_2 _34496_ (.A(_03766_),
    .B(_03767_),
    .Y(_03768_));
 sky130_as_sc_hs__or2_2 _34498_ (.A(_03760_),
    .B(_03768_),
    .Y(_03770_));
 sky130_as_sc_hs__and2_2 _34499_ (.A(_03769_),
    .B(_03770_),
    .Y(_03771_));
 sky130_as_sc_hs__or2_2 _34502_ (.A(_03771_),
    .B(_03772_),
    .Y(_03774_));
 sky130_as_sc_hs__and2_2 _34503_ (.A(_03773_),
    .B(_03774_),
    .Y(_03775_));
 sky130_as_sc_hs__or2_2 _34505_ (.A(_03759_),
    .B(_03775_),
    .Y(_03777_));
 sky130_as_sc_hs__and2_2 _34506_ (.A(_03776_),
    .B(_03777_),
    .Y(_03778_));
 sky130_as_sc_hs__or2_2 _34508_ (.A(_03757_),
    .B(_03778_),
    .Y(_03780_));
 sky130_as_sc_hs__or2_2 _34510_ (.A(_03734_),
    .B(_03781_),
    .Y(_03782_));
 sky130_as_sc_hs__and2_2 _34512_ (.A(_03782_),
    .B(_03783_),
    .Y(_03784_));
 sky130_as_sc_hs__or2_2 _34515_ (.A(_03784_),
    .B(_03785_),
    .Y(_03787_));
 sky130_as_sc_hs__and2_2 _34516_ (.A(_03786_),
    .B(_03787_),
    .Y(_03788_));
 sky130_as_sc_hs__or2_2 _34517_ (.A(_03731_),
    .B(_03733_),
    .Y(_03789_));
 sky130_as_sc_hs__and2_2 _34518_ (.A(_03734_),
    .B(_03789_),
    .Y(_03790_));
 sky130_as_sc_hs__and2_2 _34519_ (.A(net112),
    .B(net87),
    .Y(_03791_));
 sky130_as_sc_hs__and2_2 _34520_ (.A(net459),
    .B(net448),
    .Y(_03792_));
 sky130_as_sc_hs__and2_2 _34521_ (.A(net91),
    .B(net450),
    .Y(_03793_));
 sky130_as_sc_hs__or2_2 _34523_ (.A(_03792_),
    .B(_03793_),
    .Y(_03795_));
 sky130_as_sc_hs__and2_2 _34524_ (.A(_03794_),
    .B(_03795_),
    .Y(_03796_));
 sky130_as_sc_hs__or2_2 _34526_ (.A(_03791_),
    .B(_03796_),
    .Y(_03798_));
 sky130_as_sc_hs__and2_2 _34527_ (.A(_03797_),
    .B(_03798_),
    .Y(_03799_));
 sky130_as_sc_hs__and2_2 _34529_ (.A(net86),
    .B(_24814_),
    .Y(_03801_));
 sky130_as_sc_hs__and2_2 _34530_ (.A(net453),
    .B(_24808_),
    .Y(_03802_));
 sky130_as_sc_hs__or2_2 _34532_ (.A(_03801_),
    .B(_03802_),
    .Y(_03804_));
 sky130_as_sc_hs__and2_2 _34533_ (.A(_03803_),
    .B(_03804_),
    .Y(_03805_));
 sky130_as_sc_hs__and2_2 _34534_ (.A(_24501_),
    .B(_24774_),
    .Y(_03806_));
 sky130_as_sc_hs__and2_2 _34535_ (.A(net454),
    .B(_24768_),
    .Y(_03807_));
 sky130_as_sc_hs__or2_2 _34537_ (.A(_03806_),
    .B(_03807_),
    .Y(_03809_));
 sky130_as_sc_hs__or2_2 _34539_ (.A(_03703_),
    .B(_03810_),
    .Y(_03811_));
 sky130_as_sc_hs__and2_2 _34541_ (.A(_03811_),
    .B(_03812_),
    .Y(_03813_));
 sky130_as_sc_hs__or2_2 _34543_ (.A(_03805_),
    .B(_03813_),
    .Y(_03815_));
 sky130_as_sc_hs__and2_2 _34544_ (.A(_03814_),
    .B(_03815_),
    .Y(_03816_));
 sky130_as_sc_hs__and2_2 _34545_ (.A(_23712_),
    .B(net445),
    .Y(_03817_));
 sky130_as_sc_hs__and2_2 _34546_ (.A(_24229_),
    .B(_24729_),
    .Y(_03818_));
 sky130_as_sc_hs__or2_2 _34548_ (.A(_03817_),
    .B(_03818_),
    .Y(_03820_));
 sky130_as_sc_hs__or2_2 _34550_ (.A(_03794_),
    .B(_03821_),
    .Y(_03822_));
 sky130_as_sc_hs__or2_2 _34553_ (.A(_03718_),
    .B(_03824_),
    .Y(_03825_));
 sky130_as_sc_hs__and2_2 _34555_ (.A(_03825_),
    .B(_03826_),
    .Y(_03827_));
 sky130_as_sc_hs__or2_2 _34559_ (.A(_03827_),
    .B(_03829_),
    .Y(_03831_));
 sky130_as_sc_hs__and2_2 _34560_ (.A(_03830_),
    .B(_03831_),
    .Y(_03832_));
 sky130_as_sc_hs__or2_2 _34562_ (.A(_03816_),
    .B(_03832_),
    .Y(_03834_));
 sky130_as_sc_hs__and2_2 _34563_ (.A(_03833_),
    .B(_03834_),
    .Y(_03835_));
 sky130_as_sc_hs__or2_2 _34567_ (.A(_03835_),
    .B(_03837_),
    .Y(_03839_));
 sky130_as_sc_hs__and2_2 _34568_ (.A(_03838_),
    .B(_03839_),
    .Y(_03840_));
 sky130_as_sc_hs__and2_2 _34569_ (.A(net90),
    .B(net448),
    .Y(_03841_));
 sky130_as_sc_hs__and2_2 _34570_ (.A(_24053_),
    .B(net450),
    .Y(_03842_));
 sky130_as_sc_hs__or2_2 _34572_ (.A(_03841_),
    .B(_03842_),
    .Y(_03844_));
 sky130_as_sc_hs__and2_2 _34573_ (.A(_03843_),
    .B(_03844_),
    .Y(_03845_));
 sky130_as_sc_hs__and2_2 _34574_ (.A(net113),
    .B(_24537_),
    .Y(_03846_));
 sky130_as_sc_hs__and2_2 _34575_ (.A(net458),
    .B(net87),
    .Y(_03847_));
 sky130_as_sc_hs__or2_2 _34577_ (.A(_03846_),
    .B(_03847_),
    .Y(_03849_));
 sky130_as_sc_hs__and2_2 _34578_ (.A(_03848_),
    .B(_03849_),
    .Y(_03850_));
 sky130_as_sc_hs__or2_2 _34580_ (.A(_03845_),
    .B(_03850_),
    .Y(_03852_));
 sky130_as_sc_hs__or2_2 _34582_ (.A(_03797_),
    .B(_03853_),
    .Y(_03854_));
 sky130_as_sc_hs__and2_2 _34584_ (.A(_03854_),
    .B(_03855_),
    .Y(_03856_));
 sky130_as_sc_hs__or2_2 _34586_ (.A(_03840_),
    .B(_03856_),
    .Y(_03858_));
 sky130_as_sc_hs__or2_2 _34588_ (.A(_03800_),
    .B(_03859_),
    .Y(_03860_));
 sky130_as_sc_hs__and2_2 _34590_ (.A(_03860_),
    .B(_03861_),
    .Y(_03862_));
 sky130_as_sc_hs__or2_2 _34592_ (.A(_03788_),
    .B(_03862_),
    .Y(_03864_));
 sky130_as_sc_hs__and2_2 _34593_ (.A(_03863_),
    .B(_03864_),
    .Y(_03865_));
 sky130_as_sc_hs__and2_2 _34595_ (.A(_03570_),
    .B(_03866_),
    .Y(_03867_));
 sky130_as_sc_hs__or2_2 _34596_ (.A(_03712_),
    .B(_03713_),
    .Y(_03868_));
 sky130_as_sc_hs__and2_2 _34597_ (.A(_03714_),
    .B(_03868_),
    .Y(_03869_));
 sky130_as_sc_hs__or2_2 _34599_ (.A(_03790_),
    .B(_03799_),
    .Y(_03871_));
 sky130_as_sc_hs__or2_2 _34601_ (.A(_03870_),
    .B(_03872_),
    .Y(_03873_));
 sky130_as_sc_hs__and2_2 _34603_ (.A(_03873_),
    .B(_03874_),
    .Y(_03875_));
 sky130_as_sc_hs__or2_2 _34604_ (.A(_03633_),
    .B(_03693_),
    .Y(_03876_));
 sky130_as_sc_hs__and2_2 _34605_ (.A(_03694_),
    .B(_03876_),
    .Y(_03877_));
 sky130_as_sc_hs__or2_2 _34609_ (.A(_03865_),
    .B(_03879_),
    .Y(_03881_));
 sky130_as_sc_hs__and2_2 _34610_ (.A(_03880_),
    .B(_03881_),
    .Y(_03882_));
 sky130_as_sc_hs__or2_2 _34612_ (.A(_03695_),
    .B(_03882_),
    .Y(_03884_));
 sky130_as_sc_hs__and2_2 _34613_ (.A(_03883_),
    .B(_03884_),
    .Y(_03885_));
 sky130_as_sc_hs__or2_2 _34614_ (.A(_03875_),
    .B(_03877_),
    .Y(_03886_));
 sky130_as_sc_hs__and2_2 _34615_ (.A(_03878_),
    .B(_03886_),
    .Y(_03887_));
 sky130_as_sc_hs__or2_2 _34616_ (.A(_03867_),
    .B(_03869_),
    .Y(_03888_));
 sky130_as_sc_hs__and2_2 _34618_ (.A(net112),
    .B(net451),
    .Y(_03890_));
 sky130_as_sc_hs__or2_2 _34619_ (.A(_03643_),
    .B(_03645_),
    .Y(_03891_));
 sky130_as_sc_hs__and2_2 _34620_ (.A(_03646_),
    .B(_03891_),
    .Y(_03892_));
 sky130_as_sc_hs__or2_2 _34621_ (.A(_03538_),
    .B(_03539_),
    .Y(_03893_));
 sky130_as_sc_hs__and2_2 _34622_ (.A(_03540_),
    .B(_03893_),
    .Y(_03894_));
 sky130_as_sc_hs__or2_2 _34624_ (.A(_03566_),
    .B(_03568_),
    .Y(_03896_));
 sky130_as_sc_hs__or2_2 _34626_ (.A(_03895_),
    .B(_03897_),
    .Y(_03898_));
 sky130_as_sc_hs__and2_2 _34628_ (.A(_03898_),
    .B(_03899_),
    .Y(_03900_));
 sky130_as_sc_hs__or2_2 _34630_ (.A(_03889_),
    .B(_03901_),
    .Y(_03902_));
 sky130_as_sc_hs__and2_2 _34632_ (.A(_03902_),
    .B(_03903_),
    .Y(_03904_));
 sky130_as_sc_hs__or2_2 _34633_ (.A(_03670_),
    .B(_03691_),
    .Y(_03905_));
 sky130_as_sc_hs__or2_2 _34635_ (.A(_03898_),
    .B(_03906_),
    .Y(_03907_));
 sky130_as_sc_hs__and2_2 _34637_ (.A(_03907_),
    .B(_03908_),
    .Y(_03909_));
 sky130_as_sc_hs__or2_2 _34638_ (.A(_03663_),
    .B(_03665_),
    .Y(_03910_));
 sky130_as_sc_hs__and2_2 _34639_ (.A(_03666_),
    .B(_03910_),
    .Y(_03911_));
 sky130_as_sc_hs__or2_2 _34640_ (.A(_03636_),
    .B(_03637_),
    .Y(_03912_));
 sky130_as_sc_hs__and2_2 _34642_ (.A(net91),
    .B(_24774_),
    .Y(_03914_));
 sky130_as_sc_hs__and2_2 _34643_ (.A(_23712_),
    .B(_24768_),
    .Y(_03915_));
 sky130_as_sc_hs__or2_2 _34645_ (.A(_03913_),
    .B(_03916_),
    .Y(_03917_));
 sky130_as_sc_hs__or2_2 _34646_ (.A(_03651_),
    .B(_03652_),
    .Y(_03918_));
 sky130_as_sc_hs__and2_2 _34647_ (.A(_03653_),
    .B(_03918_),
    .Y(_03919_));
 sky130_as_sc_hs__and2_2 _34649_ (.A(_03917_),
    .B(_03920_),
    .Y(_03921_));
 sky130_as_sc_hs__and2_2 _34653_ (.A(_03662_),
    .B(_03924_),
    .Y(_03925_));
 sky130_as_sc_hs__or2_2 _34655_ (.A(_03659_),
    .B(_03660_),
    .Y(_03927_));
 sky130_as_sc_hs__and2_2 _34657_ (.A(_24216_),
    .B(_24814_),
    .Y(_03929_));
 sky130_as_sc_hs__and2_2 _34658_ (.A(_24229_),
    .B(_24808_),
    .Y(_03930_));
 sky130_as_sc_hs__or2_2 _34660_ (.A(_03928_),
    .B(_03931_),
    .Y(_03932_));
 sky130_as_sc_hs__and2_2 _34663_ (.A(_24501_),
    .B(_25205_),
    .Y(_03935_));
 sky130_as_sc_hs__and2_2 _34664_ (.A(_24256_),
    .B(_25211_),
    .Y(_03936_));
 sky130_as_sc_hs__or2_2 _34666_ (.A(_03934_),
    .B(_03937_),
    .Y(_03938_));
 sky130_as_sc_hs__or2_2 _34668_ (.A(_03923_),
    .B(_03925_),
    .Y(_03940_));
 sky130_as_sc_hs__and2_2 _34669_ (.A(_03926_),
    .B(_03940_),
    .Y(_03941_));
 sky130_as_sc_hs__or2_2 _34673_ (.A(_03911_),
    .B(_03943_),
    .Y(_03945_));
 sky130_as_sc_hs__and2_2 _34674_ (.A(_03944_),
    .B(_03945_),
    .Y(_03946_));
 sky130_as_sc_hs__inv_2 _34676_ (.Y(_03948_),
    .A(_03947_));
 sky130_as_sc_hs__or2_2 _34677_ (.A(_03681_),
    .B(_03683_),
    .Y(_03949_));
 sky130_as_sc_hs__and2_2 _34678_ (.A(_03684_),
    .B(_03949_),
    .Y(_03950_));
 sky130_as_sc_hs__or2_2 _34679_ (.A(_03677_),
    .B(_03678_),
    .Y(_03951_));
 sky130_as_sc_hs__and2_2 _34681_ (.A(_23636_),
    .B(_23712_),
    .Y(_03953_));
 sky130_as_sc_hs__and2_2 _34682_ (.A(net112),
    .B(net483),
    .Y(_03954_));
 sky130_as_sc_hs__or2_2 _34684_ (.A(_03952_),
    .B(_03955_),
    .Y(_03956_));
 sky130_as_sc_hs__and2_2 _34685_ (.A(net114),
    .B(net85),
    .Y(_03957_));
 sky130_as_sc_hs__and2_2 _34687_ (.A(_03956_),
    .B(_03958_),
    .Y(_03959_));
 sky130_as_sc_hs__or2_2 _34691_ (.A(_03950_),
    .B(_03961_),
    .Y(_03963_));
 sky130_as_sc_hs__and2_2 _34692_ (.A(_03962_),
    .B(_03963_),
    .Y(_03964_));
 sky130_as_sc_hs__or2_2 _34694_ (.A(_03948_),
    .B(_03964_),
    .Y(_03966_));
 sky130_as_sc_hs__and2_2 _34695_ (.A(_03965_),
    .B(_03966_),
    .Y(_03967_));
 sky130_as_sc_hs__or2_2 _34699_ (.A(_03909_),
    .B(_03969_),
    .Y(_03971_));
 sky130_as_sc_hs__and2_2 _34700_ (.A(_03970_),
    .B(_03971_),
    .Y(_03972_));
 sky130_as_sc_hs__or2_2 _34705_ (.A(_03887_),
    .B(_03974_),
    .Y(_03977_));
 sky130_as_sc_hs__and2_2 _34706_ (.A(_03975_),
    .B(_03977_),
    .Y(_03978_));
 sky130_as_sc_hs__or2_2 _34710_ (.A(_03885_),
    .B(_03980_),
    .Y(_03982_));
 sky130_as_sc_hs__and2_2 _34711_ (.A(_03981_),
    .B(_03982_),
    .Y(_03983_));
 sky130_as_sc_hs__or2_2 _34713_ (.A(_03510_),
    .B(_03983_),
    .Y(_03985_));
 sky130_as_sc_hs__or2_2 _34715_ (.A(_03976_),
    .B(_03978_),
    .Y(_03987_));
 sky130_as_sc_hs__and2_2 _34716_ (.A(_03979_),
    .B(_03987_),
    .Y(_03988_));
 sky130_as_sc_hs__or2_2 _34717_ (.A(_03904_),
    .B(_03972_),
    .Y(_03989_));
 sky130_as_sc_hs__and2_2 _34719_ (.A(net458),
    .B(_24729_),
    .Y(_03991_));
 sky130_as_sc_hs__or2_2 _34720_ (.A(_03919_),
    .B(_03921_),
    .Y(_03992_));
 sky130_as_sc_hs__and2_2 _34721_ (.A(_03922_),
    .B(_03992_),
    .Y(_03993_));
 sky130_as_sc_hs__or2_2 _34723_ (.A(_03892_),
    .B(_03894_),
    .Y(_03995_));
 sky130_as_sc_hs__or2_2 _34725_ (.A(_03994_),
    .B(_03996_),
    .Y(_03997_));
 sky130_as_sc_hs__or2_2 _34726_ (.A(_03946_),
    .B(_03967_),
    .Y(_03998_));
 sky130_as_sc_hs__or2_2 _34728_ (.A(_03997_),
    .B(_03999_),
    .Y(_04000_));
 sky130_as_sc_hs__and2_2 _34730_ (.A(_04000_),
    .B(_04001_),
    .Y(_04002_));
 sky130_as_sc_hs__or2_2 _34731_ (.A(_03939_),
    .B(_03941_),
    .Y(_04003_));
 sky130_as_sc_hs__and2_2 _34732_ (.A(_03942_),
    .B(_04003_),
    .Y(_04004_));
 sky130_as_sc_hs__or2_2 _34733_ (.A(_03914_),
    .B(_03915_),
    .Y(_04005_));
 sky130_as_sc_hs__and2_2 _34735_ (.A(net458),
    .B(_24774_),
    .Y(_04007_));
 sky130_as_sc_hs__and2_2 _34736_ (.A(_24053_),
    .B(_24768_),
    .Y(_04008_));
 sky130_as_sc_hs__or2_2 _34738_ (.A(_04006_),
    .B(_04009_),
    .Y(_04010_));
 sky130_as_sc_hs__or2_2 _34739_ (.A(_03929_),
    .B(_03930_),
    .Y(_04011_));
 sky130_as_sc_hs__and2_2 _34740_ (.A(_03931_),
    .B(_04011_),
    .Y(_04012_));
 sky130_as_sc_hs__and2_2 _34742_ (.A(_04010_),
    .B(_04013_),
    .Y(_04014_));
 sky130_as_sc_hs__and2_2 _34746_ (.A(_03938_),
    .B(_04017_),
    .Y(_04018_));
 sky130_as_sc_hs__or2_2 _34748_ (.A(_03935_),
    .B(_03936_),
    .Y(_04020_));
 sky130_as_sc_hs__and2_2 _34750_ (.A(_23712_),
    .B(_24814_),
    .Y(_04022_));
 sky130_as_sc_hs__and2_2 _34751_ (.A(_24216_),
    .B(_24808_),
    .Y(_04023_));
 sky130_as_sc_hs__or2_2 _34753_ (.A(_04021_),
    .B(_04024_),
    .Y(_04025_));
 sky130_as_sc_hs__and2_2 _34756_ (.A(_24256_),
    .B(_25205_),
    .Y(_04028_));
 sky130_as_sc_hs__and2_2 _34757_ (.A(_24229_),
    .B(_25211_),
    .Y(_04029_));
 sky130_as_sc_hs__or2_2 _34759_ (.A(_04027_),
    .B(_04030_),
    .Y(_04031_));
 sky130_as_sc_hs__or2_2 _34761_ (.A(_04016_),
    .B(_04018_),
    .Y(_04033_));
 sky130_as_sc_hs__and2_2 _34762_ (.A(_04019_),
    .B(_04033_),
    .Y(_04034_));
 sky130_as_sc_hs__or2_2 _34766_ (.A(_04004_),
    .B(_04036_),
    .Y(_04038_));
 sky130_as_sc_hs__and2_2 _34767_ (.A(_04037_),
    .B(_04038_),
    .Y(_04039_));
 sky130_as_sc_hs__inv_2 _34769_ (.Y(_04041_),
    .A(_04040_));
 sky130_as_sc_hs__or2_2 _34770_ (.A(_03957_),
    .B(_03959_),
    .Y(_04042_));
 sky130_as_sc_hs__and2_2 _34772_ (.A(net114),
    .B(net454),
    .Y(_04044_));
 sky130_as_sc_hs__or2_2 _34773_ (.A(_03953_),
    .B(_03954_),
    .Y(_04045_));
 sky130_as_sc_hs__and2_2 _34774_ (.A(_03955_),
    .B(_04045_),
    .Y(_04046_));
 sky130_as_sc_hs__or2_2 _34776_ (.A(_04043_),
    .B(_04047_),
    .Y(_04048_));
 sky130_as_sc_hs__and2_2 _34778_ (.A(_04048_),
    .B(_04049_),
    .Y(_04050_));
 sky130_as_sc_hs__or2_2 _34780_ (.A(_04041_),
    .B(_04050_),
    .Y(_04052_));
 sky130_as_sc_hs__and2_2 _34781_ (.A(_04051_),
    .B(_04052_),
    .Y(_04053_));
 sky130_as_sc_hs__or2_2 _34785_ (.A(_04002_),
    .B(_04055_),
    .Y(_04057_));
 sky130_as_sc_hs__and2_2 _34786_ (.A(_04056_),
    .B(_04057_),
    .Y(_04058_));
 sky130_as_sc_hs__or2_2 _34787_ (.A(_03890_),
    .B(_03900_),
    .Y(_04059_));
 sky130_as_sc_hs__and2_2 _34788_ (.A(_03901_),
    .B(_04059_),
    .Y(_04060_));
 sky130_as_sc_hs__or2_2 _34790_ (.A(_03990_),
    .B(_04061_),
    .Y(_04062_));
 sky130_as_sc_hs__and2_2 _34793_ (.A(_04062_),
    .B(_04064_),
    .Y(_04065_));
 sky130_as_sc_hs__or2_2 _34798_ (.A(_03988_),
    .B(_04067_),
    .Y(_04070_));
 sky130_as_sc_hs__and2_2 _34799_ (.A(_04068_),
    .B(_04070_),
    .Y(_04071_));
 sky130_as_sc_hs__and2_2 _34801_ (.A(_04068_),
    .B(_04072_),
    .Y(_04073_));
 sky130_as_sc_hs__or2_2 _34803_ (.A(_03986_),
    .B(_04073_),
    .Y(_04075_));
 sky130_as_sc_hs__or2_2 _34804_ (.A(_04069_),
    .B(_04071_),
    .Y(_04076_));
 sky130_as_sc_hs__and2_2 _34805_ (.A(_04072_),
    .B(_04076_),
    .Y(_04077_));
 sky130_as_sc_hs__or2_2 _34806_ (.A(_04063_),
    .B(_04065_),
    .Y(_04078_));
 sky130_as_sc_hs__and2_2 _34807_ (.A(_04066_),
    .B(_04078_),
    .Y(_04079_));
 sky130_as_sc_hs__or2_2 _34808_ (.A(_04058_),
    .B(_04060_),
    .Y(_04080_));
 sky130_as_sc_hs__and2_2 _34810_ (.A(net112),
    .B(_24729_),
    .Y(_04082_));
 sky130_as_sc_hs__or2_2 _34811_ (.A(_04012_),
    .B(_04014_),
    .Y(_04083_));
 sky130_as_sc_hs__and2_2 _34812_ (.A(_04015_),
    .B(_04083_),
    .Y(_04084_));
 sky130_as_sc_hs__or2_2 _34814_ (.A(_03991_),
    .B(_03993_),
    .Y(_04086_));
 sky130_as_sc_hs__or2_2 _34816_ (.A(_04085_),
    .B(_04087_),
    .Y(_04088_));
 sky130_as_sc_hs__or2_2 _34817_ (.A(_04039_),
    .B(_04053_),
    .Y(_04089_));
 sky130_as_sc_hs__or2_2 _34819_ (.A(_04088_),
    .B(_04090_),
    .Y(_04091_));
 sky130_as_sc_hs__and2_2 _34821_ (.A(_04091_),
    .B(_04092_),
    .Y(_04093_));
 sky130_as_sc_hs__or2_2 _34822_ (.A(_04032_),
    .B(_04034_),
    .Y(_04094_));
 sky130_as_sc_hs__and2_2 _34823_ (.A(_04035_),
    .B(_04094_),
    .Y(_04095_));
 sky130_as_sc_hs__or2_2 _34824_ (.A(_04007_),
    .B(_04008_),
    .Y(_04096_));
 sky130_as_sc_hs__and2_2 _34826_ (.A(net91),
    .B(_24768_),
    .Y(_04098_));
 sky130_as_sc_hs__and2_2 _34827_ (.A(net113),
    .B(_24774_),
    .Y(_04099_));
 sky130_as_sc_hs__or2_2 _34829_ (.A(_04097_),
    .B(_04100_),
    .Y(_04101_));
 sky130_as_sc_hs__and2_2 _34831_ (.A(_04101_),
    .B(_04102_),
    .Y(_04103_));
 sky130_as_sc_hs__or2_2 _34832_ (.A(_04022_),
    .B(_04023_),
    .Y(_04104_));
 sky130_as_sc_hs__and2_2 _34833_ (.A(_04024_),
    .B(_04104_),
    .Y(_04105_));
 sky130_as_sc_hs__and2_2 _34837_ (.A(_04031_),
    .B(_04108_),
    .Y(_04109_));
 sky130_as_sc_hs__or2_2 _34839_ (.A(_04028_),
    .B(_04029_),
    .Y(_04111_));
 sky130_as_sc_hs__and2_2 _34841_ (.A(_24053_),
    .B(_24814_),
    .Y(_04113_));
 sky130_as_sc_hs__and2_2 _34842_ (.A(_23712_),
    .B(_24808_),
    .Y(_04114_));
 sky130_as_sc_hs__or2_2 _34844_ (.A(_04112_),
    .B(_04115_),
    .Y(_04116_));
 sky130_as_sc_hs__and2_2 _34847_ (.A(_24229_),
    .B(_25205_),
    .Y(_04119_));
 sky130_as_sc_hs__and2_2 _34848_ (.A(_24216_),
    .B(_25211_),
    .Y(_04120_));
 sky130_as_sc_hs__or2_2 _34850_ (.A(_04118_),
    .B(_04121_),
    .Y(_04122_));
 sky130_as_sc_hs__or2_2 _34852_ (.A(_04107_),
    .B(_04109_),
    .Y(_04124_));
 sky130_as_sc_hs__and2_2 _34853_ (.A(_04110_),
    .B(_04124_),
    .Y(_04125_));
 sky130_as_sc_hs__or2_2 _34857_ (.A(_04044_),
    .B(_04046_),
    .Y(_04129_));
 sky130_as_sc_hs__and2_2 _34859_ (.A(_23636_),
    .B(_24053_),
    .Y(_04131_));
 sky130_as_sc_hs__and2_2 _34860_ (.A(net114),
    .B(_24545_),
    .Y(_04132_));
 sky130_as_sc_hs__or2_2 _34862_ (.A(_04130_),
    .B(_04133_),
    .Y(_04134_));
 sky130_as_sc_hs__and2_2 _34864_ (.A(_04134_),
    .B(_04135_),
    .Y(_04136_));
 sky130_as_sc_hs__inv_2 _34866_ (.Y(_04138_),
    .A(_04137_));
 sky130_as_sc_hs__or2_2 _34868_ (.A(_04136_),
    .B(_04138_),
    .Y(_04140_));
 sky130_as_sc_hs__and2_2 _34869_ (.A(_04139_),
    .B(_04140_),
    .Y(_04141_));
 sky130_as_sc_hs__or2_2 _34870_ (.A(_04095_),
    .B(_04127_),
    .Y(_04142_));
 sky130_as_sc_hs__and2_2 _34871_ (.A(_04128_),
    .B(_04142_),
    .Y(_04143_));
 sky130_as_sc_hs__or2_2 _34875_ (.A(_04093_),
    .B(_04145_),
    .Y(_04147_));
 sky130_as_sc_hs__and2_2 _34876_ (.A(_04146_),
    .B(_04147_),
    .Y(_04148_));
 sky130_as_sc_hs__and2_2 _34878_ (.A(_03997_),
    .B(_04149_),
    .Y(_04150_));
 sky130_as_sc_hs__or2_2 _34880_ (.A(_04081_),
    .B(_04151_),
    .Y(_04152_));
 sky130_as_sc_hs__and2_2 _34883_ (.A(_04152_),
    .B(_04154_),
    .Y(_04155_));
 sky130_as_sc_hs__or2_2 _34888_ (.A(_04079_),
    .B(_04157_),
    .Y(_04160_));
 sky130_as_sc_hs__and2_2 _34889_ (.A(_04158_),
    .B(_04160_),
    .Y(_04161_));
 sky130_as_sc_hs__or2_2 _34893_ (.A(_04159_),
    .B(_04161_),
    .Y(_04165_));
 sky130_as_sc_hs__and2_2 _34894_ (.A(_04162_),
    .B(_04165_),
    .Y(_04166_));
 sky130_as_sc_hs__or2_2 _34895_ (.A(_04153_),
    .B(_04155_),
    .Y(_04167_));
 sky130_as_sc_hs__or2_2 _34897_ (.A(_04148_),
    .B(_04150_),
    .Y(_04169_));
 sky130_as_sc_hs__and2_2 _34898_ (.A(_04151_),
    .B(_04169_),
    .Y(_04170_));
 sky130_as_sc_hs__or2_2 _34899_ (.A(_04141_),
    .B(_04143_),
    .Y(_04171_));
 sky130_as_sc_hs__and2_2 _34900_ (.A(_04144_),
    .B(_04171_),
    .Y(_04172_));
 sky130_as_sc_hs__or2_2 _34901_ (.A(_04123_),
    .B(_04125_),
    .Y(_04173_));
 sky130_as_sc_hs__and2_2 _34902_ (.A(_04126_),
    .B(_04173_),
    .Y(_04174_));
 sky130_as_sc_hs__or2_2 _34903_ (.A(_04113_),
    .B(_04114_),
    .Y(_04175_));
 sky130_as_sc_hs__and2_2 _34904_ (.A(_04115_),
    .B(_04175_),
    .Y(_04176_));
 sky130_as_sc_hs__or2_2 _34905_ (.A(_04098_),
    .B(_04099_),
    .Y(_04177_));
 sky130_as_sc_hs__and2_2 _34906_ (.A(_04100_),
    .B(_04177_),
    .Y(_04178_));
 sky130_as_sc_hs__or2_2 _34910_ (.A(_04179_),
    .B(_04181_),
    .Y(_04182_));
 sky130_as_sc_hs__or2_2 _34911_ (.A(_04119_),
    .B(_04120_),
    .Y(_04183_));
 sky130_as_sc_hs__and2_2 _34913_ (.A(net91),
    .B(_24814_),
    .Y(_04185_));
 sky130_as_sc_hs__and2_2 _34914_ (.A(_24053_),
    .B(_24808_),
    .Y(_04186_));
 sky130_as_sc_hs__or2_2 _34916_ (.A(_04184_),
    .B(_04187_),
    .Y(_04188_));
 sky130_as_sc_hs__and2_2 _34919_ (.A(_24216_),
    .B(_25205_),
    .Y(_04191_));
 sky130_as_sc_hs__and2_2 _34920_ (.A(_23712_),
    .B(_25211_),
    .Y(_04192_));
 sky130_as_sc_hs__or2_2 _34922_ (.A(_04190_),
    .B(_04193_),
    .Y(_04194_));
 sky130_as_sc_hs__and2_2 _34925_ (.A(_04182_),
    .B(_04196_),
    .Y(_04197_));
 sky130_as_sc_hs__or2_2 _34929_ (.A(_04131_),
    .B(_04132_),
    .Y(_04201_));
 sky130_as_sc_hs__and2_2 _34931_ (.A(_23636_),
    .B(net91),
    .Y(_04203_));
 sky130_as_sc_hs__and2_2 _34932_ (.A(net114),
    .B(_24501_),
    .Y(_04204_));
 sky130_as_sc_hs__or2_2 _34934_ (.A(_04202_),
    .B(_04205_),
    .Y(_04206_));
 sky130_as_sc_hs__and2_2 _34936_ (.A(_04206_),
    .B(_04207_),
    .Y(_04208_));
 sky130_as_sc_hs__inv_2 _34938_ (.Y(_04210_),
    .A(_04209_));
 sky130_as_sc_hs__or2_2 _34940_ (.A(_04208_),
    .B(_04210_),
    .Y(_04212_));
 sky130_as_sc_hs__and2_2 _34941_ (.A(_04211_),
    .B(_04212_),
    .Y(_04213_));
 sky130_as_sc_hs__or2_2 _34942_ (.A(_04174_),
    .B(_04199_),
    .Y(_04214_));
 sky130_as_sc_hs__and2_2 _34943_ (.A(_04200_),
    .B(_04214_),
    .Y(_04215_));
 sky130_as_sc_hs__or2_2 _34947_ (.A(_04172_),
    .B(_04217_),
    .Y(_04219_));
 sky130_as_sc_hs__and2_2 _34948_ (.A(_04218_),
    .B(_04219_),
    .Y(_04220_));
 sky130_as_sc_hs__and2_2 _34950_ (.A(_04088_),
    .B(_04221_),
    .Y(_04222_));
 sky130_as_sc_hs__or2_2 _34954_ (.A(_04168_),
    .B(_04225_),
    .Y(_04226_));
 sky130_as_sc_hs__and2_2 _34957_ (.A(_04226_),
    .B(_04228_),
    .Y(_04229_));
 sky130_as_sc_hs__or2_2 _34961_ (.A(_04227_),
    .B(_04229_),
    .Y(_04233_));
 sky130_as_sc_hs__and2_2 _34962_ (.A(_04230_),
    .B(_04233_),
    .Y(_04234_));
 sky130_as_sc_hs__or2_2 _34963_ (.A(_04170_),
    .B(_04224_),
    .Y(_04235_));
 sky130_as_sc_hs__or2_2 _34965_ (.A(_04220_),
    .B(_04222_),
    .Y(_04237_));
 sky130_as_sc_hs__and2_2 _34966_ (.A(_04223_),
    .B(_04237_),
    .Y(_04238_));
 sky130_as_sc_hs__or2_2 _34967_ (.A(_04213_),
    .B(_04215_),
    .Y(_04239_));
 sky130_as_sc_hs__and2_2 _34968_ (.A(_04216_),
    .B(_04239_),
    .Y(_04240_));
 sky130_as_sc_hs__or2_2 _34969_ (.A(_04195_),
    .B(_04197_),
    .Y(_04241_));
 sky130_as_sc_hs__and2_2 _34970_ (.A(_04198_),
    .B(_04241_),
    .Y(_04242_));
 sky130_as_sc_hs__and2_2 _34971_ (.A(net459),
    .B(_24768_),
    .Y(_04243_));
 sky130_as_sc_hs__or2_2 _34972_ (.A(_04185_),
    .B(_04186_),
    .Y(_04244_));
 sky130_as_sc_hs__and2_2 _34973_ (.A(_04187_),
    .B(_04244_),
    .Y(_04245_));
 sky130_as_sc_hs__or2_2 _34977_ (.A(_04246_),
    .B(_04248_),
    .Y(_04249_));
 sky130_as_sc_hs__or2_2 _34978_ (.A(_04191_),
    .B(_04192_),
    .Y(_04250_));
 sky130_as_sc_hs__and2_2 _34980_ (.A(net91),
    .B(_24808_),
    .Y(_04252_));
 sky130_as_sc_hs__and2_2 _34981_ (.A(net459),
    .B(_24814_),
    .Y(_04253_));
 sky130_as_sc_hs__or2_2 _34983_ (.A(_04251_),
    .B(_04254_),
    .Y(_04255_));
 sky130_as_sc_hs__and2_2 _34986_ (.A(_23712_),
    .B(_25205_),
    .Y(_04258_));
 sky130_as_sc_hs__and2_2 _34987_ (.A(_24053_),
    .B(_25211_),
    .Y(_04259_));
 sky130_as_sc_hs__or2_2 _34989_ (.A(_04257_),
    .B(_04260_),
    .Y(_04261_));
 sky130_as_sc_hs__and2_2 _34992_ (.A(_04249_),
    .B(_04263_),
    .Y(_04264_));
 sky130_as_sc_hs__or2_2 _34996_ (.A(_04203_),
    .B(_04204_),
    .Y(_04268_));
 sky130_as_sc_hs__and2_2 _34998_ (.A(_23636_),
    .B(net459),
    .Y(_04270_));
 sky130_as_sc_hs__and2_2 _34999_ (.A(net114),
    .B(_24256_),
    .Y(_04271_));
 sky130_as_sc_hs__or2_2 _35001_ (.A(_04269_),
    .B(_04272_),
    .Y(_04273_));
 sky130_as_sc_hs__and2_2 _35003_ (.A(_04273_),
    .B(_04274_),
    .Y(_04275_));
 sky130_as_sc_hs__inv_2 _35005_ (.Y(_04277_),
    .A(_04276_));
 sky130_as_sc_hs__or2_2 _35007_ (.A(_04275_),
    .B(_04277_),
    .Y(_04279_));
 sky130_as_sc_hs__and2_2 _35008_ (.A(_04278_),
    .B(_04279_),
    .Y(_04280_));
 sky130_as_sc_hs__or2_2 _35009_ (.A(_04242_),
    .B(_04266_),
    .Y(_04281_));
 sky130_as_sc_hs__and2_2 _35010_ (.A(_04267_),
    .B(_04281_),
    .Y(_04282_));
 sky130_as_sc_hs__or2_2 _35014_ (.A(_04240_),
    .B(_04284_),
    .Y(_04286_));
 sky130_as_sc_hs__and2_2 _35015_ (.A(_04285_),
    .B(_04286_),
    .Y(_04287_));
 sky130_as_sc_hs__or2_2 _35016_ (.A(_04082_),
    .B(_04084_),
    .Y(_04288_));
 sky130_as_sc_hs__and2_2 _35017_ (.A(_04085_),
    .B(_04288_),
    .Y(_04289_));
 sky130_as_sc_hs__or2_2 _35021_ (.A(_04236_),
    .B(_04292_),
    .Y(_04293_));
 sky130_as_sc_hs__and2_2 _35024_ (.A(_04293_),
    .B(_04295_),
    .Y(_04296_));
 sky130_as_sc_hs__or2_2 _35028_ (.A(_04234_),
    .B(_04298_),
    .Y(_04300_));
 sky130_as_sc_hs__and2_2 _35029_ (.A(_04299_),
    .B(_04300_),
    .Y(_04301_));
 sky130_as_sc_hs__or2_2 _35030_ (.A(_04294_),
    .B(_04296_),
    .Y(_04302_));
 sky130_as_sc_hs__and2_2 _35031_ (.A(_04297_),
    .B(_04302_),
    .Y(_04303_));
 sky130_as_sc_hs__or2_2 _35032_ (.A(_04287_),
    .B(_04289_),
    .Y(_04304_));
 sky130_as_sc_hs__and2_2 _35033_ (.A(_04290_),
    .B(_04304_),
    .Y(_04305_));
 sky130_as_sc_hs__or2_2 _35034_ (.A(_04280_),
    .B(_04282_),
    .Y(_04306_));
 sky130_as_sc_hs__and2_2 _35035_ (.A(_04283_),
    .B(_04306_),
    .Y(_04307_));
 sky130_as_sc_hs__or2_2 _35036_ (.A(_04262_),
    .B(_04264_),
    .Y(_04308_));
 sky130_as_sc_hs__and2_2 _35037_ (.A(_04265_),
    .B(_04308_),
    .Y(_04309_));
 sky130_as_sc_hs__and2_2 _35038_ (.A(net113),
    .B(_24768_),
    .Y(_04310_));
 sky130_as_sc_hs__or2_2 _35039_ (.A(_04252_),
    .B(_04253_),
    .Y(_04311_));
 sky130_as_sc_hs__and2_2 _35040_ (.A(_04254_),
    .B(_04311_),
    .Y(_04312_));
 sky130_as_sc_hs__or2_2 _35044_ (.A(_04313_),
    .B(_04315_),
    .Y(_04316_));
 sky130_as_sc_hs__and2_2 _35046_ (.A(_04316_),
    .B(_04317_),
    .Y(_04318_));
 sky130_as_sc_hs__or2_2 _35047_ (.A(_04258_),
    .B(_04259_),
    .Y(_04319_));
 sky130_as_sc_hs__and2_2 _35049_ (.A(net459),
    .B(_24808_),
    .Y(_04321_));
 sky130_as_sc_hs__and2_2 _35050_ (.A(net113),
    .B(_24814_),
    .Y(_04322_));
 sky130_as_sc_hs__or2_2 _35052_ (.A(_04320_),
    .B(_04323_),
    .Y(_04324_));
 sky130_as_sc_hs__and2_2 _35054_ (.A(net91),
    .B(_25211_),
    .Y(_04326_));
 sky130_as_sc_hs__and2_2 _35055_ (.A(_24053_),
    .B(_25205_),
    .Y(_04327_));
 sky130_as_sc_hs__inv_2 _35057_ (.Y(_04329_),
    .A(_04328_));
 sky130_as_sc_hs__or2_2 _35063_ (.A(_04270_),
    .B(_04271_),
    .Y(_04335_));
 sky130_as_sc_hs__and2_2 _35065_ (.A(net112),
    .B(_23636_),
    .Y(_04337_));
 sky130_as_sc_hs__and2_2 _35066_ (.A(net114),
    .B(_24229_),
    .Y(_04338_));
 sky130_as_sc_hs__or2_2 _35068_ (.A(_04336_),
    .B(_04339_),
    .Y(_04340_));
 sky130_as_sc_hs__and2_2 _35070_ (.A(_04340_),
    .B(_04341_),
    .Y(_04342_));
 sky130_as_sc_hs__or2_2 _35071_ (.A(_04309_),
    .B(_04333_),
    .Y(_04343_));
 sky130_as_sc_hs__and2_2 _35072_ (.A(_04334_),
    .B(_04343_),
    .Y(_04344_));
 sky130_as_sc_hs__or2_2 _35076_ (.A(_04307_),
    .B(_04346_),
    .Y(_04348_));
 sky130_as_sc_hs__and2_2 _35077_ (.A(_04347_),
    .B(_04348_),
    .Y(_04349_));
 sky130_as_sc_hs__or2_2 _35078_ (.A(_04103_),
    .B(_04105_),
    .Y(_04350_));
 sky130_as_sc_hs__and2_2 _35079_ (.A(_04106_),
    .B(_04350_),
    .Y(_04351_));
 sky130_as_sc_hs__or2_2 _35083_ (.A(_04238_),
    .B(_04291_),
    .Y(_04355_));
 sky130_as_sc_hs__or2_2 _35085_ (.A(_04354_),
    .B(_04356_),
    .Y(_04357_));
 sky130_as_sc_hs__and2_2 _35088_ (.A(_04357_),
    .B(_04359_),
    .Y(_04360_));
 sky130_as_sc_hs__or2_2 _35092_ (.A(_04358_),
    .B(_04360_),
    .Y(_04364_));
 sky130_as_sc_hs__and2_2 _35093_ (.A(_04361_),
    .B(_04364_),
    .Y(_04365_));
 sky130_as_sc_hs__or2_2 _35094_ (.A(_04305_),
    .B(_04353_),
    .Y(_04366_));
 sky130_as_sc_hs__or2_2 _35096_ (.A(_04349_),
    .B(_04351_),
    .Y(_04368_));
 sky130_as_sc_hs__and2_2 _35097_ (.A(_04352_),
    .B(_04368_),
    .Y(_04369_));
 sky130_as_sc_hs__or2_2 _35098_ (.A(_04342_),
    .B(_04344_),
    .Y(_04370_));
 sky130_as_sc_hs__and2_2 _35099_ (.A(_04345_),
    .B(_04370_),
    .Y(_04371_));
 sky130_as_sc_hs__or2_2 _35100_ (.A(_04318_),
    .B(_04331_),
    .Y(_04372_));
 sky130_as_sc_hs__and2_2 _35101_ (.A(_04332_),
    .B(_04372_),
    .Y(_04373_));
 sky130_as_sc_hs__and2_2 _35102_ (.A(_04324_),
    .B(_04325_),
    .Y(_04374_));
 sky130_as_sc_hs__and2_2 _35103_ (.A(net459),
    .B(_25211_),
    .Y(_04375_));
 sky130_as_sc_hs__and2_2 _35104_ (.A(net91),
    .B(_25205_),
    .Y(_04376_));
 sky130_as_sc_hs__and2_2 _35105_ (.A(_04375_),
    .B(_04376_),
    .Y(_04377_));
 sky130_as_sc_hs__and2_2 _35106_ (.A(_04328_),
    .B(_04377_),
    .Y(_04378_));
 sky130_as_sc_hs__and2_2 _35107_ (.A(_04374_),
    .B(_04378_),
    .Y(_04379_));
 sky130_as_sc_hs__or2_2 _35109_ (.A(_04337_),
    .B(_04338_),
    .Y(_04381_));
 sky130_as_sc_hs__and2_2 _35110_ (.A(_04339_),
    .B(_04381_),
    .Y(_04382_));
 sky130_as_sc_hs__or2_2 _35111_ (.A(_04373_),
    .B(_04379_),
    .Y(_04383_));
 sky130_as_sc_hs__and2_2 _35112_ (.A(_04380_),
    .B(_04383_),
    .Y(_04384_));
 sky130_as_sc_hs__or2_2 _35116_ (.A(_04371_),
    .B(_04386_),
    .Y(_04388_));
 sky130_as_sc_hs__and2_2 _35117_ (.A(_04387_),
    .B(_04388_),
    .Y(_04389_));
 sky130_as_sc_hs__or2_2 _35118_ (.A(_04176_),
    .B(_04178_),
    .Y(_04390_));
 sky130_as_sc_hs__and2_2 _35119_ (.A(_04179_),
    .B(_04390_),
    .Y(_04391_));
 sky130_as_sc_hs__or2_2 _35123_ (.A(_04367_),
    .B(_04394_),
    .Y(_04395_));
 sky130_as_sc_hs__and2_2 _35126_ (.A(_04395_),
    .B(_04397_),
    .Y(_04398_));
 sky130_as_sc_hs__or2_2 _35130_ (.A(_04396_),
    .B(_04398_),
    .Y(_04402_));
 sky130_as_sc_hs__and2_2 _35131_ (.A(_04399_),
    .B(_04402_),
    .Y(_04403_));
 sky130_as_sc_hs__or2_2 _35132_ (.A(_04369_),
    .B(_04393_),
    .Y(_04404_));
 sky130_as_sc_hs__or2_2 _35134_ (.A(_04389_),
    .B(_04391_),
    .Y(_04406_));
 sky130_as_sc_hs__and2_2 _35135_ (.A(_04392_),
    .B(_04406_),
    .Y(_04407_));
 sky130_as_sc_hs__or2_2 _35136_ (.A(_04382_),
    .B(_04384_),
    .Y(_04408_));
 sky130_as_sc_hs__and2_2 _35137_ (.A(_04385_),
    .B(_04408_),
    .Y(_04409_));
 sky130_as_sc_hs__and2_2 _35138_ (.A(net113),
    .B(_25211_),
    .Y(_04410_));
 sky130_as_sc_hs__and2_2 _35139_ (.A(net459),
    .B(_25205_),
    .Y(_04411_));
 sky130_as_sc_hs__or2_2 _35141_ (.A(_04377_),
    .B(_04412_),
    .Y(_04413_));
 sky130_as_sc_hs__or2_2 _35142_ (.A(_04328_),
    .B(_04377_),
    .Y(_04414_));
 sky130_as_sc_hs__nor2_2 _35143_ (.A(_04326_),
    .B(_04327_),
    .Y(_04415_));
 sky130_as_sc_hs__nor2_2 _35144_ (.A(_04378_),
    .B(_04415_),
    .Y(_04416_));
 sky130_as_sc_hs__or2_2 _35146_ (.A(_04413_),
    .B(_04417_),
    .Y(_04418_));
 sky130_as_sc_hs__or2_2 _35147_ (.A(_04329_),
    .B(_04377_),
    .Y(_04419_));
 sky130_as_sc_hs__or2_2 _35149_ (.A(_04374_),
    .B(_04419_),
    .Y(_04421_));
 sky130_as_sc_hs__or2_2 _35151_ (.A(_04418_),
    .B(_04422_),
    .Y(_04423_));
 sky130_as_sc_hs__and2_2 _35152_ (.A(net114),
    .B(_24216_),
    .Y(_04424_));
 sky130_as_sc_hs__and2_2 _35154_ (.A(_04423_),
    .B(_04425_),
    .Y(_04426_));
 sky130_as_sc_hs__or2_2 _35158_ (.A(_04409_),
    .B(_04428_),
    .Y(_04430_));
 sky130_as_sc_hs__and2_2 _35159_ (.A(_04429_),
    .B(_04430_),
    .Y(_04431_));
 sky130_as_sc_hs__or2_2 _35160_ (.A(_04243_),
    .B(_04245_),
    .Y(_04432_));
 sky130_as_sc_hs__and2_2 _35161_ (.A(_04246_),
    .B(_04432_),
    .Y(_04433_));
 sky130_as_sc_hs__or2_2 _35165_ (.A(_04405_),
    .B(_04436_),
    .Y(_04437_));
 sky130_as_sc_hs__or2_2 _35168_ (.A(_04340_),
    .B(_04439_),
    .Y(_04440_));
 sky130_as_sc_hs__or2_2 _35171_ (.A(_04403_),
    .B(_04441_),
    .Y(_04443_));
 sky130_as_sc_hs__and2_2 _35172_ (.A(_04442_),
    .B(_04443_),
    .Y(_04444_));
 sky130_as_sc_hs__and2_2 _35174_ (.A(_04440_),
    .B(_04445_),
    .Y(_04446_));
 sky130_as_sc_hs__or2_2 _35175_ (.A(_04407_),
    .B(_04435_),
    .Y(_04447_));
 sky130_as_sc_hs__or2_2 _35177_ (.A(_04431_),
    .B(_04433_),
    .Y(_04449_));
 sky130_as_sc_hs__and2_2 _35178_ (.A(_04434_),
    .B(_04449_),
    .Y(_04450_));
 sky130_as_sc_hs__or2_2 _35179_ (.A(_04424_),
    .B(_04426_),
    .Y(_04451_));
 sky130_as_sc_hs__and2_2 _35181_ (.A(net114),
    .B(_23712_),
    .Y(_04453_));
 sky130_as_sc_hs__and2_2 _35183_ (.A(_04418_),
    .B(_04454_),
    .Y(_04455_));
 sky130_as_sc_hs__or2_2 _35185_ (.A(_04452_),
    .B(_04456_),
    .Y(_04457_));
 sky130_as_sc_hs__and2_2 _35187_ (.A(_04457_),
    .B(_04458_),
    .Y(_04459_));
 sky130_as_sc_hs__or2_2 _35188_ (.A(_04310_),
    .B(_04312_),
    .Y(_04460_));
 sky130_as_sc_hs__and2_2 _35189_ (.A(_04313_),
    .B(_04460_),
    .Y(_04461_));
 sky130_as_sc_hs__nor2_2 _35193_ (.A(_04448_),
    .B(_04464_),
    .Y(_04465_));
 sky130_as_sc_hs__or2_2 _35195_ (.A(_04446_),
    .B(_04465_),
    .Y(_04467_));
 sky130_as_sc_hs__and2_2 _35196_ (.A(_04466_),
    .B(_04467_),
    .Y(_04468_));
 sky130_as_sc_hs__or2_2 _35197_ (.A(_04450_),
    .B(_04463_),
    .Y(_04469_));
 sky130_as_sc_hs__or2_2 _35199_ (.A(_04459_),
    .B(_04461_),
    .Y(_04471_));
 sky130_as_sc_hs__and2_2 _35200_ (.A(_04462_),
    .B(_04471_),
    .Y(_04472_));
 sky130_as_sc_hs__or2_2 _35201_ (.A(_04453_),
    .B(_04455_),
    .Y(_04473_));
 sky130_as_sc_hs__or2_2 _35205_ (.A(_04375_),
    .B(_04376_),
    .Y(_04477_));
 sky130_as_sc_hs__nand3_2 _35206_ (.A(_04413_),
    .B(_04476_),
    .C(_04477_),
    .Y(_04478_));
 sky130_as_sc_hs__or2_2 _35207_ (.A(_04475_),
    .B(_04478_),
    .Y(_04479_));
 sky130_as_sc_hs__or2_2 _35208_ (.A(_04474_),
    .B(_04479_),
    .Y(_04480_));
 sky130_as_sc_hs__and2_2 _35210_ (.A(_04480_),
    .B(_04481_),
    .Y(_04482_));
 sky130_as_sc_hs__or2_2 _35211_ (.A(_04321_),
    .B(_04322_),
    .Y(_04483_));
 sky130_as_sc_hs__and2_2 _35212_ (.A(_04323_),
    .B(_04483_),
    .Y(_04484_));
 sky130_as_sc_hs__or2_2 _35216_ (.A(_04470_),
    .B(_04487_),
    .Y(_04488_));
 sky130_as_sc_hs__and2_2 _35218_ (.A(_04488_),
    .B(_04489_),
    .Y(_04490_));
 sky130_as_sc_hs__or2_2 _35219_ (.A(_04472_),
    .B(_04486_),
    .Y(_04491_));
 sky130_as_sc_hs__or2_2 _35221_ (.A(_04482_),
    .B(_04484_),
    .Y(_04493_));
 sky130_as_sc_hs__and2_2 _35222_ (.A(_04485_),
    .B(_04493_),
    .Y(_04494_));
 sky130_as_sc_hs__and2_2 _35225_ (.A(net116),
    .B(net91),
    .Y(_04497_));
 sky130_as_sc_hs__or2_2 _35226_ (.A(_04410_),
    .B(_04411_),
    .Y(_04498_));
 sky130_as_sc_hs__and2_2 _35227_ (.A(_04412_),
    .B(_04498_),
    .Y(_04499_));
 sky130_as_sc_hs__or2_2 _35229_ (.A(_04496_),
    .B(_04500_),
    .Y(_04501_));
 sky130_as_sc_hs__inv_2 _35231_ (.Y(_04503_),
    .A(_04502_));
 sky130_as_sc_hs__and2_2 _35233_ (.A(_04501_),
    .B(_04504_),
    .Y(_04505_));
 sky130_as_sc_hs__nor2_2 _35237_ (.A(_04492_),
    .B(_04508_),
    .Y(_04509_));
 sky130_as_sc_hs__or2_2 _35238_ (.A(_04497_),
    .B(_04499_),
    .Y(_04510_));
 sky130_as_sc_hs__or2_2 _35242_ (.A(_04512_),
    .B(_04513_),
    .Y(_04514_));
 sky130_as_sc_hs__nor2_2 _35243_ (.A(_04511_),
    .B(_04514_),
    .Y(_04515_));
 sky130_as_sc_hs__or2_2 _35244_ (.A(_04503_),
    .B(_04505_),
    .Y(_04516_));
 sky130_as_sc_hs__and2_2 _35245_ (.A(_04506_),
    .B(_04516_),
    .Y(_04517_));
 sky130_as_sc_hs__and2_2 _35246_ (.A(_04515_),
    .B(_04517_),
    .Y(_04518_));
 sky130_as_sc_hs__or2_2 _35247_ (.A(_04494_),
    .B(_04507_),
    .Y(_04519_));
 sky130_as_sc_hs__and2_2 _35248_ (.A(_04508_),
    .B(_04519_),
    .Y(_04520_));
 sky130_as_sc_hs__and2_2 _35249_ (.A(_04518_),
    .B(_04520_),
    .Y(_04521_));
 sky130_as_sc_hs__inv_2 _35250_ (.Y(_04522_),
    .A(_04521_));
 sky130_as_sc_hs__nor2_2 _35251_ (.A(_04492_),
    .B(_04522_),
    .Y(_04523_));
 sky130_as_sc_hs__or2_2 _35252_ (.A(_04509_),
    .B(_04523_),
    .Y(_04524_));
 sky130_as_sc_hs__nand3_2 _35253_ (.A(_04488_),
    .B(_04489_),
    .C(_04524_),
    .Y(_04525_));
 sky130_as_sc_hs__inv_2 _35254_ (.Y(_04526_),
    .A(_04525_));
 sky130_as_sc_hs__and2_2 _35255_ (.A(_04464_),
    .B(_04488_),
    .Y(_04527_));
 sky130_as_sc_hs__or2_2 _35256_ (.A(_04448_),
    .B(_04527_),
    .Y(_04528_));
 sky130_as_sc_hs__nand3_2 _35259_ (.A(_04526_),
    .B(_04528_),
    .C(_04529_),
    .Y(_04531_));
 sky130_as_sc_hs__or2_2 _35260_ (.A(_04448_),
    .B(_04488_),
    .Y(_04532_));
 sky130_as_sc_hs__nand3_2 _35262_ (.A(_04466_),
    .B(_04467_),
    .C(_04533_),
    .Y(_04534_));
 sky130_as_sc_hs__nand3_2 _35264_ (.A(_04442_),
    .B(_04443_),
    .C(_04535_),
    .Y(_04536_));
 sky130_as_sc_hs__or2_2 _35266_ (.A(_04365_),
    .B(_04400_),
    .Y(_04538_));
 sky130_as_sc_hs__and2_2 _35267_ (.A(_04401_),
    .B(_04538_),
    .Y(_04539_));
 sky130_as_sc_hs__or2_2 _35270_ (.A(_04303_),
    .B(_04362_),
    .Y(_04542_));
 sky130_as_sc_hs__or2_2 _35275_ (.A(_04166_),
    .B(_04231_),
    .Y(_04547_));
 sky130_as_sc_hs__or2_2 _35278_ (.A(_04077_),
    .B(_04163_),
    .Y(_04550_));
 sky130_as_sc_hs__and2_2 _35279_ (.A(_04164_),
    .B(_04550_),
    .Y(_04551_));
 sky130_as_sc_hs__and2_2 _35281_ (.A(_04164_),
    .B(_04552_),
    .Y(_04553_));
 sky130_as_sc_hs__nand3_2 _35282_ (.A(_04075_),
    .B(_04164_),
    .C(_04552_),
    .Y(_04554_));
 sky130_as_sc_hs__and2_2 _35283_ (.A(_04074_),
    .B(_04554_),
    .Y(_04555_));
 sky130_as_sc_hs__or2_2 _35284_ (.A(_03462_),
    .B(_03464_),
    .Y(_04556_));
 sky130_as_sc_hs__or2_2 _35286_ (.A(_03317_),
    .B(_03339_),
    .Y(_04558_));
 sky130_as_sc_hs__or2_2 _35288_ (.A(_03171_),
    .B(_03172_),
    .Y(_04560_));
 sky130_as_sc_hs__and2_2 _35289_ (.A(_03173_),
    .B(_04560_),
    .Y(_04561_));
 sky130_as_sc_hs__or2_2 _35290_ (.A(_03332_),
    .B(_03334_),
    .Y(_04562_));
 sky130_as_sc_hs__and2_2 _35291_ (.A(_03335_),
    .B(_04562_),
    .Y(_04563_));
 sky130_as_sc_hs__nand3_2 _35292_ (.A(net458),
    .B(_24535_),
    .C(_24536_),
    .Y(_04564_));
 sky130_as_sc_hs__or2_2 _35294_ (.A(_04564_),
    .B(_04565_),
    .Y(_04566_));
 sky130_as_sc_hs__and2_2 _35295_ (.A(net90),
    .B(net87),
    .Y(_04567_));
 sky130_as_sc_hs__and2_2 _35297_ (.A(_04566_),
    .B(_04568_),
    .Y(_04569_));
 sky130_as_sc_hs__or2_2 _35300_ (.A(_03323_),
    .B(_03325_),
    .Y(_04572_));
 sky130_as_sc_hs__and2_2 _35301_ (.A(_03326_),
    .B(_04572_),
    .Y(_04573_));
 sky130_as_sc_hs__or2_2 _35303_ (.A(_03348_),
    .B(_03349_),
    .Y(_04575_));
 sky130_as_sc_hs__and2_2 _35304_ (.A(_03350_),
    .B(_04575_),
    .Y(_04576_));
 sky130_as_sc_hs__or2_2 _35305_ (.A(_04571_),
    .B(_04573_),
    .Y(_04577_));
 sky130_as_sc_hs__and2_2 _35306_ (.A(_04574_),
    .B(_04577_),
    .Y(_04578_));
 sky130_as_sc_hs__or2_2 _35310_ (.A(_04563_),
    .B(_04580_),
    .Y(_04582_));
 sky130_as_sc_hs__and2_2 _35311_ (.A(_04581_),
    .B(_04582_),
    .Y(_04583_));
 sky130_as_sc_hs__or2_2 _35313_ (.A(_04559_),
    .B(_04584_),
    .Y(_04585_));
 sky130_as_sc_hs__and2_2 _35315_ (.A(_04585_),
    .B(_04586_),
    .Y(_04587_));
 sky130_as_sc_hs__and2_2 _35317_ (.A(_03357_),
    .B(_04588_),
    .Y(_04589_));
 sky130_as_sc_hs__or2_2 _35318_ (.A(_03354_),
    .B(_03355_),
    .Y(_04590_));
 sky130_as_sc_hs__and2_2 _35320_ (.A(_24053_),
    .B(net448),
    .Y(_04592_));
 sky130_as_sc_hs__and2_2 _35321_ (.A(_23712_),
    .B(net450),
    .Y(_04593_));
 sky130_as_sc_hs__or2_2 _35323_ (.A(_04591_),
    .B(_04594_),
    .Y(_04595_));
 sky130_as_sc_hs__and2_2 _35326_ (.A(_24216_),
    .B(net445),
    .Y(_04598_));
 sky130_as_sc_hs__and2_2 _35327_ (.A(_24256_),
    .B(_24729_),
    .Y(_04599_));
 sky130_as_sc_hs__or2_2 _35329_ (.A(_04597_),
    .B(_04600_),
    .Y(_04601_));
 sky130_as_sc_hs__or2_2 _35332_ (.A(_04589_),
    .B(_04602_),
    .Y(_04604_));
 sky130_as_sc_hs__and2_2 _35333_ (.A(_04603_),
    .B(_04604_),
    .Y(_04605_));
 sky130_as_sc_hs__or2_2 _35334_ (.A(_03390_),
    .B(_03392_),
    .Y(_04606_));
 sky130_as_sc_hs__and2_2 _35335_ (.A(_03393_),
    .B(_04606_),
    .Y(_04607_));
 sky130_as_sc_hs__or2_2 _35338_ (.A(_03361_),
    .B(_03363_),
    .Y(_04610_));
 sky130_as_sc_hs__or2_2 _35340_ (.A(_04581_),
    .B(_04611_),
    .Y(_04612_));
 sky130_as_sc_hs__and2_2 _35342_ (.A(_04612_),
    .B(_04613_),
    .Y(_04614_));
 sky130_as_sc_hs__or2_2 _35344_ (.A(_04609_),
    .B(_04614_),
    .Y(_04616_));
 sky130_as_sc_hs__and2_2 _35345_ (.A(_04615_),
    .B(_04616_),
    .Y(_04617_));
 sky130_as_sc_hs__or2_2 _35348_ (.A(_03343_),
    .B(_03373_),
    .Y(_04620_));
 sky130_as_sc_hs__and2_2 _35349_ (.A(_03374_),
    .B(_04620_),
    .Y(_04621_));
 sky130_as_sc_hs__or2_2 _35351_ (.A(_04619_),
    .B(_04621_),
    .Y(_04623_));
 sky130_as_sc_hs__and2_2 _35352_ (.A(_04622_),
    .B(_04623_),
    .Y(_04624_));
 sky130_as_sc_hs__or2_2 _35353_ (.A(_03410_),
    .B(_03412_),
    .Y(_04625_));
 sky130_as_sc_hs__and2_2 _35354_ (.A(_03413_),
    .B(_04625_),
    .Y(_04626_));
 sky130_as_sc_hs__or2_2 _35355_ (.A(_03385_),
    .B(_03386_),
    .Y(_04627_));
 sky130_as_sc_hs__and2_2 _35357_ (.A(_24545_),
    .B(_24774_),
    .Y(_04629_));
 sky130_as_sc_hs__and2_2 _35358_ (.A(net86),
    .B(_24768_),
    .Y(_04630_));
 sky130_as_sc_hs__or2_2 _35360_ (.A(_04628_),
    .B(_04631_),
    .Y(_04632_));
 sky130_as_sc_hs__or2_2 _35361_ (.A(_03400_),
    .B(_03401_),
    .Y(_04633_));
 sky130_as_sc_hs__and2_2 _35362_ (.A(_03402_),
    .B(_04633_),
    .Y(_04634_));
 sky130_as_sc_hs__and2_2 _35364_ (.A(_04632_),
    .B(_04635_),
    .Y(_04636_));
 sky130_as_sc_hs__and2_2 _35368_ (.A(_03409_),
    .B(_04639_),
    .Y(_04640_));
 sky130_as_sc_hs__nand2b_2 _35370_ (.B(_03407_),
    .Y(_04642_),
    .A(_03406_));
 sky130_as_sc_hs__and2_2 _35372_ (.A(net453),
    .B(_24814_),
    .Y(_04644_));
 sky130_as_sc_hs__and2_2 _35373_ (.A(net447),
    .B(_24808_),
    .Y(_04645_));
 sky130_as_sc_hs__or2_2 _35375_ (.A(_04643_),
    .B(_04646_),
    .Y(_04647_));
 sky130_as_sc_hs__and2_2 _35378_ (.A(net79),
    .B(_25211_),
    .Y(_04650_));
 sky130_as_sc_hs__and2_2 _35379_ (.A(net443),
    .B(_25205_),
    .Y(_04651_));
 sky130_as_sc_hs__or2_2 _35381_ (.A(_04649_),
    .B(_04652_),
    .Y(_04653_));
 sky130_as_sc_hs__or2_2 _35383_ (.A(_04638_),
    .B(_04640_),
    .Y(_04655_));
 sky130_as_sc_hs__and2_2 _35384_ (.A(_04641_),
    .B(_04655_),
    .Y(_04656_));
 sky130_as_sc_hs__or2_2 _35388_ (.A(_04626_),
    .B(_04658_),
    .Y(_04660_));
 sky130_as_sc_hs__and2_2 _35389_ (.A(_04659_),
    .B(_04660_),
    .Y(_04661_));
 sky130_as_sc_hs__and2_2 _35390_ (.A(_23702_),
    .B(net86),
    .Y(_04662_));
 sky130_as_sc_hs__or2_2 _35391_ (.A(_03427_),
    .B(_03429_),
    .Y(_04663_));
 sky130_as_sc_hs__and2_2 _35392_ (.A(_03430_),
    .B(_04663_),
    .Y(_04664_));
 sky130_as_sc_hs__or2_2 _35393_ (.A(_03423_),
    .B(_03424_),
    .Y(_04665_));
 sky130_as_sc_hs__and2_2 _35395_ (.A(net482),
    .B(_24256_),
    .Y(_04667_));
 sky130_as_sc_hs__and2_2 _35396_ (.A(_23636_),
    .B(net85),
    .Y(_04668_));
 sky130_as_sc_hs__or2_2 _35398_ (.A(_04666_),
    .B(_04669_),
    .Y(_04670_));
 sky130_as_sc_hs__and2_2 _35399_ (.A(net114),
    .B(net477),
    .Y(_04671_));
 sky130_as_sc_hs__and2_2 _35401_ (.A(_04670_),
    .B(_04672_),
    .Y(_04673_));
 sky130_as_sc_hs__or2_2 _35405_ (.A(_04664_),
    .B(_04675_),
    .Y(_04677_));
 sky130_as_sc_hs__and2_2 _35406_ (.A(_04676_),
    .B(_04677_),
    .Y(_04678_));
 sky130_as_sc_hs__or2_2 _35408_ (.A(_04662_),
    .B(_04678_),
    .Y(_04680_));
 sky130_as_sc_hs__and2_2 _35409_ (.A(_04679_),
    .B(_04680_),
    .Y(_04681_));
 sky130_as_sc_hs__or2_2 _35413_ (.A(_03417_),
    .B(_03437_),
    .Y(_04685_));
 sky130_as_sc_hs__and2_2 _35414_ (.A(_03438_),
    .B(_04685_),
    .Y(_04686_));
 sky130_as_sc_hs__or2_2 _35416_ (.A(_04684_),
    .B(_04686_),
    .Y(_04688_));
 sky130_as_sc_hs__and2_2 _35417_ (.A(_04687_),
    .B(_04688_),
    .Y(_04689_));
 sky130_as_sc_hs__or2_2 _35419_ (.A(_04683_),
    .B(_04689_),
    .Y(_04691_));
 sky130_as_sc_hs__and2_2 _35420_ (.A(_04690_),
    .B(_04691_),
    .Y(_04692_));
 sky130_as_sc_hs__or2_2 _35423_ (.A(_03380_),
    .B(_03448_),
    .Y(_04695_));
 sky130_as_sc_hs__and2_2 _35424_ (.A(_03449_),
    .B(_04695_),
    .Y(_04696_));
 sky130_as_sc_hs__or2_2 _35427_ (.A(_04694_),
    .B(_04696_),
    .Y(_04699_));
 sky130_as_sc_hs__and2_2 _35428_ (.A(_04697_),
    .B(_04699_),
    .Y(_04700_));
 sky130_as_sc_hs__or2_2 _35431_ (.A(_03454_),
    .B(_03456_),
    .Y(_04703_));
 sky130_as_sc_hs__and2_2 _35432_ (.A(_03457_),
    .B(_04703_),
    .Y(_04704_));
 sky130_as_sc_hs__or2_2 _35435_ (.A(_04702_),
    .B(_04704_),
    .Y(_04707_));
 sky130_as_sc_hs__and2_2 _35436_ (.A(_04705_),
    .B(_04707_),
    .Y(_04708_));
 sky130_as_sc_hs__and2_2 _35438_ (.A(_04705_),
    .B(_04709_),
    .Y(_04710_));
 sky130_as_sc_hs__or2_2 _35439_ (.A(_04557_),
    .B(_04710_),
    .Y(_04711_));
 sky130_as_sc_hs__and2_2 _35441_ (.A(_04711_),
    .B(_04712_),
    .Y(_04713_));
 sky130_as_sc_hs__or2_2 _35442_ (.A(_04706_),
    .B(_04708_),
    .Y(_04714_));
 sky130_as_sc_hs__and2_2 _35443_ (.A(_04709_),
    .B(_04714_),
    .Y(_04715_));
 sky130_as_sc_hs__or2_2 _35444_ (.A(_04561_),
    .B(_04583_),
    .Y(_04716_));
 sky130_as_sc_hs__and2_2 _35446_ (.A(net113),
    .B(net461),
    .Y(_04718_));
 sky130_as_sc_hs__or2_2 _35447_ (.A(_04576_),
    .B(_04578_),
    .Y(_04719_));
 sky130_as_sc_hs__and2_2 _35448_ (.A(_04579_),
    .B(_04719_),
    .Y(_04720_));
 sky130_as_sc_hs__or2_2 _35449_ (.A(_04567_),
    .B(_04569_),
    .Y(_04721_));
 sky130_as_sc_hs__or2_2 _35451_ (.A(_03848_),
    .B(_04722_),
    .Y(_04723_));
 sky130_as_sc_hs__and2_2 _35453_ (.A(_04723_),
    .B(_04724_),
    .Y(_04725_));
 sky130_as_sc_hs__or2_2 _35454_ (.A(_04592_),
    .B(_04593_),
    .Y(_04726_));
 sky130_as_sc_hs__and2_2 _35455_ (.A(_04594_),
    .B(_04726_),
    .Y(_04727_));
 sky130_as_sc_hs__or2_2 _35459_ (.A(_04720_),
    .B(_04729_),
    .Y(_04731_));
 sky130_as_sc_hs__and2_2 _35460_ (.A(_04730_),
    .B(_04731_),
    .Y(_04732_));
 sky130_as_sc_hs__or2_2 _35462_ (.A(_04717_),
    .B(_04733_),
    .Y(_04734_));
 sky130_as_sc_hs__and2_2 _35464_ (.A(_04734_),
    .B(_04735_),
    .Y(_04736_));
 sky130_as_sc_hs__and2_2 _35466_ (.A(_04601_),
    .B(_04737_),
    .Y(_04738_));
 sky130_as_sc_hs__or2_2 _35467_ (.A(_04598_),
    .B(_04599_),
    .Y(_04739_));
 sky130_as_sc_hs__or2_2 _35469_ (.A(_03843_),
    .B(_04740_),
    .Y(_04741_));
 sky130_as_sc_hs__or2_2 _35472_ (.A(_03819_),
    .B(_04743_),
    .Y(_04744_));
 sky130_as_sc_hs__or2_2 _35475_ (.A(_04738_),
    .B(_04745_),
    .Y(_04747_));
 sky130_as_sc_hs__and2_2 _35476_ (.A(_04746_),
    .B(_04747_),
    .Y(_04748_));
 sky130_as_sc_hs__or2_2 _35477_ (.A(_04634_),
    .B(_04636_),
    .Y(_04749_));
 sky130_as_sc_hs__and2_2 _35478_ (.A(_04637_),
    .B(_04749_),
    .Y(_04750_));
 sky130_as_sc_hs__or2_2 _35481_ (.A(_04605_),
    .B(_04607_),
    .Y(_04753_));
 sky130_as_sc_hs__or2_2 _35483_ (.A(_04730_),
    .B(_04754_),
    .Y(_04755_));
 sky130_as_sc_hs__and2_2 _35485_ (.A(_04755_),
    .B(_04756_),
    .Y(_04757_));
 sky130_as_sc_hs__or2_2 _35487_ (.A(_04752_),
    .B(_04757_),
    .Y(_04759_));
 sky130_as_sc_hs__and2_2 _35488_ (.A(_04758_),
    .B(_04759_),
    .Y(_04760_));
 sky130_as_sc_hs__or2_2 _35491_ (.A(_04587_),
    .B(_04617_),
    .Y(_04763_));
 sky130_as_sc_hs__and2_2 _35492_ (.A(_04618_),
    .B(_04763_),
    .Y(_04764_));
 sky130_as_sc_hs__or2_2 _35494_ (.A(_04762_),
    .B(_04764_),
    .Y(_04766_));
 sky130_as_sc_hs__and2_2 _35495_ (.A(_04765_),
    .B(_04766_),
    .Y(_04767_));
 sky130_as_sc_hs__or2_2 _35496_ (.A(_04654_),
    .B(_04656_),
    .Y(_04768_));
 sky130_as_sc_hs__and2_2 _35497_ (.A(_04657_),
    .B(_04768_),
    .Y(_04769_));
 sky130_as_sc_hs__or2_2 _35498_ (.A(_04629_),
    .B(_04630_),
    .Y(_04770_));
 sky130_as_sc_hs__or2_2 _35500_ (.A(_03808_),
    .B(_04771_),
    .Y(_04772_));
 sky130_as_sc_hs__or2_2 _35501_ (.A(_04644_),
    .B(_04645_),
    .Y(_04773_));
 sky130_as_sc_hs__and2_2 _35502_ (.A(_04646_),
    .B(_04773_),
    .Y(_04774_));
 sky130_as_sc_hs__and2_2 _35504_ (.A(_04772_),
    .B(_04775_),
    .Y(_04776_));
 sky130_as_sc_hs__and2_2 _35508_ (.A(_04653_),
    .B(_04779_),
    .Y(_04780_));
 sky130_as_sc_hs__or2_2 _35510_ (.A(_04650_),
    .B(_04651_),
    .Y(_04782_));
 sky130_as_sc_hs__or2_2 _35512_ (.A(_03803_),
    .B(_04783_),
    .Y(_04784_));
 sky130_as_sc_hs__or2_2 _35515_ (.A(_03739_),
    .B(_04786_),
    .Y(_04787_));
 sky130_as_sc_hs__or2_2 _35517_ (.A(_04778_),
    .B(_04780_),
    .Y(_04789_));
 sky130_as_sc_hs__and2_2 _35518_ (.A(_04781_),
    .B(_04789_),
    .Y(_04790_));
 sky130_as_sc_hs__or2_2 _35522_ (.A(_04769_),
    .B(_04792_),
    .Y(_04794_));
 sky130_as_sc_hs__and2_2 _35523_ (.A(_04793_),
    .B(_04794_),
    .Y(_04795_));
 sky130_as_sc_hs__and2_2 _35524_ (.A(_23702_),
    .B(net455),
    .Y(_04796_));
 sky130_as_sc_hs__or2_2 _35525_ (.A(_04671_),
    .B(_04673_),
    .Y(_04797_));
 sky130_as_sc_hs__and2_2 _35526_ (.A(_04674_),
    .B(_04797_),
    .Y(_04798_));
 sky130_as_sc_hs__or2_2 _35527_ (.A(_04667_),
    .B(_04668_),
    .Y(_04799_));
 sky130_as_sc_hs__and2_2 _35529_ (.A(net483),
    .B(_24229_),
    .Y(_04801_));
 sky130_as_sc_hs__and2_2 _35530_ (.A(_23636_),
    .B(net454),
    .Y(_04802_));
 sky130_as_sc_hs__or2_2 _35532_ (.A(_04800_),
    .B(_04803_),
    .Y(_04804_));
 sky130_as_sc_hs__and2_2 _35533_ (.A(net114),
    .B(net481),
    .Y(_04805_));
 sky130_as_sc_hs__and2_2 _35535_ (.A(_04804_),
    .B(_04806_),
    .Y(_04807_));
 sky130_as_sc_hs__or2_2 _35539_ (.A(_04798_),
    .B(_04809_),
    .Y(_04811_));
 sky130_as_sc_hs__and2_2 _35540_ (.A(_04810_),
    .B(_04811_),
    .Y(_04812_));
 sky130_as_sc_hs__or2_2 _35542_ (.A(_04796_),
    .B(_04812_),
    .Y(_04814_));
 sky130_as_sc_hs__and2_2 _35543_ (.A(_04813_),
    .B(_04814_),
    .Y(_04815_));
 sky130_as_sc_hs__or2_2 _35547_ (.A(_04661_),
    .B(_04681_),
    .Y(_04819_));
 sky130_as_sc_hs__and2_2 _35548_ (.A(_04682_),
    .B(_04819_),
    .Y(_04820_));
 sky130_as_sc_hs__or2_2 _35550_ (.A(_04818_),
    .B(_04820_),
    .Y(_04822_));
 sky130_as_sc_hs__and2_2 _35551_ (.A(_04821_),
    .B(_04822_),
    .Y(_04823_));
 sky130_as_sc_hs__or2_2 _35553_ (.A(_04817_),
    .B(_04823_),
    .Y(_04825_));
 sky130_as_sc_hs__and2_2 _35554_ (.A(_04824_),
    .B(_04825_),
    .Y(_04826_));
 sky130_as_sc_hs__or2_2 _35557_ (.A(_04624_),
    .B(_04692_),
    .Y(_04829_));
 sky130_as_sc_hs__and2_2 _35558_ (.A(_04693_),
    .B(_04829_),
    .Y(_04830_));
 sky130_as_sc_hs__or2_2 _35561_ (.A(_04828_),
    .B(_04830_),
    .Y(_04833_));
 sky130_as_sc_hs__and2_2 _35562_ (.A(_04831_),
    .B(_04833_),
    .Y(_04834_));
 sky130_as_sc_hs__or2_2 _35565_ (.A(_04698_),
    .B(_04700_),
    .Y(_04837_));
 sky130_as_sc_hs__and2_2 _35566_ (.A(_04701_),
    .B(_04837_),
    .Y(_04838_));
 sky130_as_sc_hs__or2_2 _35569_ (.A(_04836_),
    .B(_04838_),
    .Y(_04841_));
 sky130_as_sc_hs__and2_2 _35570_ (.A(_04839_),
    .B(_04841_),
    .Y(_04842_));
 sky130_as_sc_hs__or2_2 _35574_ (.A(_04715_),
    .B(_04844_),
    .Y(_04846_));
 sky130_as_sc_hs__and2_2 _35575_ (.A(_04845_),
    .B(_04846_),
    .Y(_04847_));
 sky130_as_sc_hs__and2_2 _35576_ (.A(_04713_),
    .B(_04847_),
    .Y(_04848_));
 sky130_as_sc_hs__or2_2 _35577_ (.A(_04840_),
    .B(_04842_),
    .Y(_04849_));
 sky130_as_sc_hs__or2_2 _35579_ (.A(_04736_),
    .B(_04760_),
    .Y(_04851_));
 sky130_as_sc_hs__and2_2 _35582_ (.A(_04744_),
    .B(_04853_),
    .Y(_04854_));
 sky130_as_sc_hs__or2_2 _35585_ (.A(_04854_),
    .B(_04855_),
    .Y(_04857_));
 sky130_as_sc_hs__and2_2 _35586_ (.A(_04856_),
    .B(_04857_),
    .Y(_04858_));
 sky130_as_sc_hs__or2_2 _35587_ (.A(_04774_),
    .B(_04776_),
    .Y(_04859_));
 sky130_as_sc_hs__and2_2 _35588_ (.A(_04777_),
    .B(_04859_),
    .Y(_04860_));
 sky130_as_sc_hs__or2_2 _35591_ (.A(_04725_),
    .B(_04727_),
    .Y(_04863_));
 sky130_as_sc_hs__or2_2 _35593_ (.A(_03851_),
    .B(_04864_),
    .Y(_04865_));
 sky130_as_sc_hs__or2_2 _35594_ (.A(_04748_),
    .B(_04750_),
    .Y(_04866_));
 sky130_as_sc_hs__or2_2 _35596_ (.A(_04865_),
    .B(_04867_),
    .Y(_04868_));
 sky130_as_sc_hs__and2_2 _35598_ (.A(_04868_),
    .B(_04869_),
    .Y(_04870_));
 sky130_as_sc_hs__or2_2 _35600_ (.A(_04862_),
    .B(_04870_),
    .Y(_04872_));
 sky130_as_sc_hs__and2_2 _35601_ (.A(_04871_),
    .B(_04872_),
    .Y(_04873_));
 sky130_as_sc_hs__or2_2 _35602_ (.A(_04718_),
    .B(_04732_),
    .Y(_04874_));
 sky130_as_sc_hs__and2_2 _35603_ (.A(_04733_),
    .B(_04874_),
    .Y(_04875_));
 sky130_as_sc_hs__or2_2 _35605_ (.A(_04852_),
    .B(_04876_),
    .Y(_04877_));
 sky130_as_sc_hs__and2_2 _35607_ (.A(_04877_),
    .B(_04878_),
    .Y(_04879_));
 sky130_as_sc_hs__or2_2 _35609_ (.A(_04795_),
    .B(_04815_),
    .Y(_04881_));
 sky130_as_sc_hs__and2_2 _35610_ (.A(_04816_),
    .B(_04881_),
    .Y(_04882_));
 sky130_as_sc_hs__or2_2 _35612_ (.A(_04880_),
    .B(_04882_),
    .Y(_04884_));
 sky130_as_sc_hs__and2_2 _35613_ (.A(_04883_),
    .B(_04884_),
    .Y(_04885_));
 sky130_as_sc_hs__or2_2 _35614_ (.A(_04788_),
    .B(_04790_),
    .Y(_04886_));
 sky130_as_sc_hs__and2_2 _35615_ (.A(_04791_),
    .B(_04886_),
    .Y(_04887_));
 sky130_as_sc_hs__and2_2 _35618_ (.A(_04787_),
    .B(_04889_),
    .Y(_04890_));
 sky130_as_sc_hs__or2_2 _35621_ (.A(_04888_),
    .B(_04890_),
    .Y(_04893_));
 sky130_as_sc_hs__and2_2 _35622_ (.A(_04891_),
    .B(_04893_),
    .Y(_04894_));
 sky130_as_sc_hs__nand3_2 _35623_ (.A(_04891_),
    .B(_04892_),
    .C(_04893_),
    .Y(_04895_));
 sky130_as_sc_hs__or2_2 _35626_ (.A(_04887_),
    .B(_04896_),
    .Y(_04898_));
 sky130_as_sc_hs__and2_2 _35627_ (.A(_04897_),
    .B(_04898_),
    .Y(_04899_));
 sky130_as_sc_hs__and2_2 _35628_ (.A(_23702_),
    .B(_24545_),
    .Y(_04900_));
 sky130_as_sc_hs__or2_2 _35629_ (.A(_04805_),
    .B(_04807_),
    .Y(_04901_));
 sky130_as_sc_hs__and2_2 _35630_ (.A(_04808_),
    .B(_04901_),
    .Y(_04902_));
 sky130_as_sc_hs__or2_2 _35631_ (.A(_04801_),
    .B(_04802_),
    .Y(_04903_));
 sky130_as_sc_hs__or2_2 _35633_ (.A(_03763_),
    .B(_04904_),
    .Y(_04905_));
 sky130_as_sc_hs__and2_2 _35634_ (.A(net116),
    .B(_23674_),
    .Y(_04906_));
 sky130_as_sc_hs__and2_2 _35636_ (.A(_04905_),
    .B(_04907_),
    .Y(_04908_));
 sky130_as_sc_hs__or2_2 _35640_ (.A(_04902_),
    .B(_04910_),
    .Y(_04912_));
 sky130_as_sc_hs__and2_2 _35641_ (.A(_04911_),
    .B(_04912_),
    .Y(_04913_));
 sky130_as_sc_hs__or2_2 _35643_ (.A(_04900_),
    .B(_04913_),
    .Y(_04915_));
 sky130_as_sc_hs__and2_2 _35644_ (.A(_04914_),
    .B(_04915_),
    .Y(_04916_));
 sky130_as_sc_hs__or2_2 _35648_ (.A(_04885_),
    .B(_04918_),
    .Y(_04920_));
 sky130_as_sc_hs__and2_2 _35649_ (.A(_04919_),
    .B(_04920_),
    .Y(_04921_));
 sky130_as_sc_hs__or2_2 _35652_ (.A(_04767_),
    .B(_04826_),
    .Y(_04924_));
 sky130_as_sc_hs__and2_2 _35653_ (.A(_04827_),
    .B(_04924_),
    .Y(_04925_));
 sky130_as_sc_hs__or2_2 _35656_ (.A(_04923_),
    .B(_04925_),
    .Y(_04928_));
 sky130_as_sc_hs__and2_2 _35657_ (.A(_04926_),
    .B(_04928_),
    .Y(_04929_));
 sky130_as_sc_hs__or2_2 _35660_ (.A(_04832_),
    .B(_04834_),
    .Y(_04932_));
 sky130_as_sc_hs__and2_2 _35661_ (.A(_04835_),
    .B(_04932_),
    .Y(_04933_));
 sky130_as_sc_hs__or2_2 _35664_ (.A(_04931_),
    .B(_04933_),
    .Y(_04936_));
 sky130_as_sc_hs__and2_2 _35665_ (.A(_04934_),
    .B(_04936_),
    .Y(_04937_));
 sky130_as_sc_hs__and2_2 _35667_ (.A(_04934_),
    .B(_04938_),
    .Y(_04939_));
 sky130_as_sc_hs__or2_2 _35669_ (.A(_04850_),
    .B(_04939_),
    .Y(_04941_));
 sky130_as_sc_hs__and2_2 _35670_ (.A(_04940_),
    .B(_04941_),
    .Y(_04942_));
 sky130_as_sc_hs__or2_2 _35671_ (.A(_04935_),
    .B(_04937_),
    .Y(_04943_));
 sky130_as_sc_hs__and2_2 _35672_ (.A(_04938_),
    .B(_04943_),
    .Y(_04944_));
 sky130_as_sc_hs__or2_2 _35673_ (.A(_04873_),
    .B(_04875_),
    .Y(_04945_));
 sky130_as_sc_hs__or2_2 _35676_ (.A(_04858_),
    .B(_04860_),
    .Y(_04948_));
 sky130_as_sc_hs__or2_2 _35678_ (.A(_03854_),
    .B(_04949_),
    .Y(_04950_));
 sky130_as_sc_hs__and2_2 _35680_ (.A(_04950_),
    .B(_04951_),
    .Y(_04952_));
 sky130_as_sc_hs__or2_2 _35682_ (.A(_04947_),
    .B(_04952_),
    .Y(_04954_));
 sky130_as_sc_hs__and2_2 _35683_ (.A(_04953_),
    .B(_04954_),
    .Y(_04955_));
 sky130_as_sc_hs__and2_2 _35685_ (.A(_04865_),
    .B(_04956_),
    .Y(_04957_));
 sky130_as_sc_hs__or2_2 _35687_ (.A(_04946_),
    .B(_04958_),
    .Y(_04959_));
 sky130_as_sc_hs__and2_2 _35689_ (.A(_04959_),
    .B(_04960_),
    .Y(_04961_));
 sky130_as_sc_hs__or2_2 _35691_ (.A(_04899_),
    .B(_04916_),
    .Y(_04963_));
 sky130_as_sc_hs__and2_2 _35692_ (.A(_04917_),
    .B(_04963_),
    .Y(_04964_));
 sky130_as_sc_hs__or2_2 _35694_ (.A(_04962_),
    .B(_04964_),
    .Y(_04966_));
 sky130_as_sc_hs__and2_2 _35695_ (.A(_04965_),
    .B(_04966_),
    .Y(_04967_));
 sky130_as_sc_hs__or2_2 _35696_ (.A(_04892_),
    .B(_04894_),
    .Y(_04968_));
 sky130_as_sc_hs__and2_2 _35697_ (.A(_04895_),
    .B(_04968_),
    .Y(_04969_));
 sky130_as_sc_hs__or2_2 _35700_ (.A(_04969_),
    .B(_04970_),
    .Y(_04972_));
 sky130_as_sc_hs__and2_2 _35701_ (.A(_04971_),
    .B(_04972_),
    .Y(_04973_));
 sky130_as_sc_hs__and2_2 _35702_ (.A(_23702_),
    .B(_24501_),
    .Y(_04974_));
 sky130_as_sc_hs__or2_2 _35703_ (.A(_04906_),
    .B(_04908_),
    .Y(_04975_));
 sky130_as_sc_hs__and2_2 _35704_ (.A(_04909_),
    .B(_04975_),
    .Y(_04976_));
 sky130_as_sc_hs__or2_2 _35707_ (.A(_04976_),
    .B(_04977_),
    .Y(_04979_));
 sky130_as_sc_hs__and2_2 _35708_ (.A(_04978_),
    .B(_04979_),
    .Y(_04980_));
 sky130_as_sc_hs__or2_2 _35710_ (.A(_04974_),
    .B(_04980_),
    .Y(_04982_));
 sky130_as_sc_hs__and2_2 _35711_ (.A(_04981_),
    .B(_04982_),
    .Y(_04983_));
 sky130_as_sc_hs__or2_2 _35715_ (.A(_04967_),
    .B(_04985_),
    .Y(_04987_));
 sky130_as_sc_hs__and2_2 _35716_ (.A(_04986_),
    .B(_04987_),
    .Y(_04988_));
 sky130_as_sc_hs__or2_2 _35719_ (.A(_04879_),
    .B(_04921_),
    .Y(_04991_));
 sky130_as_sc_hs__and2_2 _35720_ (.A(_04922_),
    .B(_04991_),
    .Y(_04992_));
 sky130_as_sc_hs__or2_2 _35723_ (.A(_04990_),
    .B(_04992_),
    .Y(_04995_));
 sky130_as_sc_hs__and2_2 _35724_ (.A(_04993_),
    .B(_04995_),
    .Y(_04996_));
 sky130_as_sc_hs__or2_2 _35727_ (.A(_04927_),
    .B(_04929_),
    .Y(_04999_));
 sky130_as_sc_hs__and2_2 _35728_ (.A(_04930_),
    .B(_04999_),
    .Y(_05000_));
 sky130_as_sc_hs__or2_2 _35731_ (.A(_04998_),
    .B(_05000_),
    .Y(_05003_));
 sky130_as_sc_hs__and2_2 _35732_ (.A(_05001_),
    .B(_05003_),
    .Y(_05004_));
 sky130_as_sc_hs__or2_2 _35736_ (.A(_04944_),
    .B(_05006_),
    .Y(_05008_));
 sky130_as_sc_hs__and2_2 _35737_ (.A(_05007_),
    .B(_05008_),
    .Y(_05009_));
 sky130_as_sc_hs__and2_2 _35738_ (.A(_04942_),
    .B(_05009_),
    .Y(_05010_));
 sky130_as_sc_hs__and2_2 _35739_ (.A(_04848_),
    .B(_05010_),
    .Y(_05011_));
 sky130_as_sc_hs__or2_2 _35740_ (.A(_05002_),
    .B(_05004_),
    .Y(_05012_));
 sky130_as_sc_hs__or2_2 _35742_ (.A(_04994_),
    .B(_04996_),
    .Y(_05014_));
 sky130_as_sc_hs__and2_2 _35743_ (.A(_04997_),
    .B(_05014_),
    .Y(_05015_));
 sky130_as_sc_hs__or2_2 _35744_ (.A(_04961_),
    .B(_04988_),
    .Y(_05016_));
 sky130_as_sc_hs__and2_2 _35745_ (.A(_04989_),
    .B(_05016_),
    .Y(_05017_));
 sky130_as_sc_hs__or2_2 _35746_ (.A(_04955_),
    .B(_04957_),
    .Y(_05018_));
 sky130_as_sc_hs__or2_2 _35748_ (.A(_03857_),
    .B(_05019_),
    .Y(_05020_));
 sky130_as_sc_hs__or2_2 _35749_ (.A(_04973_),
    .B(_04983_),
    .Y(_05021_));
 sky130_as_sc_hs__or2_2 _35751_ (.A(_03838_),
    .B(_05022_),
    .Y(_05023_));
 sky130_as_sc_hs__and2_2 _35753_ (.A(_05023_),
    .B(_05024_),
    .Y(_05025_));
 sky130_as_sc_hs__or2_2 _35756_ (.A(_05025_),
    .B(_05026_),
    .Y(_05028_));
 sky130_as_sc_hs__and2_2 _35757_ (.A(_05027_),
    .B(_05028_),
    .Y(_05029_));
 sky130_as_sc_hs__and2_2 _35759_ (.A(_05020_),
    .B(_05030_),
    .Y(_05031_));
 sky130_as_sc_hs__or2_2 _35764_ (.A(_05017_),
    .B(_05033_),
    .Y(_05036_));
 sky130_as_sc_hs__and2_2 _35765_ (.A(_05034_),
    .B(_05036_),
    .Y(_05037_));
 sky130_as_sc_hs__nand3_2 _35766_ (.A(_05034_),
    .B(_05035_),
    .C(_05036_),
    .Y(_05038_));
 sky130_as_sc_hs__or2_2 _35770_ (.A(_05015_),
    .B(_05039_),
    .Y(_05042_));
 sky130_as_sc_hs__and2_2 _35771_ (.A(_05040_),
    .B(_05042_),
    .Y(_05043_));
 sky130_as_sc_hs__and2_2 _35773_ (.A(_05040_),
    .B(_05044_),
    .Y(_05045_));
 sky130_as_sc_hs__or2_2 _35774_ (.A(_05013_),
    .B(_05045_),
    .Y(_05046_));
 sky130_as_sc_hs__and2_2 _35776_ (.A(_05046_),
    .B(_05047_),
    .Y(_05048_));
 sky130_as_sc_hs__or2_2 _35777_ (.A(_05041_),
    .B(_05043_),
    .Y(_05049_));
 sky130_as_sc_hs__and2_2 _35778_ (.A(_05044_),
    .B(_05049_),
    .Y(_05050_));
 sky130_as_sc_hs__or2_2 _35779_ (.A(_05035_),
    .B(_05037_),
    .Y(_05051_));
 sky130_as_sc_hs__and2_2 _35780_ (.A(_05038_),
    .B(_05051_),
    .Y(_05052_));
 sky130_as_sc_hs__or2_2 _35781_ (.A(_05029_),
    .B(_05031_),
    .Y(_05053_));
 sky130_as_sc_hs__and2_2 _35782_ (.A(_05032_),
    .B(_05053_),
    .Y(_05054_));
 sky130_as_sc_hs__or2_2 _35786_ (.A(_05054_),
    .B(_05055_),
    .Y(_05058_));
 sky130_as_sc_hs__and2_2 _35787_ (.A(_05056_),
    .B(_05058_),
    .Y(_05059_));
 sky130_as_sc_hs__or2_2 _35792_ (.A(_05052_),
    .B(_05061_),
    .Y(_05064_));
 sky130_as_sc_hs__and2_2 _35793_ (.A(_05062_),
    .B(_05064_),
    .Y(_05065_));
 sky130_as_sc_hs__nand3_2 _35794_ (.A(_05062_),
    .B(_05063_),
    .C(_05064_),
    .Y(_05066_));
 sky130_as_sc_hs__or2_2 _35797_ (.A(_05050_),
    .B(_05067_),
    .Y(_05069_));
 sky130_as_sc_hs__and2_2 _35798_ (.A(_05068_),
    .B(_05069_),
    .Y(_05070_));
 sky130_as_sc_hs__and2_2 _35799_ (.A(_05048_),
    .B(_05070_),
    .Y(_05071_));
 sky130_as_sc_hs__or2_2 _35800_ (.A(_05063_),
    .B(_05065_),
    .Y(_05072_));
 sky130_as_sc_hs__and2_2 _35801_ (.A(_05066_),
    .B(_05072_),
    .Y(_05073_));
 sky130_as_sc_hs__or2_2 _35802_ (.A(_05057_),
    .B(_05059_),
    .Y(_05074_));
 sky130_as_sc_hs__and2_2 _35803_ (.A(_05060_),
    .B(_05074_),
    .Y(_05075_));
 sky130_as_sc_hs__or2_2 _35807_ (.A(_05075_),
    .B(_05076_),
    .Y(_05079_));
 sky130_as_sc_hs__and2_2 _35808_ (.A(_05077_),
    .B(_05079_),
    .Y(_05080_));
 sky130_as_sc_hs__nand3_2 _35809_ (.A(_05077_),
    .B(_05078_),
    .C(_05079_),
    .Y(_05081_));
 sky130_as_sc_hs__or2_2 _35811_ (.A(_05073_),
    .B(_05082_),
    .Y(_05083_));
 sky130_as_sc_hs__nand3_2 _35812_ (.A(_05066_),
    .B(_05072_),
    .C(_05082_),
    .Y(_05084_));
 sky130_as_sc_hs__and2_2 _35813_ (.A(_05083_),
    .B(_05084_),
    .Y(_05085_));
 sky130_as_sc_hs__or2_2 _35814_ (.A(_05078_),
    .B(_05080_),
    .Y(_05086_));
 sky130_as_sc_hs__and2_2 _35815_ (.A(_05081_),
    .B(_05086_),
    .Y(_05087_));
 sky130_as_sc_hs__nand3_2 _35817_ (.A(_05081_),
    .B(_05086_),
    .C(_05088_),
    .Y(_05089_));
 sky130_as_sc_hs__or2_2 _35818_ (.A(_05087_),
    .B(_05088_),
    .Y(_05090_));
 sky130_as_sc_hs__and2_2 _35819_ (.A(_05089_),
    .B(_05090_),
    .Y(_05091_));
 sky130_as_sc_hs__and2_2 _35820_ (.A(_05085_),
    .B(_05091_),
    .Y(_05092_));
 sky130_as_sc_hs__and2_2 _35821_ (.A(_05071_),
    .B(_05092_),
    .Y(_05093_));
 sky130_as_sc_hs__nand3_2 _35822_ (.A(_04555_),
    .B(_05011_),
    .C(_05093_),
    .Y(_05094_));
 sky130_as_sc_hs__and2_2 _35824_ (.A(_05083_),
    .B(_05095_),
    .Y(_05096_));
 sky130_as_sc_hs__nand2b_2 _35826_ (.B(_05047_),
    .Y(_05098_),
    .A(_05068_));
 sky130_as_sc_hs__nand3_2 _35827_ (.A(_05046_),
    .B(_05097_),
    .C(_05098_),
    .Y(_05099_));
 sky130_as_sc_hs__inv_2 _35828_ (.Y(_05100_),
    .A(_05099_));
 sky130_as_sc_hs__nand3_2 _35829_ (.A(_04848_),
    .B(_05010_),
    .C(_05099_),
    .Y(_05101_));
 sky130_as_sc_hs__and2_2 _35831_ (.A(_04940_),
    .B(_05102_),
    .Y(_05103_));
 sky130_as_sc_hs__nand2b_2 _35833_ (.B(_04712_),
    .Y(_05105_),
    .A(_04845_));
 sky130_as_sc_hs__and2_2 _35834_ (.A(_04711_),
    .B(_05105_),
    .Y(_05106_));
 sky130_as_sc_hs__nand3_2 _35835_ (.A(_05101_),
    .B(_05104_),
    .C(_05106_),
    .Y(_05107_));
 sky130_as_sc_hs__nand2b_2 _35836_ (.B(_05094_),
    .Y(_05108_),
    .A(_05107_));
 sky130_as_sc_hs__or2_2 _35839_ (.A(_02783_),
    .B(_05110_),
    .Y(_05111_));
 sky130_as_sc_hs__nand2b_2 _35840_ (.B(_02775_),
    .Y(_05112_),
    .A(_02780_));
 sky130_as_sc_hs__nand3_2 _35841_ (.A(_02774_),
    .B(_05111_),
    .C(_05112_),
    .Y(_05113_));
 sky130_as_sc_hs__nand3_2 _35843_ (.A(_03148_),
    .B(_03473_),
    .C(_05114_),
    .Y(_05115_));
 sky130_as_sc_hs__nand2b_2 _35844_ (.B(_02965_),
    .Y(_05116_),
    .A(_03145_));
 sky130_as_sc_hs__and2_2 _35845_ (.A(_02964_),
    .B(_05116_),
    .Y(_05117_));
 sky130_as_sc_hs__and2_2 _35846_ (.A(_05115_),
    .B(_05117_),
    .Y(_05118_));
 sky130_as_sc_hs__or2_2 _35847_ (.A(_02784_),
    .B(_05118_),
    .Y(_05119_));
 sky130_as_sc_hs__or2_2 _35848_ (.A(_03477_),
    .B(_05094_),
    .Y(_05120_));
 sky130_as_sc_hs__nor2b_2 _35849_ (.A(_03477_),
    .Y(_05121_),
    .B(_05107_));
 sky130_as_sc_hs__nor2_2 _35850_ (.A(_05113_),
    .B(_05121_),
    .Y(_05122_));
 sky130_as_sc_hs__nand3_2 _35851_ (.A(_05119_),
    .B(_05120_),
    .C(_05122_),
    .Y(_05123_));
 sky130_as_sc_hs__and2_2 _35856_ (.A(net483),
    .B(net475),
    .Y(_05128_));
 sky130_as_sc_hs__and2_2 _35857_ (.A(_23636_),
    .B(net428),
    .Y(_05129_));
 sky130_as_sc_hs__and2_2 _35858_ (.A(_24053_),
    .B(net422),
    .Y(_05130_));
 sky130_as_sc_hs__or2_2 _35859_ (.A(_05129_),
    .B(_05130_),
    .Y(_05131_));
 sky130_as_sc_hs__and2_2 _35861_ (.A(_05131_),
    .B(_05132_),
    .Y(_05133_));
 sky130_as_sc_hs__or2_2 _35863_ (.A(_05128_),
    .B(_05133_),
    .Y(_05135_));
 sky130_as_sc_hs__and2_2 _35864_ (.A(_05134_),
    .B(_05135_),
    .Y(_05136_));
 sky130_as_sc_hs__or2_2 _35867_ (.A(_05136_),
    .B(_05137_),
    .Y(_05139_));
 sky130_as_sc_hs__and2_2 _35868_ (.A(_05138_),
    .B(_05139_),
    .Y(_05140_));
 sky130_as_sc_hs__or2_2 _35871_ (.A(_05140_),
    .B(_05141_),
    .Y(_05143_));
 sky130_as_sc_hs__and2_2 _35872_ (.A(_05142_),
    .B(_05143_),
    .Y(_05144_));
 sky130_as_sc_hs__and2_2 _35873_ (.A(_23702_),
    .B(net432),
    .Y(_05145_));
 sky130_as_sc_hs__or2_2 _35875_ (.A(_05144_),
    .B(_05145_),
    .Y(_05147_));
 sky130_as_sc_hs__and2_2 _35876_ (.A(_05146_),
    .B(_05147_),
    .Y(_05148_));
 sky130_as_sc_hs__or2_2 _35884_ (.A(_05153_),
    .B(_05154_),
    .Y(_05156_));
 sky130_as_sc_hs__and2_2 _35885_ (.A(_05155_),
    .B(_05156_),
    .Y(_05157_));
 sky130_as_sc_hs__and2_2 _35886_ (.A(_25205_),
    .B(net75),
    .Y(_05158_));
 sky130_as_sc_hs__or2_2 _35888_ (.A(_05157_),
    .B(_05158_),
    .Y(_05160_));
 sky130_as_sc_hs__and2_2 _35889_ (.A(_05159_),
    .B(_05160_),
    .Y(_05161_));
 sky130_as_sc_hs__or2_2 _35891_ (.A(_05152_),
    .B(_05161_),
    .Y(_05163_));
 sky130_as_sc_hs__and2_2 _35892_ (.A(_05162_),
    .B(_05163_),
    .Y(_05164_));
 sky130_as_sc_hs__or2_2 _35894_ (.A(_05151_),
    .B(_05164_),
    .Y(_05166_));
 sky130_as_sc_hs__and2_2 _35895_ (.A(_05165_),
    .B(_05166_),
    .Y(_05167_));
 sky130_as_sc_hs__or2_2 _35897_ (.A(_05150_),
    .B(_05167_),
    .Y(_05169_));
 sky130_as_sc_hs__and2_2 _35898_ (.A(_05168_),
    .B(_05169_),
    .Y(_05170_));
 sky130_as_sc_hs__or2_2 _35900_ (.A(_05149_),
    .B(_05170_),
    .Y(_05172_));
 sky130_as_sc_hs__and2_2 _35901_ (.A(_05171_),
    .B(_05172_),
    .Y(_05173_));
 sky130_as_sc_hs__or2_2 _35904_ (.A(_05173_),
    .B(_05174_),
    .Y(_05176_));
 sky130_as_sc_hs__and2_2 _35905_ (.A(_05175_),
    .B(_05176_),
    .Y(_05177_));
 sky130_as_sc_hs__or2_2 _35907_ (.A(_05148_),
    .B(_05177_),
    .Y(_05179_));
 sky130_as_sc_hs__and2_2 _35908_ (.A(_05178_),
    .B(_05179_),
    .Y(_05180_));
 sky130_as_sc_hs__or2_2 _35910_ (.A(_05127_),
    .B(_05180_),
    .Y(_05182_));
 sky130_as_sc_hs__and2_2 _35911_ (.A(_05181_),
    .B(_05182_),
    .Y(_05183_));
 sky130_as_sc_hs__or2_2 _35913_ (.A(_05126_),
    .B(_05183_),
    .Y(_05185_));
 sky130_as_sc_hs__and2_2 _35914_ (.A(_05184_),
    .B(_05185_),
    .Y(_05186_));
 sky130_as_sc_hs__or2_2 _35920_ (.A(_05189_),
    .B(_05190_),
    .Y(_05192_));
 sky130_as_sc_hs__and2_2 _35921_ (.A(_05191_),
    .B(_05192_),
    .Y(_05193_));
 sky130_as_sc_hs__and2_2 _35922_ (.A(_24808_),
    .B(net424),
    .Y(_05194_));
 sky130_as_sc_hs__or2_2 _35924_ (.A(_05193_),
    .B(_05194_),
    .Y(_05196_));
 sky130_as_sc_hs__and2_2 _35925_ (.A(_05195_),
    .B(_05196_),
    .Y(_05197_));
 sky130_as_sc_hs__and2_2 _35926_ (.A(_24774_),
    .B(net430),
    .Y(_05198_));
 sky130_as_sc_hs__and2_2 _35927_ (.A(_24501_),
    .B(net441),
    .Y(_05199_));
 sky130_as_sc_hs__or2_2 _35928_ (.A(_05198_),
    .B(_05199_),
    .Y(_05200_));
 sky130_as_sc_hs__and2_2 _35930_ (.A(_05200_),
    .B(_05201_),
    .Y(_05202_));
 sky130_as_sc_hs__and2_2 _35931_ (.A(net121),
    .B(_24768_),
    .Y(_05203_));
 sky130_as_sc_hs__or2_2 _35933_ (.A(_05202_),
    .B(_05203_),
    .Y(_05205_));
 sky130_as_sc_hs__and2_2 _35934_ (.A(_05204_),
    .B(_05205_),
    .Y(_05206_));
 sky130_as_sc_hs__or2_2 _35937_ (.A(_05206_),
    .B(_05207_),
    .Y(_05209_));
 sky130_as_sc_hs__and2_2 _35938_ (.A(_05208_),
    .B(_05209_),
    .Y(_05210_));
 sky130_as_sc_hs__or2_2 _35940_ (.A(_05197_),
    .B(_05210_),
    .Y(_05212_));
 sky130_as_sc_hs__and2_2 _35941_ (.A(_05211_),
    .B(_05212_),
    .Y(_05213_));
 sky130_as_sc_hs__and2_2 _35944_ (.A(net479),
    .B(net444),
    .Y(_05216_));
 sky130_as_sc_hs__and2_2 _35945_ (.A(_24229_),
    .B(net435),
    .Y(_05217_));
 sky130_as_sc_hs__or2_2 _35946_ (.A(_05216_),
    .B(_05217_),
    .Y(_05218_));
 sky130_as_sc_hs__and2_2 _35948_ (.A(_05218_),
    .B(_05219_),
    .Y(_05220_));
 sky130_as_sc_hs__and2_2 _35949_ (.A(_24729_),
    .B(net84),
    .Y(_05221_));
 sky130_as_sc_hs__or2_2 _35951_ (.A(_05220_),
    .B(_05221_),
    .Y(_05223_));
 sky130_as_sc_hs__and2_2 _35952_ (.A(_05222_),
    .B(_05223_),
    .Y(_05224_));
 sky130_as_sc_hs__or2_2 _35954_ (.A(_05215_),
    .B(_05224_),
    .Y(_05226_));
 sky130_as_sc_hs__and2_2 _35955_ (.A(_05225_),
    .B(_05226_),
    .Y(_05227_));
 sky130_as_sc_hs__or2_2 _35957_ (.A(_05214_),
    .B(_05227_),
    .Y(_05229_));
 sky130_as_sc_hs__and2_2 _35958_ (.A(_05228_),
    .B(_05229_),
    .Y(_05230_));
 sky130_as_sc_hs__or2_2 _35961_ (.A(_05230_),
    .B(_05231_),
    .Y(_05233_));
 sky130_as_sc_hs__and2_2 _35962_ (.A(_05232_),
    .B(_05233_),
    .Y(_05234_));
 sky130_as_sc_hs__or2_2 _35964_ (.A(_05213_),
    .B(_05234_),
    .Y(_05236_));
 sky130_as_sc_hs__and2_2 _35965_ (.A(_05235_),
    .B(_05236_),
    .Y(_05237_));
 sky130_as_sc_hs__or2_2 _35967_ (.A(_05188_),
    .B(_05237_),
    .Y(_05239_));
 sky130_as_sc_hs__and2_2 _35968_ (.A(_05238_),
    .B(_05239_),
    .Y(_05240_));
 sky130_as_sc_hs__or2_2 _35970_ (.A(_05187_),
    .B(_05240_),
    .Y(_05242_));
 sky130_as_sc_hs__and2_2 _35971_ (.A(_05241_),
    .B(_05242_),
    .Y(_05243_));
 sky130_as_sc_hs__and2_2 _35974_ (.A(net449),
    .B(net439),
    .Y(_05246_));
 sky130_as_sc_hs__and2_2 _35975_ (.A(_23712_),
    .B(net426),
    .Y(_05247_));
 sky130_as_sc_hs__or2_2 _35976_ (.A(_05246_),
    .B(_05247_),
    .Y(_05248_));
 sky130_as_sc_hs__and2_2 _35978_ (.A(_05248_),
    .B(_05249_),
    .Y(_05250_));
 sky130_as_sc_hs__and2_2 _35979_ (.A(net473),
    .B(net451),
    .Y(_05251_));
 sky130_as_sc_hs__or2_2 _35981_ (.A(_05250_),
    .B(_05251_),
    .Y(_05253_));
 sky130_as_sc_hs__and2_2 _35982_ (.A(_05252_),
    .B(_05253_),
    .Y(_05254_));
 sky130_as_sc_hs__and2_2 _35983_ (.A(_23674_),
    .B(_24527_),
    .Y(_05255_));
 sky130_as_sc_hs__and2_2 _35984_ (.A(net480),
    .B(net89),
    .Y(_05256_));
 sky130_as_sc_hs__or2_2 _35985_ (.A(_05255_),
    .B(_05256_),
    .Y(_05257_));
 sky130_as_sc_hs__and2_2 _35987_ (.A(_05257_),
    .B(_05258_),
    .Y(_05259_));
 sky130_as_sc_hs__and2_2 _35988_ (.A(net477),
    .B(net88),
    .Y(_05260_));
 sky130_as_sc_hs__or2_2 _35990_ (.A(_05259_),
    .B(_05260_),
    .Y(_05262_));
 sky130_as_sc_hs__and2_2 _35991_ (.A(_05261_),
    .B(_05262_),
    .Y(_05263_));
 sky130_as_sc_hs__or2_2 _35994_ (.A(_05263_),
    .B(_05264_),
    .Y(_05266_));
 sky130_as_sc_hs__and2_2 _35995_ (.A(_05265_),
    .B(_05266_),
    .Y(_05267_));
 sky130_as_sc_hs__or2_2 _35997_ (.A(_05254_),
    .B(_05267_),
    .Y(_05269_));
 sky130_as_sc_hs__and2_2 _35998_ (.A(_05268_),
    .B(_05269_),
    .Y(_05270_));
 sky130_as_sc_hs__or2_2 _36000_ (.A(_05245_),
    .B(_05270_),
    .Y(_05272_));
 sky130_as_sc_hs__and2_2 _36001_ (.A(_05271_),
    .B(_05272_),
    .Y(_05273_));
 sky130_as_sc_hs__or2_2 _36003_ (.A(_05244_),
    .B(_05273_),
    .Y(_05275_));
 sky130_as_sc_hs__and2_2 _36004_ (.A(_05274_),
    .B(_05275_),
    .Y(_05276_));
 sky130_as_sc_hs__and2_2 _36007_ (.A(net464),
    .B(net446),
    .Y(_05279_));
 sky130_as_sc_hs__and2_2 _36008_ (.A(net462),
    .B(net78),
    .Y(_05280_));
 sky130_as_sc_hs__or2_2 _36009_ (.A(_05279_),
    .B(_05280_),
    .Y(_05281_));
 sky130_as_sc_hs__and2_2 _36011_ (.A(_05281_),
    .B(_05282_),
    .Y(_05283_));
 sky130_as_sc_hs__and2_2 _36012_ (.A(net460),
    .B(net442),
    .Y(_05284_));
 sky130_as_sc_hs__or2_2 _36014_ (.A(_05283_),
    .B(_05284_),
    .Y(_05286_));
 sky130_as_sc_hs__and2_2 _36015_ (.A(_05285_),
    .B(_05286_),
    .Y(_05287_));
 sky130_as_sc_hs__or2_2 _36017_ (.A(_05278_),
    .B(_05287_),
    .Y(_05289_));
 sky130_as_sc_hs__and2_2 _36018_ (.A(_05288_),
    .B(_05289_),
    .Y(_05290_));
 sky130_as_sc_hs__or2_2 _36020_ (.A(_05277_),
    .B(_05290_),
    .Y(_05292_));
 sky130_as_sc_hs__and2_2 _36021_ (.A(_05291_),
    .B(_05292_),
    .Y(_05293_));
 sky130_as_sc_hs__and2_2 _36022_ (.A(net467),
    .B(net454),
    .Y(_05294_));
 sky130_as_sc_hs__and2_2 _36023_ (.A(net469),
    .B(net85),
    .Y(_05295_));
 sky130_as_sc_hs__or2_2 _36024_ (.A(_05294_),
    .B(_05295_),
    .Y(_05296_));
 sky130_as_sc_hs__and2_2 _36026_ (.A(_05296_),
    .B(_05297_),
    .Y(_05298_));
 sky130_as_sc_hs__and2_2 _36027_ (.A(net470),
    .B(net452),
    .Y(_05299_));
 sky130_as_sc_hs__or2_2 _36029_ (.A(_05298_),
    .B(_05299_),
    .Y(_05301_));
 sky130_as_sc_hs__and2_2 _36030_ (.A(_05300_),
    .B(_05301_),
    .Y(_05302_));
 sky130_as_sc_hs__and2_2 _36031_ (.A(_24256_),
    .B(net456),
    .Y(_05303_));
 sky130_as_sc_hs__nand3_2 _36032_ (.A(_24216_),
    .B(_25033_),
    .C(_25034_),
    .Y(_05304_));
 sky130_as_sc_hs__nand3_2 _36033_ (.A(_23598_),
    .B(net458),
    .C(_02549_),
    .Y(_05305_));
 sky130_as_sc_hs__or2_2 _36035_ (.A(_05304_),
    .B(_05305_),
    .Y(_05307_));
 sky130_as_sc_hs__and2_2 _36036_ (.A(_05306_),
    .B(_05307_),
    .Y(_05308_));
 sky130_as_sc_hs__or2_2 _36038_ (.A(_05303_),
    .B(_05308_),
    .Y(_05310_));
 sky130_as_sc_hs__and2_2 _36039_ (.A(_05309_),
    .B(_05310_),
    .Y(_05311_));
 sky130_as_sc_hs__or2_2 _36042_ (.A(_05311_),
    .B(_05312_),
    .Y(_05314_));
 sky130_as_sc_hs__and2_2 _36043_ (.A(_05313_),
    .B(_05314_),
    .Y(_05315_));
 sky130_as_sc_hs__or2_2 _36045_ (.A(_05302_),
    .B(_05315_),
    .Y(_05317_));
 sky130_as_sc_hs__and2_2 _36046_ (.A(_05316_),
    .B(_05317_),
    .Y(_05318_));
 sky130_as_sc_hs__or2_2 _36049_ (.A(_05318_),
    .B(_05319_),
    .Y(_05321_));
 sky130_as_sc_hs__and2_2 _36050_ (.A(_05320_),
    .B(_05321_),
    .Y(_05322_));
 sky130_as_sc_hs__or2_2 _36052_ (.A(_05293_),
    .B(_05322_),
    .Y(_05324_));
 sky130_as_sc_hs__and2_2 _36053_ (.A(_05323_),
    .B(_05324_),
    .Y(_05325_));
 sky130_as_sc_hs__or2_2 _36056_ (.A(_05325_),
    .B(_05326_),
    .Y(_05328_));
 sky130_as_sc_hs__and2_2 _36057_ (.A(_05327_),
    .B(_05328_),
    .Y(_05329_));
 sky130_as_sc_hs__or2_2 _36059_ (.A(_05276_),
    .B(_05329_),
    .Y(_05331_));
 sky130_as_sc_hs__and2_2 _36060_ (.A(_05330_),
    .B(_05331_),
    .Y(_05332_));
 sky130_as_sc_hs__or2_2 _36063_ (.A(_05332_),
    .B(_05333_),
    .Y(_05335_));
 sky130_as_sc_hs__and2_2 _36064_ (.A(_05334_),
    .B(_05335_),
    .Y(_05336_));
 sky130_as_sc_hs__or2_2 _36066_ (.A(_05243_),
    .B(_05336_),
    .Y(_05338_));
 sky130_as_sc_hs__and2_2 _36067_ (.A(_05337_),
    .B(_05338_),
    .Y(_05339_));
 sky130_as_sc_hs__or2_2 _36070_ (.A(_05339_),
    .B(_05340_),
    .Y(_05342_));
 sky130_as_sc_hs__and2_2 _36071_ (.A(_05341_),
    .B(_05342_),
    .Y(_05343_));
 sky130_as_sc_hs__or2_2 _36073_ (.A(_05186_),
    .B(_05343_),
    .Y(_05345_));
 sky130_as_sc_hs__and2_2 _36074_ (.A(_05344_),
    .B(_05345_),
    .Y(_05346_));
 sky130_as_sc_hs__or2_2 _36077_ (.A(_05346_),
    .B(_05347_),
    .Y(_05349_));
 sky130_as_sc_hs__and2_2 _36078_ (.A(_05348_),
    .B(_05349_),
    .Y(_05350_));
 sky130_as_sc_hs__or2_2 _36080_ (.A(_05125_),
    .B(_05350_),
    .Y(_05352_));
 sky130_as_sc_hs__and2_2 _36081_ (.A(_05351_),
    .B(_05352_),
    .Y(_05353_));
 sky130_as_sc_hs__or2_2 _36084_ (.A(_05353_),
    .B(_05354_),
    .Y(_05356_));
 sky130_as_sc_hs__and2_2 _36085_ (.A(_05355_),
    .B(_05356_),
    .Y(_05357_));
 sky130_as_sc_hs__nand3_2 _36086_ (.A(_05124_),
    .B(_05355_),
    .C(_05356_),
    .Y(_05358_));
 sky130_as_sc_hs__or2_2 _36087_ (.A(_05124_),
    .B(_05357_),
    .Y(_05359_));
 sky130_as_sc_hs__and2_2 _36088_ (.A(_05358_),
    .B(_05359_),
    .Y(_05360_));
 sky130_as_sc_hs__nand3_2 _36090_ (.A(_05358_),
    .B(_05359_),
    .C(_05361_),
    .Y(_05362_));
 sky130_as_sc_hs__or2_2 _36091_ (.A(_05360_),
    .B(_05361_),
    .Y(_05363_));
 sky130_as_sc_hs__and2_2 _36092_ (.A(_05362_),
    .B(_05363_),
    .Y(_05364_));
 sky130_as_sc_hs__or2_2 _36094_ (.A(_05123_),
    .B(_05364_),
    .Y(_05366_));
 sky130_as_sc_hs__nand3_2 _36096_ (.A(_04074_),
    .B(_04554_),
    .C(_05093_),
    .Y(_05368_));
 sky130_as_sc_hs__and2_2 _36098_ (.A(_05010_),
    .B(_05369_),
    .Y(_05370_));
 sky130_as_sc_hs__or2_2 _36099_ (.A(_05103_),
    .B(_05370_),
    .Y(_05371_));
 sky130_as_sc_hs__or2_2 _36101_ (.A(_04847_),
    .B(_05371_),
    .Y(_05373_));
 sky130_as_sc_hs__nand3_2 _36103_ (.A(_04074_),
    .B(_04554_),
    .C(_05091_),
    .Y(_05375_));
 sky130_as_sc_hs__or2_2 _36104_ (.A(_04555_),
    .B(_05091_),
    .Y(_05376_));
 sky130_as_sc_hs__or2_2 _36108_ (.A(_05085_),
    .B(_05378_),
    .Y(_05380_));
 sky130_as_sc_hs__and2_2 _36110_ (.A(_05377_),
    .B(_05381_),
    .Y(_05382_));
 sky130_as_sc_hs__or2_2 _36111_ (.A(_04549_),
    .B(_04551_),
    .Y(_05383_));
 sky130_as_sc_hs__or2_2 _36113_ (.A(_04301_),
    .B(_04544_),
    .Y(_05385_));
 sky130_as_sc_hs__or2_2 _36115_ (.A(_04537_),
    .B(_04539_),
    .Y(_05387_));
 sky130_as_sc_hs__or2_2 _36117_ (.A(_04444_),
    .B(_04535_),
    .Y(_05389_));
 sky130_as_sc_hs__or2_2 _36119_ (.A(_04468_),
    .B(_04533_),
    .Y(_05391_));
 sky130_as_sc_hs__or2_2 _36123_ (.A(_04490_),
    .B(_04524_),
    .Y(_05395_));
 sky130_as_sc_hs__and2_2 _36125_ (.A(net116),
    .B(net113),
    .Y(_05397_));
 sky130_as_sc_hs__nor2_2 _36127_ (.A(_05397_),
    .B(_05398_),
    .Y(_05399_));
 sky130_as_sc_hs__and2_2 _36128_ (.A(_04511_),
    .B(_05399_),
    .Y(_05400_));
 sky130_as_sc_hs__nor2b_2 _36129_ (.A(_04517_),
    .Y(_05401_),
    .B(_05400_));
 sky130_as_sc_hs__nand2b_2 _36130_ (.B(_05401_),
    .Y(_05402_),
    .A(_04520_));
 sky130_as_sc_hs__inv_2 _36131_ (.Y(_05403_),
    .A(_05402_));
 sky130_as_sc_hs__and2_2 _36132_ (.A(_04492_),
    .B(_04508_),
    .Y(_05404_));
 sky130_as_sc_hs__or2_2 _36133_ (.A(_04509_),
    .B(_05404_),
    .Y(_05405_));
 sky130_as_sc_hs__and2_2 _36134_ (.A(_05403_),
    .B(_05405_),
    .Y(_05406_));
 sky130_as_sc_hs__and2_2 _36135_ (.A(_05396_),
    .B(_05406_),
    .Y(_05407_));
 sky130_as_sc_hs__and2_2 _36136_ (.A(_05394_),
    .B(_05407_),
    .Y(_05408_));
 sky130_as_sc_hs__and2_2 _36137_ (.A(_05392_),
    .B(_05408_),
    .Y(_05409_));
 sky130_as_sc_hs__and2_2 _36138_ (.A(_05390_),
    .B(_05409_),
    .Y(_05410_));
 sky130_as_sc_hs__inv_2 _36140_ (.Y(_05412_),
    .A(_05411_));
 sky130_as_sc_hs__or2_2 _36142_ (.A(_04541_),
    .B(_05413_),
    .Y(_05414_));
 sky130_as_sc_hs__and2_2 _36144_ (.A(_05414_),
    .B(_05415_),
    .Y(_05416_));
 sky130_as_sc_hs__and2_2 _36145_ (.A(_05412_),
    .B(_05416_),
    .Y(_05417_));
 sky130_as_sc_hs__inv_2 _36147_ (.Y(_05419_),
    .A(_05418_));
 sky130_as_sc_hs__or2_2 _36149_ (.A(_04546_),
    .B(_05420_),
    .Y(_05421_));
 sky130_as_sc_hs__and2_2 _36151_ (.A(_05421_),
    .B(_05422_),
    .Y(_05423_));
 sky130_as_sc_hs__and2_2 _36152_ (.A(_05419_),
    .B(_05423_),
    .Y(_05424_));
 sky130_as_sc_hs__and2_2 _36153_ (.A(_05384_),
    .B(_05424_),
    .Y(_05425_));
 sky130_as_sc_hs__or2_2 _36156_ (.A(_04553_),
    .B(_05426_),
    .Y(_05428_));
 sky130_as_sc_hs__and2_2 _36158_ (.A(_05425_),
    .B(_05429_),
    .Y(_05430_));
 sky130_as_sc_hs__nand3_2 _36159_ (.A(_04074_),
    .B(_04554_),
    .C(_05092_),
    .Y(_05431_));
 sky130_as_sc_hs__nand2b_2 _36160_ (.B(_05431_),
    .Y(_05432_),
    .A(_05096_));
 sky130_as_sc_hs__or2_2 _36162_ (.A(_05070_),
    .B(_05432_),
    .Y(_05434_));
 sky130_as_sc_hs__and2_2 _36164_ (.A(_05430_),
    .B(_05435_),
    .Y(_05436_));
 sky130_as_sc_hs__and2_2 _36165_ (.A(_05382_),
    .B(_05436_),
    .Y(_05437_));
 sky130_as_sc_hs__or2_2 _36168_ (.A(_05048_),
    .B(_05438_),
    .Y(_05440_));
 sky130_as_sc_hs__and2_2 _36170_ (.A(_05437_),
    .B(_05441_),
    .Y(_05442_));
 sky130_as_sc_hs__or2_2 _36172_ (.A(_05009_),
    .B(_05369_),
    .Y(_05444_));
 sky130_as_sc_hs__or2_2 _36176_ (.A(_04942_),
    .B(_05446_),
    .Y(_05448_));
 sky130_as_sc_hs__and2_2 _36178_ (.A(_05445_),
    .B(_05449_),
    .Y(_05450_));
 sky130_as_sc_hs__nand3_2 _36180_ (.A(_05374_),
    .B(_05442_),
    .C(_05450_),
    .Y(_05452_));
 sky130_as_sc_hs__or2_2 _36183_ (.A(_04713_),
    .B(_05453_),
    .Y(_05455_));
 sky130_as_sc_hs__and2_2 _36184_ (.A(_05454_),
    .B(_05455_),
    .Y(_05456_));
 sky130_as_sc_hs__nor2_2 _36185_ (.A(_05452_),
    .B(_05456_),
    .Y(_05457_));
 sky130_as_sc_hs__nand2b_2 _36187_ (.B(_05458_),
    .Y(_05459_),
    .A(_05114_));
 sky130_as_sc_hs__and2_2 _36188_ (.A(_03473_),
    .B(_05459_),
    .Y(_05460_));
 sky130_as_sc_hs__nand3_2 _36189_ (.A(_03147_),
    .B(_03473_),
    .C(_05459_),
    .Y(_05461_));
 sky130_as_sc_hs__or2_2 _36192_ (.A(_02966_),
    .B(_05462_),
    .Y(_05464_));
 sky130_as_sc_hs__or2_2 _36194_ (.A(_03147_),
    .B(_05460_),
    .Y(_05466_));
 sky130_as_sc_hs__nor2_2 _36196_ (.A(_03469_),
    .B(_05108_),
    .Y(_05468_));
 sky130_as_sc_hs__inv_2 _36197_ (.Y(_05469_),
    .A(_05468_));
 sky130_as_sc_hs__or2_2 _36201_ (.A(_03475_),
    .B(_05471_),
    .Y(_05473_));
 sky130_as_sc_hs__and2_2 _36203_ (.A(_05470_),
    .B(_05474_),
    .Y(_05475_));
 sky130_as_sc_hs__and2_2 _36204_ (.A(_05467_),
    .B(_05475_),
    .Y(_05476_));
 sky130_as_sc_hs__nand3_2 _36205_ (.A(_05457_),
    .B(_05465_),
    .C(_05476_),
    .Y(_05477_));
 sky130_as_sc_hs__nand2b_2 _36206_ (.B(_05108_),
    .Y(_05478_),
    .A(_03476_));
 sky130_as_sc_hs__and2_2 _36208_ (.A(_02155_),
    .B(_05479_),
    .Y(_05480_));
 sky130_as_sc_hs__nor2_2 _36210_ (.A(_02155_),
    .B(_05479_),
    .Y(_05482_));
 sky130_as_sc_hs__or2_2 _36211_ (.A(_05480_),
    .B(_05482_),
    .Y(_05483_));
 sky130_as_sc_hs__or2_2 _36214_ (.A(_01966_),
    .B(_05484_),
    .Y(_05486_));
 sky130_as_sc_hs__nor2_2 _36217_ (.A(_05477_),
    .B(_05488_),
    .Y(_05489_));
 sky130_as_sc_hs__or2_2 _36223_ (.A(_02776_),
    .B(_05493_),
    .Y(_05495_));
 sky130_as_sc_hs__or2_2 _36225_ (.A(_02782_),
    .B(_05491_),
    .Y(_05497_));
 sky130_as_sc_hs__inv_2 _36227_ (.Y(_05499_),
    .A(_05498_));
 sky130_as_sc_hs__nand3_2 _36228_ (.A(_05489_),
    .B(_05496_),
    .C(_05498_),
    .Y(_05500_));
 sky130_as_sc_hs__inv_2 _36229_ (.Y(_05501_),
    .A(_05500_));
 sky130_as_sc_hs__and2_2 _36232_ (.A(_05502_),
    .B(_05503_),
    .Y(_05504_));
 sky130_as_sc_hs__or2_2 _36236_ (.A(_05367_),
    .B(_05506_),
    .Y(_05508_));
 sky130_as_sc_hs__nor2_2 _36237_ (.A(net411),
    .B(_19988_),
    .Y(_05509_));
 sky130_as_sc_hs__and2_2 _36238_ (.A(_23604_),
    .B(_05509_),
    .Y(_05510_));
 sky130_as_sc_hs__nand3_2 _36239_ (.A(_05507_),
    .B(_05508_),
    .C(net142),
    .Y(_05511_));
 sky130_as_sc_hs__and2_2 _36240_ (.A(\tholin_riscv.Jimm[13] ),
    .B(_19487_),
    .Y(_05512_));
 sky130_as_sc_hs__and2_2 _36241_ (.A(_19968_),
    .B(_19980_),
    .Y(_05513_));
 sky130_as_sc_hs__and2_2 _36243_ (.A(net334),
    .B(net417),
    .Y(_05515_));
 sky130_as_sc_hs__and2_2 _36244_ (.A(_23598_),
    .B(_05514_),
    .Y(_05516_));
 sky130_as_sc_hs__nor2_2 _36245_ (.A(net149),
    .B(_05516_),
    .Y(_05517_));
 sky130_as_sc_hs__nor2_2 _36246_ (.A(_19474_),
    .B(_19948_),
    .Y(_05518_));
 sky130_as_sc_hs__or2_2 _36247_ (.A(_19474_),
    .B(_19948_),
    .Y(_05519_));
 sky130_as_sc_hs__inv_2 _36251_ (.Y(_05523_),
    .A(_05522_));
 sky130_as_sc_hs__and2_2 _36252_ (.A(_05517_),
    .B(_05523_),
    .Y(_05524_));
 sky130_as_sc_hs__nor2_2 _36253_ (.A(_05517_),
    .B(_05523_),
    .Y(_05525_));
 sky130_as_sc_hs__or2_2 _36254_ (.A(_05524_),
    .B(_05525_),
    .Y(_05526_));
 sky130_as_sc_hs__and2_2 _36255_ (.A(_02381_),
    .B(_05514_),
    .Y(_05527_));
 sky130_as_sc_hs__or2_2 _36256_ (.A(net149),
    .B(_05527_),
    .Y(_05528_));
 sky130_as_sc_hs__inv_2 _36257_ (.Y(_05529_),
    .A(_05528_));
 sky130_as_sc_hs__or2_2 _36259_ (.A(_02474_),
    .B(net126),
    .Y(_05531_));
 sky130_as_sc_hs__and2_2 _36261_ (.A(_05529_),
    .B(_05532_),
    .Y(_05533_));
 sky130_as_sc_hs__and2_2 _36262_ (.A(_05528_),
    .B(_05532_),
    .Y(_05534_));
 sky130_as_sc_hs__nor2_2 _36263_ (.A(_05528_),
    .B(_05532_),
    .Y(_05535_));
 sky130_as_sc_hs__or2_2 _36264_ (.A(_05534_),
    .B(_05535_),
    .Y(_05536_));
 sky130_as_sc_hs__nor2_2 _36265_ (.A(_01723_),
    .B(net416),
    .Y(_05537_));
 sky130_as_sc_hs__or2_2 _36266_ (.A(net149),
    .B(_05537_),
    .Y(_05538_));
 sky130_as_sc_hs__or2_2 _36268_ (.A(_25868_),
    .B(_05518_),
    .Y(_05540_));
 sky130_as_sc_hs__nand2b_2 _36270_ (.B(_05541_),
    .Y(_05542_),
    .A(_05538_));
 sky130_as_sc_hs__or2_2 _36272_ (.A(_05538_),
    .B(_05541_),
    .Y(_05544_));
 sky130_as_sc_hs__nor2_2 _36274_ (.A(_25487_),
    .B(net416),
    .Y(_05546_));
 sky130_as_sc_hs__or2_2 _36275_ (.A(net149),
    .B(_05546_),
    .Y(_05547_));
 sky130_as_sc_hs__nand2b_2 _36279_ (.B(_05550_),
    .Y(_05551_),
    .A(_05547_));
 sky130_as_sc_hs__nand2b_2 _36280_ (.B(_05545_),
    .Y(_05552_),
    .A(_05551_));
 sky130_as_sc_hs__and2_2 _36282_ (.A(_05536_),
    .B(_05553_),
    .Y(_05554_));
 sky130_as_sc_hs__or2_2 _36283_ (.A(_05533_),
    .B(_05554_),
    .Y(_05555_));
 sky130_as_sc_hs__nor2_2 _36285_ (.A(_25027_),
    .B(net416),
    .Y(_05557_));
 sky130_as_sc_hs__or2_2 _36286_ (.A(_05515_),
    .B(_05557_),
    .Y(_05558_));
 sky130_as_sc_hs__nand2b_2 _36290_ (.B(_05561_),
    .Y(_05562_),
    .A(_05558_));
 sky130_as_sc_hs__or2_2 _36292_ (.A(_05558_),
    .B(_05561_),
    .Y(_05564_));
 sky130_as_sc_hs__nor2_2 _36294_ (.A(_24898_),
    .B(net416),
    .Y(_05566_));
 sky130_as_sc_hs__or2_2 _36295_ (.A(net149),
    .B(_05566_),
    .Y(_05567_));
 sky130_as_sc_hs__or2_2 _36297_ (.A(_23397_),
    .B(net126),
    .Y(_05569_));
 sky130_as_sc_hs__nand2b_2 _36299_ (.B(_05570_),
    .Y(_05571_),
    .A(_05567_));
 sky130_as_sc_hs__or2_2 _36301_ (.A(_05567_),
    .B(_05570_),
    .Y(_05573_));
 sky130_as_sc_hs__and2_2 _36303_ (.A(_24337_),
    .B(_05514_),
    .Y(_05575_));
 sky130_as_sc_hs__or2_2 _36304_ (.A(net149),
    .B(_05575_),
    .Y(_05576_));
 sky130_as_sc_hs__or2_2 _36306_ (.A(_23461_),
    .B(net126),
    .Y(_05578_));
 sky130_as_sc_hs__nand2b_2 _36308_ (.B(_05579_),
    .Y(_05580_),
    .A(_05576_));
 sky130_as_sc_hs__or2_2 _36310_ (.A(_05576_),
    .B(_05579_),
    .Y(_05582_));
 sky130_as_sc_hs__nor2_2 _36312_ (.A(_24471_),
    .B(net417),
    .Y(_05584_));
 sky130_as_sc_hs__or2_2 _36313_ (.A(net149),
    .B(_05584_),
    .Y(_05585_));
 sky130_as_sc_hs__or2_2 _36315_ (.A(_23525_),
    .B(net127),
    .Y(_05587_));
 sky130_as_sc_hs__nand2b_2 _36317_ (.B(_05588_),
    .Y(_05589_),
    .A(_05585_));
 sky130_as_sc_hs__nor2_2 _36318_ (.A(_24403_),
    .B(net416),
    .Y(_05590_));
 sky130_as_sc_hs__or2_2 _36319_ (.A(net149),
    .B(_05590_),
    .Y(_05591_));
 sky130_as_sc_hs__nand2b_2 _36323_ (.B(_05594_),
    .Y(_05595_),
    .A(_05591_));
 sky130_as_sc_hs__or2_2 _36325_ (.A(_05591_),
    .B(_05594_),
    .Y(_05597_));
 sky130_as_sc_hs__and2_2 _36326_ (.A(_05596_),
    .B(_05597_),
    .Y(_05598_));
 sky130_as_sc_hs__nor2_2 _36328_ (.A(_24191_),
    .B(net416),
    .Y(_05600_));
 sky130_as_sc_hs__or2_2 _36329_ (.A(_05515_),
    .B(_05600_),
    .Y(_05601_));
 sky130_as_sc_hs__and2_2 _36330_ (.A(\tholin_riscv.PC[22] ),
    .B(net127),
    .Y(_05602_));
 sky130_as_sc_hs__nor2_2 _36331_ (.A(_23077_),
    .B(net126),
    .Y(_05603_));
 sky130_as_sc_hs__or2_2 _36332_ (.A(_05602_),
    .B(_05603_),
    .Y(_05604_));
 sky130_as_sc_hs__nand2b_2 _36333_ (.B(_05604_),
    .Y(_05605_),
    .A(_05601_));
 sky130_as_sc_hs__or2_2 _36335_ (.A(_05601_),
    .B(_05604_),
    .Y(_05607_));
 sky130_as_sc_hs__and2_2 _36336_ (.A(_05606_),
    .B(_05607_),
    .Y(_05608_));
 sky130_as_sc_hs__nor2_2 _36338_ (.A(_24116_),
    .B(net417),
    .Y(_05610_));
 sky130_as_sc_hs__or2_2 _36339_ (.A(_05515_),
    .B(_05610_),
    .Y(_05611_));
 sky130_as_sc_hs__and2_2 _36340_ (.A(\tholin_riscv.PC[21] ),
    .B(net126),
    .Y(_05612_));
 sky130_as_sc_hs__nor2_2 _36341_ (.A(_23204_),
    .B(net126),
    .Y(_05613_));
 sky130_as_sc_hs__or2_2 _36342_ (.A(_05612_),
    .B(_05613_),
    .Y(_05614_));
 sky130_as_sc_hs__nand2b_2 _36343_ (.B(_05614_),
    .Y(_05615_),
    .A(_05611_));
 sky130_as_sc_hs__or2_2 _36345_ (.A(_05611_),
    .B(_05614_),
    .Y(_05617_));
 sky130_as_sc_hs__and2_2 _36346_ (.A(_05616_),
    .B(_05617_),
    .Y(_05618_));
 sky130_as_sc_hs__nor2_2 _36348_ (.A(_23775_),
    .B(net417),
    .Y(_05620_));
 sky130_as_sc_hs__or2_2 _36349_ (.A(_05515_),
    .B(_05620_),
    .Y(_05621_));
 sky130_as_sc_hs__and2_2 _36350_ (.A(\tholin_riscv.PC[20] ),
    .B(net126),
    .Y(_05622_));
 sky130_as_sc_hs__nor2_2 _36351_ (.A(_23268_),
    .B(net126),
    .Y(_05623_));
 sky130_as_sc_hs__or2_2 _36352_ (.A(_05622_),
    .B(_05623_),
    .Y(_05624_));
 sky130_as_sc_hs__nand2b_2 _36353_ (.B(_05624_),
    .Y(_05625_),
    .A(_05621_));
 sky130_as_sc_hs__or2_2 _36355_ (.A(_05621_),
    .B(_05624_),
    .Y(_05627_));
 sky130_as_sc_hs__and2_2 _36356_ (.A(_05626_),
    .B(_05627_),
    .Y(_05628_));
 sky130_as_sc_hs__nor2_2 _36358_ (.A(_23839_),
    .B(net416),
    .Y(_05630_));
 sky130_as_sc_hs__or2_2 _36359_ (.A(_05515_),
    .B(_05630_),
    .Y(_05631_));
 sky130_as_sc_hs__and2_2 _36360_ (.A(\tholin_riscv.PC[19] ),
    .B(net127),
    .Y(_05632_));
 sky130_as_sc_hs__nor2_2 _36361_ (.A(_21786_),
    .B(net126),
    .Y(_05633_));
 sky130_as_sc_hs__or2_2 _36362_ (.A(_05632_),
    .B(_05633_),
    .Y(_05634_));
 sky130_as_sc_hs__nand2b_2 _36363_ (.B(_05634_),
    .Y(_05635_),
    .A(_05631_));
 sky130_as_sc_hs__or2_2 _36365_ (.A(_05631_),
    .B(_05634_),
    .Y(_05637_));
 sky130_as_sc_hs__and2_2 _36366_ (.A(_05636_),
    .B(_05637_),
    .Y(_05638_));
 sky130_as_sc_hs__nor2_2 _36368_ (.A(_23902_),
    .B(net416),
    .Y(_05640_));
 sky130_as_sc_hs__or2_2 _36369_ (.A(net149),
    .B(_05640_),
    .Y(_05641_));
 sky130_as_sc_hs__and2_2 _36370_ (.A(\tholin_riscv.PC[18] ),
    .B(net126),
    .Y(_05642_));
 sky130_as_sc_hs__nor2_2 _36371_ (.A(_23011_),
    .B(net126),
    .Y(_05643_));
 sky130_as_sc_hs__or2_2 _36372_ (.A(_05642_),
    .B(_05643_),
    .Y(_05644_));
 sky130_as_sc_hs__nand2b_2 _36373_ (.B(_05644_),
    .Y(_05645_),
    .A(_05641_));
 sky130_as_sc_hs__or2_2 _36375_ (.A(_05641_),
    .B(_05644_),
    .Y(_05647_));
 sky130_as_sc_hs__and2_2 _36376_ (.A(_05646_),
    .B(_05647_),
    .Y(_05648_));
 sky130_as_sc_hs__nor2_2 _36378_ (.A(_23966_),
    .B(net416),
    .Y(_05650_));
 sky130_as_sc_hs__or2_2 _36379_ (.A(net149),
    .B(_05650_),
    .Y(_05651_));
 sky130_as_sc_hs__and2_2 _36380_ (.A(\tholin_riscv.PC[17] ),
    .B(net126),
    .Y(_05652_));
 sky130_as_sc_hs__nor2_2 _36381_ (.A(_21850_),
    .B(net126),
    .Y(_05653_));
 sky130_as_sc_hs__or2_2 _36382_ (.A(_05652_),
    .B(_05653_),
    .Y(_05654_));
 sky130_as_sc_hs__nand2b_2 _36383_ (.B(_05654_),
    .Y(_05655_),
    .A(_05651_));
 sky130_as_sc_hs__or2_2 _36385_ (.A(_05651_),
    .B(_05654_),
    .Y(_05657_));
 sky130_as_sc_hs__nor2_2 _36387_ (.A(_24037_),
    .B(net416),
    .Y(_05659_));
 sky130_as_sc_hs__or2_2 _36388_ (.A(net149),
    .B(_05659_),
    .Y(_05660_));
 sky130_as_sc_hs__and2_2 _36389_ (.A(\tholin_riscv.PC[16] ),
    .B(net127),
    .Y(_05661_));
 sky130_as_sc_hs__nor2_2 _36390_ (.A(_22945_),
    .B(net126),
    .Y(_05662_));
 sky130_as_sc_hs__or2_2 _36391_ (.A(_05661_),
    .B(_05662_),
    .Y(_05663_));
 sky130_as_sc_hs__or2_2 _36393_ (.A(_05660_),
    .B(_05663_),
    .Y(_05665_));
 sky130_as_sc_hs__and2_2 _36395_ (.A(_20707_),
    .B(_05514_),
    .Y(_05667_));
 sky130_as_sc_hs__or2_2 _36396_ (.A(net149),
    .B(_05667_),
    .Y(_05668_));
 sky130_as_sc_hs__inv_2 _36397_ (.Y(_05669_),
    .A(_05668_));
 sky130_as_sc_hs__or2_2 _36399_ (.A(_22750_),
    .B(net127),
    .Y(_05671_));
 sky130_as_sc_hs__or2_2 _36403_ (.A(_05668_),
    .B(_05672_),
    .Y(_05675_));
 sky130_as_sc_hs__and2_2 _36405_ (.A(_20622_),
    .B(_05514_),
    .Y(_05677_));
 sky130_as_sc_hs__or2_2 _36406_ (.A(net149),
    .B(_05677_),
    .Y(_05678_));
 sky130_as_sc_hs__inv_2 _36407_ (.Y(_05679_),
    .A(_05678_));
 sky130_as_sc_hs__or2_2 _36413_ (.A(_05678_),
    .B(_05682_),
    .Y(_05685_));
 sky130_as_sc_hs__nor2_2 _36415_ (.A(_20535_),
    .B(net416),
    .Y(_05687_));
 sky130_as_sc_hs__or2_2 _36416_ (.A(net149),
    .B(_05687_),
    .Y(_05688_));
 sky130_as_sc_hs__inv_2 _36417_ (.Y(_05689_),
    .A(_05688_));
 sky130_as_sc_hs__or2_2 _36419_ (.A(_22815_),
    .B(_05518_),
    .Y(_05691_));
 sky130_as_sc_hs__or2_2 _36423_ (.A(_05688_),
    .B(_05692_),
    .Y(_05695_));
 sky130_as_sc_hs__nor2_2 _36425_ (.A(_20449_),
    .B(net416),
    .Y(_05697_));
 sky130_as_sc_hs__or2_2 _36426_ (.A(net149),
    .B(_05697_),
    .Y(_05698_));
 sky130_as_sc_hs__inv_2 _36427_ (.Y(_05699_),
    .A(_05698_));
 sky130_as_sc_hs__or2_2 _36429_ (.A(_22879_),
    .B(net126),
    .Y(_05701_));
 sky130_as_sc_hs__or2_2 _36433_ (.A(_05698_),
    .B(_05702_),
    .Y(_05705_));
 sky130_as_sc_hs__nor2_2 _36435_ (.A(_20363_),
    .B(net416),
    .Y(_05707_));
 sky130_as_sc_hs__or2_2 _36436_ (.A(net149),
    .B(_05707_),
    .Y(_05708_));
 sky130_as_sc_hs__nand2b_2 _36440_ (.B(_05711_),
    .Y(_05712_),
    .A(_05708_));
 sky130_as_sc_hs__or2_2 _36442_ (.A(_05708_),
    .B(_05711_),
    .Y(_05714_));
 sky130_as_sc_hs__and2_2 _36447_ (.A(\tholin_riscv.Bimm[10] ),
    .B(net417),
    .Y(_05719_));
 sky130_as_sc_hs__nor2_2 _36448_ (.A(_20277_),
    .B(net416),
    .Y(_05720_));
 sky130_as_sc_hs__nor2_2 _36449_ (.A(_05719_),
    .B(_05720_),
    .Y(_05721_));
 sky130_as_sc_hs__inv_2 _36450_ (.Y(_05722_),
    .A(_05721_));
 sky130_as_sc_hs__or2_2 _36453_ (.A(_05718_),
    .B(_05722_),
    .Y(_05725_));
 sky130_as_sc_hs__and2_2 _36458_ (.A(\tholin_riscv.Bimm[9] ),
    .B(net417),
    .Y(_05730_));
 sky130_as_sc_hs__nor2_2 _36459_ (.A(_20191_),
    .B(net416),
    .Y(_05731_));
 sky130_as_sc_hs__nor2_2 _36460_ (.A(_05730_),
    .B(_05731_),
    .Y(_05732_));
 sky130_as_sc_hs__inv_2 _36461_ (.Y(_05733_),
    .A(_05732_));
 sky130_as_sc_hs__or2_2 _36464_ (.A(_05729_),
    .B(_05733_),
    .Y(_05736_));
 sky130_as_sc_hs__and2_2 _36465_ (.A(_05735_),
    .B(_05736_),
    .Y(_05737_));
 sky130_as_sc_hs__inv_2 _36466_ (.Y(_05738_),
    .A(_05737_));
 sky130_as_sc_hs__and2_2 _36470_ (.A(\tholin_riscv.Bimm[8] ),
    .B(net417),
    .Y(_05742_));
 sky130_as_sc_hs__nor2_2 _36471_ (.A(_20105_),
    .B(net416),
    .Y(_05743_));
 sky130_as_sc_hs__nor2_2 _36472_ (.A(_05742_),
    .B(_05743_),
    .Y(_05744_));
 sky130_as_sc_hs__inv_2 _36473_ (.Y(_05745_),
    .A(_05744_));
 sky130_as_sc_hs__and2_2 _36475_ (.A(\tholin_riscv.PC[7] ),
    .B(net127),
    .Y(_05747_));
 sky130_as_sc_hs__and2_2 _36476_ (.A(_22301_),
    .B(_05519_),
    .Y(_05748_));
 sky130_as_sc_hs__or2_2 _36477_ (.A(_05747_),
    .B(_05748_),
    .Y(_05749_));
 sky130_as_sc_hs__and2_2 _36478_ (.A(\tholin_riscv.Bimm[7] ),
    .B(net417),
    .Y(_05750_));
 sky130_as_sc_hs__nor2_2 _36479_ (.A(_21534_),
    .B(net417),
    .Y(_05751_));
 sky130_as_sc_hs__nor2_2 _36480_ (.A(_05750_),
    .B(_05751_),
    .Y(_05752_));
 sky130_as_sc_hs__inv_2 _36481_ (.Y(_05753_),
    .A(_05752_));
 sky130_as_sc_hs__or2_2 _36484_ (.A(_05749_),
    .B(_05753_),
    .Y(_05756_));
 sky130_as_sc_hs__inv_2 _36489_ (.Y(_05761_),
    .A(_05760_));
 sky130_as_sc_hs__and2_2 _36492_ (.A(_05762_),
    .B(_05763_),
    .Y(_05764_));
 sky130_as_sc_hs__or2_2 _36494_ (.A(_05761_),
    .B(_05764_),
    .Y(_05766_));
 sky130_as_sc_hs__inv_2 _36500_ (.Y(_05772_),
    .A(_05771_));
 sky130_as_sc_hs__and2_2 _36503_ (.A(_05773_),
    .B(_05774_),
    .Y(_05775_));
 sky130_as_sc_hs__or2_2 _36505_ (.A(_05772_),
    .B(_05775_),
    .Y(_05777_));
 sky130_as_sc_hs__and2_2 _36507_ (.A(_05777_),
    .B(_05778_),
    .Y(_05779_));
 sky130_as_sc_hs__inv_2 _36508_ (.Y(_05780_),
    .A(_05779_));
 sky130_as_sc_hs__or2_2 _36517_ (.A(\tholin_riscv.Bimm[4] ),
    .B(_05784_),
    .Y(_05789_));
 sky130_as_sc_hs__and2_2 _36518_ (.A(_05788_),
    .B(_05789_),
    .Y(_05790_));
 sky130_as_sc_hs__inv_2 _36519_ (.Y(_05791_),
    .A(_05790_));
 sky130_as_sc_hs__nor2_2 _36521_ (.A(_05783_),
    .B(_05790_),
    .Y(_05793_));
 sky130_as_sc_hs__inv_2 _36522_ (.Y(_05794_),
    .A(_05793_));
 sky130_as_sc_hs__and2_2 _36524_ (.A(\tholin_riscv.PC[3] ),
    .B(net127),
    .Y(_05796_));
 sky130_as_sc_hs__and2_2 _36525_ (.A(_21977_),
    .B(_05519_),
    .Y(_05797_));
 sky130_as_sc_hs__or2_2 _36526_ (.A(_05796_),
    .B(_05797_),
    .Y(_05798_));
 sky130_as_sc_hs__or2_2 _36531_ (.A(\tholin_riscv.Bimm[3] ),
    .B(_05784_),
    .Y(_05803_));
 sky130_as_sc_hs__and2_2 _36532_ (.A(_05802_),
    .B(_05803_),
    .Y(_05804_));
 sky130_as_sc_hs__inv_2 _36533_ (.Y(_05805_),
    .A(_05804_));
 sky130_as_sc_hs__nor2_2 _36536_ (.A(_05798_),
    .B(_05804_),
    .Y(_05808_));
 sky130_as_sc_hs__inv_2 _36537_ (.Y(_05809_),
    .A(_05808_));
 sky130_as_sc_hs__and2_2 _36542_ (.A(_21037_),
    .B(_05514_),
    .Y(_05814_));
 sky130_as_sc_hs__nor2_2 _36543_ (.A(\tholin_riscv.Iimm[2] ),
    .B(_05514_),
    .Y(_05815_));
 sky130_as_sc_hs__or2_2 _36544_ (.A(_05814_),
    .B(_05815_),
    .Y(_05816_));
 sky130_as_sc_hs__or2_2 _36546_ (.A(\tholin_riscv.Bimm[2] ),
    .B(_05784_),
    .Y(_05818_));
 sky130_as_sc_hs__and2_2 _36547_ (.A(_05817_),
    .B(_05818_),
    .Y(_05819_));
 sky130_as_sc_hs__inv_2 _36548_ (.Y(_05820_),
    .A(_05819_));
 sky130_as_sc_hs__and2_2 _36550_ (.A(_05813_),
    .B(_05819_),
    .Y(_05822_));
 sky130_as_sc_hs__nor2_2 _36551_ (.A(_05813_),
    .B(_05819_),
    .Y(_05823_));
 sky130_as_sc_hs__or2_2 _36552_ (.A(_05822_),
    .B(_05823_),
    .Y(_05824_));
 sky130_as_sc_hs__and2_2 _36553_ (.A(\tholin_riscv.PC[1] ),
    .B(net127),
    .Y(_05825_));
 sky130_as_sc_hs__nor2_2 _36554_ (.A(_22104_),
    .B(net126),
    .Y(_05826_));
 sky130_as_sc_hs__or2_2 _36555_ (.A(_05825_),
    .B(_05826_),
    .Y(_05827_));
 sky130_as_sc_hs__nand3_2 _36558_ (.A(_05784_),
    .B(_05828_),
    .C(_05829_),
    .Y(_05830_));
 sky130_as_sc_hs__nand3_2 _36559_ (.A(\tholin_riscv.instr[5] ),
    .B(\tholin_riscv.Bimm[1] ),
    .C(_19971_),
    .Y(_05831_));
 sky130_as_sc_hs__nand3_2 _36561_ (.A(_05827_),
    .B(_05830_),
    .C(_05831_),
    .Y(_05833_));
 sky130_as_sc_hs__and2_2 _36562_ (.A(_05827_),
    .B(_05832_),
    .Y(_05834_));
 sky130_as_sc_hs__nor2_2 _36563_ (.A(_05827_),
    .B(_05832_),
    .Y(_05835_));
 sky130_as_sc_hs__or2_2 _36564_ (.A(_05834_),
    .B(_05835_),
    .Y(_05836_));
 sky130_as_sc_hs__and2_2 _36565_ (.A(\tholin_riscv.PC[0] ),
    .B(net127),
    .Y(_05837_));
 sky130_as_sc_hs__and2_2 _36566_ (.A(net113),
    .B(_05519_),
    .Y(_05838_));
 sky130_as_sc_hs__nor2_2 _36567_ (.A(_05837_),
    .B(_05838_),
    .Y(_05839_));
 sky130_as_sc_hs__or2_2 _36568_ (.A(_05837_),
    .B(_05838_),
    .Y(_05840_));
 sky130_as_sc_hs__and2_2 _36569_ (.A(_20826_),
    .B(_05514_),
    .Y(_05841_));
 sky130_as_sc_hs__nor2_2 _36570_ (.A(\tholin_riscv.Iimm[0] ),
    .B(_05514_),
    .Y(_05842_));
 sky130_as_sc_hs__or2_2 _36571_ (.A(_05841_),
    .B(_05842_),
    .Y(_05843_));
 sky130_as_sc_hs__or2_2 _36573_ (.A(\tholin_riscv.Bimm[11] ),
    .B(_05784_),
    .Y(_05845_));
 sky130_as_sc_hs__and2_2 _36574_ (.A(_05844_),
    .B(_05845_),
    .Y(_05846_));
 sky130_as_sc_hs__and2_2 _36584_ (.A(_05854_),
    .B(_05855_),
    .Y(_05856_));
 sky130_as_sc_hs__or2_2 _36585_ (.A(_05779_),
    .B(_05856_),
    .Y(_05857_));
 sky130_as_sc_hs__or2_2 _36592_ (.A(_05741_),
    .B(_05745_),
    .Y(_05864_));
 sky130_as_sc_hs__and2_2 _36595_ (.A(_05746_),
    .B(_05866_),
    .Y(_05867_));
 sky130_as_sc_hs__or2_2 _36596_ (.A(_05737_),
    .B(_05867_),
    .Y(_05868_));
 sky130_as_sc_hs__nand2b_2 _36611_ (.B(_05663_),
    .Y(_05883_),
    .A(_05660_));
 sky130_as_sc_hs__or2_2 _36628_ (.A(_05585_),
    .B(_05588_),
    .Y(_05900_));
 sky130_as_sc_hs__or2_2 _36639_ (.A(_05547_),
    .B(_05550_),
    .Y(_05911_));
 sky130_as_sc_hs__and2_2 _36641_ (.A(_05545_),
    .B(_05912_),
    .Y(_05913_));
 sky130_as_sc_hs__nand3_2 _36642_ (.A(_05526_),
    .B(_05536_),
    .C(_05913_),
    .Y(_05914_));
 sky130_as_sc_hs__inv_2 _36643_ (.Y(_05915_),
    .A(_05914_));
 sky130_as_sc_hs__nand3_2 _36645_ (.A(_05526_),
    .B(_05556_),
    .C(_05916_),
    .Y(_05917_));
 sky130_as_sc_hs__nand3_2 _36649_ (.A(_05556_),
    .B(_05916_),
    .C(_05918_),
    .Y(_05921_));
 sky130_as_sc_hs__or2_2 _36650_ (.A(_21657_),
    .B(_05921_),
    .Y(_05922_));
 sky130_as_sc_hs__nor2_2 _36652_ (.A(net411),
    .B(_19987_),
    .Y(_05924_));
 sky130_as_sc_hs__and2_2 _36654_ (.A(_19988_),
    .B(_23601_),
    .Y(_05926_));
 sky130_as_sc_hs__inv_2 _36658_ (.Y(_05930_),
    .A(_05929_));
 sky130_as_sc_hs__and2_2 _36659_ (.A(\tholin_riscv.Bimm[10] ),
    .B(_05522_),
    .Y(_05931_));
 sky130_as_sc_hs__inv_2 _36664_ (.Y(_05936_),
    .A(_05935_));
 sky130_as_sc_hs__and2_2 _36666_ (.A(_19979_),
    .B(_21036_),
    .Y(_05938_));
 sky130_as_sc_hs__and2_2 _36667_ (.A(\tholin_riscv.Iimm[2] ),
    .B(_19980_),
    .Y(_05939_));
 sky130_as_sc_hs__or2_2 _36668_ (.A(_05938_),
    .B(_05939_),
    .Y(_05940_));
 sky130_as_sc_hs__nor2_2 _36669_ (.A(_05938_),
    .B(_05939_),
    .Y(_05941_));
 sky130_as_sc_hs__and2_2 _36671_ (.A(_19979_),
    .B(_20931_),
    .Y(_05943_));
 sky130_as_sc_hs__and2_2 _36672_ (.A(\tholin_riscv.Iimm[1] ),
    .B(_19980_),
    .Y(_05944_));
 sky130_as_sc_hs__or2_2 _36673_ (.A(_05943_),
    .B(_05944_),
    .Y(_05945_));
 sky130_as_sc_hs__nor2_2 _36674_ (.A(_05943_),
    .B(_05944_),
    .Y(_05946_));
 sky130_as_sc_hs__and2_2 _36675_ (.A(_05931_),
    .B(net82),
    .Y(_05947_));
 sky130_as_sc_hs__and2_2 _36676_ (.A(_19979_),
    .B(net116),
    .Y(_05948_));
 sky130_as_sc_hs__and2_2 _36677_ (.A(\tholin_riscv.Iimm[0] ),
    .B(_19980_),
    .Y(_05949_));
 sky130_as_sc_hs__or2_2 _36678_ (.A(_05948_),
    .B(_05949_),
    .Y(_05950_));
 sky130_as_sc_hs__nor2_2 _36679_ (.A(_05948_),
    .B(_05949_),
    .Y(_05951_));
 sky130_as_sc_hs__and2_2 _36686_ (.A(_05946_),
    .B(_05957_),
    .Y(_05958_));
 sky130_as_sc_hs__nor2_2 _36687_ (.A(_05947_),
    .B(_05958_),
    .Y(_05959_));
 sky130_as_sc_hs__or2_2 _36688_ (.A(_05940_),
    .B(_05959_),
    .Y(_05960_));
 sky130_as_sc_hs__and2_2 _36694_ (.A(_05926_),
    .B(_05965_),
    .Y(_05966_));
 sky130_as_sc_hs__and2_2 _36695_ (.A(net411),
    .B(_19988_),
    .Y(_05967_));
 sky130_as_sc_hs__and2_2 _36696_ (.A(_23599_),
    .B(_05967_),
    .Y(_05968_));
 sky130_as_sc_hs__or2_2 _36701_ (.A(_23602_),
    .B(_05522_),
    .Y(_05973_));
 sky130_as_sc_hs__nand3_2 _36703_ (.A(_05951_),
    .B(_05973_),
    .C(_05974_),
    .Y(_05975_));
 sky130_as_sc_hs__nand3_2 _36704_ (.A(_05946_),
    .B(_05972_),
    .C(_05975_),
    .Y(_05976_));
 sky130_as_sc_hs__and2_2 _36713_ (.A(_05980_),
    .B(_05984_),
    .Y(_05985_));
 sky130_as_sc_hs__and2_2 _36723_ (.A(_05990_),
    .B(_05994_),
    .Y(_05995_));
 sky130_as_sc_hs__or2_2 _36734_ (.A(net82),
    .B(_06005_),
    .Y(_06006_));
 sky130_as_sc_hs__and2_2 _36735_ (.A(_05996_),
    .B(_06006_),
    .Y(_06007_));
 sky130_as_sc_hs__nand3_2 _36737_ (.A(_05941_),
    .B(_05976_),
    .C(_05986_),
    .Y(_06009_));
 sky130_as_sc_hs__nand3_2 _36738_ (.A(_05935_),
    .B(_06008_),
    .C(_06009_),
    .Y(_06010_));
 sky130_as_sc_hs__and2_2 _36747_ (.A(_06014_),
    .B(_06018_),
    .Y(_06019_));
 sky130_as_sc_hs__or2_2 _36758_ (.A(net82),
    .B(_06029_),
    .Y(_06030_));
 sky130_as_sc_hs__or2_2 _36760_ (.A(_05940_),
    .B(_06031_),
    .Y(_06032_));
 sky130_as_sc_hs__and2_2 _36764_ (.A(_05950_),
    .B(_06035_),
    .Y(_06036_));
 sky130_as_sc_hs__and2_2 _36768_ (.A(_05951_),
    .B(_06039_),
    .Y(_06040_));
 sky130_as_sc_hs__or2_2 _36769_ (.A(_06036_),
    .B(_06040_),
    .Y(_06041_));
 sky130_as_sc_hs__and2_2 _36778_ (.A(_06045_),
    .B(_06049_),
    .Y(_06050_));
 sky130_as_sc_hs__or2_2 _36779_ (.A(net82),
    .B(_06050_),
    .Y(_06051_));
 sky130_as_sc_hs__and2_2 _36783_ (.A(_06032_),
    .B(_06054_),
    .Y(_06055_));
 sky130_as_sc_hs__and2_2 _36795_ (.A(_06062_),
    .B(_06066_),
    .Y(_06067_));
 sky130_as_sc_hs__or2_2 _36806_ (.A(net82),
    .B(_06077_),
    .Y(_06078_));
 sky130_as_sc_hs__and2_2 _36807_ (.A(_06068_),
    .B(_06078_),
    .Y(_06079_));
 sky130_as_sc_hs__and2_2 _36817_ (.A(_06084_),
    .B(_06088_),
    .Y(_06089_));
 sky130_as_sc_hs__and2_2 _36827_ (.A(_06094_),
    .B(_06098_),
    .Y(_06099_));
 sky130_as_sc_hs__and2_2 _36829_ (.A(_06090_),
    .B(_06100_),
    .Y(_06101_));
 sky130_as_sc_hs__and2_2 _36841_ (.A(_06108_),
    .B(_06112_),
    .Y(_06113_));
 sky130_as_sc_hs__and2_2 _36851_ (.A(_06118_),
    .B(_06122_),
    .Y(_06123_));
 sky130_as_sc_hs__and2_2 _36853_ (.A(_06114_),
    .B(_06124_),
    .Y(_06125_));
 sky130_as_sc_hs__and2_2 _36855_ (.A(_05950_),
    .B(_05954_),
    .Y(_06127_));
 sky130_as_sc_hs__and2_2 _36859_ (.A(_05951_),
    .B(_06130_),
    .Y(_06131_));
 sky130_as_sc_hs__or2_2 _36860_ (.A(_06127_),
    .B(_06131_),
    .Y(_06132_));
 sky130_as_sc_hs__and2_2 _36869_ (.A(_06136_),
    .B(_06140_),
    .Y(_06141_));
 sky130_as_sc_hs__or2_2 _36870_ (.A(net82),
    .B(_06141_),
    .Y(_06142_));
 sky130_as_sc_hs__or2_2 _36877_ (.A(_05929_),
    .B(_06148_),
    .Y(_06149_));
 sky130_as_sc_hs__and2_2 _36878_ (.A(_06058_),
    .B(_06149_),
    .Y(_06150_));
 sky130_as_sc_hs__and2_2 _36880_ (.A(_05840_),
    .B(_05846_),
    .Y(_06152_));
 sky130_as_sc_hs__nor2_2 _36882_ (.A(_05840_),
    .B(_05846_),
    .Y(_06154_));
 sky130_as_sc_hs__nor2_2 _36883_ (.A(_06152_),
    .B(_06154_),
    .Y(_06155_));
 sky130_as_sc_hs__nand3_2 _36884_ (.A(_19988_),
    .B(_23603_),
    .C(_06155_),
    .Y(_06156_));
 sky130_as_sc_hs__and2_2 _36885_ (.A(_05512_),
    .B(_05967_),
    .Y(_06157_));
 sky130_as_sc_hs__nor2_2 _36887_ (.A(_06154_),
    .B(_06158_),
    .Y(_06159_));
 sky130_as_sc_hs__and2_2 _36888_ (.A(_21656_),
    .B(_05967_),
    .Y(_06160_));
 sky130_as_sc_hs__and2_2 _36891_ (.A(_23603_),
    .B(_05509_),
    .Y(_06163_));
 sky130_as_sc_hs__and2_2 _36893_ (.A(net411),
    .B(_19987_),
    .Y(_06165_));
 sky130_as_sc_hs__or2_2 _36894_ (.A(\tholin_riscv.Jimm[13] ),
    .B(\tholin_riscv.div_res[0] ),
    .Y(_06166_));
 sky130_as_sc_hs__nand3_2 _36896_ (.A(_06165_),
    .B(_06166_),
    .C(_06167_),
    .Y(_06168_));
 sky130_as_sc_hs__nand3_2 _36897_ (.A(net413),
    .B(_06164_),
    .C(_06168_),
    .Y(_06169_));
 sky130_as_sc_hs__nor2_2 _36898_ (.A(_06159_),
    .B(_06169_),
    .Y(_06170_));
 sky130_as_sc_hs__nand3_2 _36899_ (.A(_06156_),
    .B(_06162_),
    .C(_06170_),
    .Y(_06171_));
 sky130_as_sc_hs__nor2_2 _36900_ (.A(_05966_),
    .B(_06171_),
    .Y(_06172_));
 sky130_as_sc_hs__and2_2 _36901_ (.A(_06151_),
    .B(_06172_),
    .Y(_06173_));
 sky130_as_sc_hs__nand3_2 _36902_ (.A(_05511_),
    .B(_05925_),
    .C(_06173_),
    .Y(_06174_));
 sky130_as_sc_hs__inv_2 _36906_ (.Y(_06178_),
    .A(_06177_));
 sky130_as_sc_hs__or2_2 _36908_ (.A(net735),
    .B(_21586_),
    .Y(_06180_));
 sky130_as_sc_hs__and2_2 _36909_ (.A(_06179_),
    .B(net736),
    .Y(_00021_));
 sky130_as_sc_hs__and2_2 _36915_ (.A(_23636_),
    .B(net121),
    .Y(_06186_));
 sky130_as_sc_hs__and2_2 _36916_ (.A(_23712_),
    .B(net422),
    .Y(_06187_));
 sky130_as_sc_hs__or2_2 _36917_ (.A(_06186_),
    .B(_06187_),
    .Y(_06188_));
 sky130_as_sc_hs__and2_2 _36919_ (.A(_06188_),
    .B(_06189_),
    .Y(_06190_));
 sky130_as_sc_hs__and2_2 _36920_ (.A(net482),
    .B(net84),
    .Y(_06191_));
 sky130_as_sc_hs__or2_2 _36922_ (.A(_06190_),
    .B(_06191_),
    .Y(_06193_));
 sky130_as_sc_hs__and2_2 _36923_ (.A(_06192_),
    .B(_06193_),
    .Y(_06194_));
 sky130_as_sc_hs__or2_2 _36926_ (.A(_06194_),
    .B(_06195_),
    .Y(_06197_));
 sky130_as_sc_hs__or2_2 _36928_ (.A(_05138_),
    .B(_06198_),
    .Y(_06199_));
 sky130_as_sc_hs__and2_2 _36930_ (.A(_06199_),
    .B(_06200_),
    .Y(_06201_));
 sky130_as_sc_hs__and2_2 _36931_ (.A(_23702_),
    .B(net430),
    .Y(_06202_));
 sky130_as_sc_hs__or2_2 _36933_ (.A(_06201_),
    .B(_06202_),
    .Y(_06204_));
 sky130_as_sc_hs__and2_2 _36934_ (.A(_06203_),
    .B(_06204_),
    .Y(_06205_));
 sky130_as_sc_hs__and2_2 _36939_ (.A(_25211_),
    .B(net75),
    .Y(_06210_));
 sky130_as_sc_hs__and2_2 _36940_ (.A(_24053_),
    .B(net129),
    .Y(_06211_));
 sky130_as_sc_hs__or2_2 _36942_ (.A(_06210_),
    .B(_06211_),
    .Y(_06213_));
 sky130_as_sc_hs__and2_2 _36943_ (.A(_06212_),
    .B(_06213_),
    .Y(_06214_));
 sky130_as_sc_hs__or2_2 _36945_ (.A(_06209_),
    .B(_06214_),
    .Y(_06216_));
 sky130_as_sc_hs__and2_2 _36946_ (.A(_06215_),
    .B(_06216_),
    .Y(_06217_));
 sky130_as_sc_hs__or2_2 _36948_ (.A(_06208_),
    .B(_06217_),
    .Y(_06219_));
 sky130_as_sc_hs__and2_2 _36949_ (.A(_06218_),
    .B(_06219_),
    .Y(_06220_));
 sky130_as_sc_hs__or2_2 _36951_ (.A(_06207_),
    .B(_06220_),
    .Y(_06222_));
 sky130_as_sc_hs__and2_2 _36952_ (.A(_06221_),
    .B(_06222_),
    .Y(_06223_));
 sky130_as_sc_hs__nand3_2 _36953_ (.A(_06206_),
    .B(_06221_),
    .C(_06222_),
    .Y(_06224_));
 sky130_as_sc_hs__or2_2 _36954_ (.A(_06206_),
    .B(_06223_),
    .Y(_06225_));
 sky130_as_sc_hs__and2_2 _36955_ (.A(_06224_),
    .B(_06225_),
    .Y(_06226_));
 sky130_as_sc_hs__or2_2 _36958_ (.A(_06226_),
    .B(_06227_),
    .Y(_06229_));
 sky130_as_sc_hs__and2_2 _36959_ (.A(_06228_),
    .B(_06229_),
    .Y(_06230_));
 sky130_as_sc_hs__or2_2 _36961_ (.A(_06205_),
    .B(_06230_),
    .Y(_06232_));
 sky130_as_sc_hs__and2_2 _36962_ (.A(_06231_),
    .B(_06232_),
    .Y(_06233_));
 sky130_as_sc_hs__or2_2 _36964_ (.A(_06185_),
    .B(_06233_),
    .Y(_06235_));
 sky130_as_sc_hs__and2_2 _36965_ (.A(_06234_),
    .B(_06235_),
    .Y(_06236_));
 sky130_as_sc_hs__or2_2 _36967_ (.A(_06184_),
    .B(_06236_),
    .Y(_06238_));
 sky130_as_sc_hs__and2_2 _36968_ (.A(_06237_),
    .B(_06238_),
    .Y(_06239_));
 sky130_as_sc_hs__nand3_2 _36972_ (.A(net455),
    .B(_24818_),
    .C(_24819_),
    .Y(_06243_));
 sky130_as_sc_hs__or2_2 _36974_ (.A(_06242_),
    .B(_06243_),
    .Y(_06245_));
 sky130_as_sc_hs__and2_2 _36975_ (.A(_06244_),
    .B(_06245_),
    .Y(_06246_));
 sky130_as_sc_hs__and2_2 _36976_ (.A(_24808_),
    .B(net420),
    .Y(_06247_));
 sky130_as_sc_hs__or2_2 _36978_ (.A(_06246_),
    .B(_06247_),
    .Y(_06249_));
 sky130_as_sc_hs__and2_2 _36979_ (.A(_06248_),
    .B(_06249_),
    .Y(_06250_));
 sky130_as_sc_hs__and2_2 _36980_ (.A(_24774_),
    .B(net428),
    .Y(_06251_));
 sky130_as_sc_hs__and2_2 _36981_ (.A(_24545_),
    .B(net441),
    .Y(_06252_));
 sky130_as_sc_hs__or2_2 _36982_ (.A(_06251_),
    .B(_06252_),
    .Y(_06253_));
 sky130_as_sc_hs__and2_2 _36984_ (.A(_06253_),
    .B(_06254_),
    .Y(_06255_));
 sky130_as_sc_hs__and2_2 _36985_ (.A(net123),
    .B(_24768_),
    .Y(_06256_));
 sky130_as_sc_hs__or2_2 _36987_ (.A(_06255_),
    .B(_06256_),
    .Y(_06258_));
 sky130_as_sc_hs__and2_2 _36988_ (.A(_06257_),
    .B(_06258_),
    .Y(_06259_));
 sky130_as_sc_hs__or2_2 _36991_ (.A(_06259_),
    .B(_06260_),
    .Y(_06262_));
 sky130_as_sc_hs__and2_2 _36992_ (.A(_06261_),
    .B(_06262_),
    .Y(_06263_));
 sky130_as_sc_hs__or2_2 _36994_ (.A(_06250_),
    .B(_06263_),
    .Y(_06265_));
 sky130_as_sc_hs__and2_2 _36995_ (.A(_06264_),
    .B(_06265_),
    .Y(_06266_));
 sky130_as_sc_hs__and2_2 _36998_ (.A(net475),
    .B(net445),
    .Y(_06269_));
 sky130_as_sc_hs__and2_2 _36999_ (.A(_24256_),
    .B(net435),
    .Y(_06270_));
 sky130_as_sc_hs__or2_2 _37000_ (.A(_06269_),
    .B(_06270_),
    .Y(_06271_));
 sky130_as_sc_hs__and2_2 _37002_ (.A(_06271_),
    .B(_06272_),
    .Y(_06273_));
 sky130_as_sc_hs__and2_2 _37003_ (.A(_24729_),
    .B(net432),
    .Y(_06274_));
 sky130_as_sc_hs__or2_2 _37005_ (.A(_06273_),
    .B(_06274_),
    .Y(_06276_));
 sky130_as_sc_hs__and2_2 _37006_ (.A(_06275_),
    .B(_06276_),
    .Y(_06277_));
 sky130_as_sc_hs__or2_2 _37008_ (.A(_06268_),
    .B(_06277_),
    .Y(_06279_));
 sky130_as_sc_hs__and2_2 _37009_ (.A(_06278_),
    .B(_06279_),
    .Y(_06280_));
 sky130_as_sc_hs__or2_2 _37011_ (.A(_06267_),
    .B(_06280_),
    .Y(_06282_));
 sky130_as_sc_hs__and2_2 _37012_ (.A(_06281_),
    .B(_06282_),
    .Y(_06283_));
 sky130_as_sc_hs__or2_2 _37015_ (.A(_06283_),
    .B(_06284_),
    .Y(_06286_));
 sky130_as_sc_hs__and2_2 _37016_ (.A(_06285_),
    .B(_06286_),
    .Y(_06287_));
 sky130_as_sc_hs__or2_2 _37018_ (.A(_06266_),
    .B(_06287_),
    .Y(_06289_));
 sky130_as_sc_hs__and2_2 _37019_ (.A(_06288_),
    .B(_06289_),
    .Y(_06290_));
 sky130_as_sc_hs__or2_2 _37021_ (.A(_06241_),
    .B(_06290_),
    .Y(_06292_));
 sky130_as_sc_hs__and2_2 _37022_ (.A(_06291_),
    .B(_06292_),
    .Y(_06293_));
 sky130_as_sc_hs__or2_2 _37024_ (.A(_06240_),
    .B(_06293_),
    .Y(_06295_));
 sky130_as_sc_hs__and2_2 _37025_ (.A(_06294_),
    .B(_06295_),
    .Y(_06296_));
 sky130_as_sc_hs__and2_2 _37028_ (.A(net473),
    .B(net449),
    .Y(_06299_));
 sky130_as_sc_hs__and2_2 _37029_ (.A(_24216_),
    .B(net426),
    .Y(_06300_));
 sky130_as_sc_hs__or2_2 _37030_ (.A(_06299_),
    .B(_06300_),
    .Y(_06301_));
 sky130_as_sc_hs__and2_2 _37032_ (.A(_06301_),
    .B(_06302_),
    .Y(_06303_));
 sky130_as_sc_hs__and2_2 _37033_ (.A(net479),
    .B(net451),
    .Y(_06304_));
 sky130_as_sc_hs__or2_2 _37035_ (.A(_06303_),
    .B(_06304_),
    .Y(_06306_));
 sky130_as_sc_hs__and2_2 _37036_ (.A(_06305_),
    .B(_06306_),
    .Y(_06307_));
 sky130_as_sc_hs__and2_2 _37037_ (.A(net480),
    .B(_24527_),
    .Y(_06308_));
 sky130_as_sc_hs__and2_2 _37038_ (.A(net477),
    .B(net89),
    .Y(_06309_));
 sky130_as_sc_hs__or2_2 _37039_ (.A(_06308_),
    .B(_06309_),
    .Y(_06310_));
 sky130_as_sc_hs__and2_2 _37041_ (.A(_06310_),
    .B(_06311_),
    .Y(_06312_));
 sky130_as_sc_hs__and2_2 _37042_ (.A(net88),
    .B(net439),
    .Y(_06313_));
 sky130_as_sc_hs__or2_2 _37044_ (.A(_06312_),
    .B(_06313_),
    .Y(_06315_));
 sky130_as_sc_hs__and2_2 _37045_ (.A(_06314_),
    .B(_06315_),
    .Y(_06316_));
 sky130_as_sc_hs__or2_2 _37048_ (.A(_06316_),
    .B(_06317_),
    .Y(_06319_));
 sky130_as_sc_hs__and2_2 _37049_ (.A(_06318_),
    .B(_06319_),
    .Y(_06320_));
 sky130_as_sc_hs__or2_2 _37051_ (.A(_06307_),
    .B(_06320_),
    .Y(_06322_));
 sky130_as_sc_hs__and2_2 _37052_ (.A(_06321_),
    .B(_06322_),
    .Y(_06323_));
 sky130_as_sc_hs__or2_2 _37054_ (.A(_06298_),
    .B(_06323_),
    .Y(_06325_));
 sky130_as_sc_hs__and2_2 _37055_ (.A(_06324_),
    .B(_06325_),
    .Y(_06326_));
 sky130_as_sc_hs__or2_2 _37057_ (.A(_06297_),
    .B(_06326_),
    .Y(_06328_));
 sky130_as_sc_hs__and2_2 _37058_ (.A(_06327_),
    .B(_06328_),
    .Y(_06329_));
 sky130_as_sc_hs__and2_2 _37061_ (.A(net464),
    .B(net78),
    .Y(_06332_));
 sky130_as_sc_hs__and2_2 _37062_ (.A(net462),
    .B(net443),
    .Y(_06333_));
 sky130_as_sc_hs__or2_2 _37063_ (.A(_06332_),
    .B(_06333_),
    .Y(_06334_));
 sky130_as_sc_hs__and2_2 _37065_ (.A(_06334_),
    .B(_06335_),
    .Y(_06336_));
 sky130_as_sc_hs__and2_2 _37066_ (.A(_23674_),
    .B(net461),
    .Y(_06337_));
 sky130_as_sc_hs__or2_2 _37068_ (.A(_06336_),
    .B(_06337_),
    .Y(_06339_));
 sky130_as_sc_hs__and2_2 _37069_ (.A(_06338_),
    .B(_06339_),
    .Y(_06340_));
 sky130_as_sc_hs__or2_2 _37071_ (.A(_06331_),
    .B(_06340_),
    .Y(_06342_));
 sky130_as_sc_hs__and2_2 _37072_ (.A(_06341_),
    .B(_06342_),
    .Y(_06343_));
 sky130_as_sc_hs__or2_2 _37074_ (.A(_06330_),
    .B(_06343_),
    .Y(_06345_));
 sky130_as_sc_hs__and2_2 _37075_ (.A(_06344_),
    .B(_06345_),
    .Y(_06346_));
 sky130_as_sc_hs__and2_2 _37076_ (.A(net470),
    .B(net446),
    .Y(_06347_));
 sky130_as_sc_hs__and2_2 _37077_ (.A(net467),
    .B(net85),
    .Y(_06348_));
 sky130_as_sc_hs__and2_2 _37078_ (.A(net469),
    .B(net452),
    .Y(_06349_));
 sky130_as_sc_hs__or2_2 _37079_ (.A(_06348_),
    .B(_06349_),
    .Y(_06350_));
 sky130_as_sc_hs__and2_2 _37081_ (.A(_06350_),
    .B(_06351_),
    .Y(_06352_));
 sky130_as_sc_hs__or2_2 _37083_ (.A(_06347_),
    .B(_06352_),
    .Y(_06354_));
 sky130_as_sc_hs__and2_2 _37084_ (.A(_06353_),
    .B(_06354_),
    .Y(_06355_));
 sky130_as_sc_hs__and2_2 _37085_ (.A(net456),
    .B(_24501_),
    .Y(_06356_));
 sky130_as_sc_hs__nand3_2 _37086_ (.A(_23598_),
    .B(net90),
    .C(_02549_),
    .Y(_06357_));
 sky130_as_sc_hs__nand3_2 _37087_ (.A(_24229_),
    .B(_25033_),
    .C(_25034_),
    .Y(_06358_));
 sky130_as_sc_hs__or2_2 _37089_ (.A(_06357_),
    .B(_06358_),
    .Y(_06360_));
 sky130_as_sc_hs__and2_2 _37090_ (.A(_06359_),
    .B(_06360_),
    .Y(_06361_));
 sky130_as_sc_hs__or2_2 _37092_ (.A(_06356_),
    .B(_06361_),
    .Y(_06363_));
 sky130_as_sc_hs__and2_2 _37093_ (.A(_06362_),
    .B(_06363_),
    .Y(_06364_));
 sky130_as_sc_hs__or2_2 _37096_ (.A(_06364_),
    .B(_06365_),
    .Y(_06367_));
 sky130_as_sc_hs__and2_2 _37097_ (.A(_06366_),
    .B(_06367_),
    .Y(_06368_));
 sky130_as_sc_hs__or2_2 _37099_ (.A(_06355_),
    .B(_06368_),
    .Y(_06370_));
 sky130_as_sc_hs__and2_2 _37100_ (.A(_06369_),
    .B(_06370_),
    .Y(_06371_));
 sky130_as_sc_hs__or2_2 _37103_ (.A(_06371_),
    .B(_06372_),
    .Y(_06374_));
 sky130_as_sc_hs__and2_2 _37104_ (.A(_06373_),
    .B(_06374_),
    .Y(_06375_));
 sky130_as_sc_hs__or2_2 _37106_ (.A(_06346_),
    .B(_06375_),
    .Y(_06377_));
 sky130_as_sc_hs__and2_2 _37107_ (.A(_06376_),
    .B(_06377_),
    .Y(_06378_));
 sky130_as_sc_hs__or2_2 _37110_ (.A(_06378_),
    .B(_06379_),
    .Y(_06381_));
 sky130_as_sc_hs__and2_2 _37111_ (.A(_06380_),
    .B(_06381_),
    .Y(_06382_));
 sky130_as_sc_hs__or2_2 _37113_ (.A(_06329_),
    .B(_06382_),
    .Y(_06384_));
 sky130_as_sc_hs__and2_2 _37114_ (.A(_06383_),
    .B(_06384_),
    .Y(_06385_));
 sky130_as_sc_hs__or2_2 _37117_ (.A(_06385_),
    .B(_06386_),
    .Y(_06388_));
 sky130_as_sc_hs__and2_2 _37118_ (.A(_06387_),
    .B(_06388_),
    .Y(_06389_));
 sky130_as_sc_hs__or2_2 _37120_ (.A(_06296_),
    .B(_06389_),
    .Y(_06391_));
 sky130_as_sc_hs__and2_2 _37121_ (.A(_06390_),
    .B(_06391_),
    .Y(_06392_));
 sky130_as_sc_hs__or2_2 _37124_ (.A(_06392_),
    .B(_06393_),
    .Y(_06395_));
 sky130_as_sc_hs__and2_2 _37125_ (.A(_06394_),
    .B(_06395_),
    .Y(_06396_));
 sky130_as_sc_hs__nand3_2 _37126_ (.A(_06237_),
    .B(_06238_),
    .C(_06396_),
    .Y(_06397_));
 sky130_as_sc_hs__or2_2 _37127_ (.A(_06239_),
    .B(_06396_),
    .Y(_06398_));
 sky130_as_sc_hs__and2_2 _37128_ (.A(_06397_),
    .B(_06398_),
    .Y(_06399_));
 sky130_as_sc_hs__or2_2 _37131_ (.A(_06399_),
    .B(_06400_),
    .Y(_06402_));
 sky130_as_sc_hs__and2_2 _37132_ (.A(_06401_),
    .B(_06402_),
    .Y(_06403_));
 sky130_as_sc_hs__nand3_2 _37133_ (.A(_06183_),
    .B(_06401_),
    .C(_06402_),
    .Y(_06404_));
 sky130_as_sc_hs__or2_2 _37134_ (.A(_06183_),
    .B(_06403_),
    .Y(_06405_));
 sky130_as_sc_hs__and2_2 _37135_ (.A(_06404_),
    .B(_06405_),
    .Y(_06406_));
 sky130_as_sc_hs__or2_2 _37138_ (.A(_06406_),
    .B(_06407_),
    .Y(_06409_));
 sky130_as_sc_hs__and2_2 _37139_ (.A(_06408_),
    .B(_06409_),
    .Y(_06410_));
 sky130_as_sc_hs__nand3_2 _37140_ (.A(_06182_),
    .B(_06408_),
    .C(_06409_),
    .Y(_06411_));
 sky130_as_sc_hs__or2_2 _37141_ (.A(_06182_),
    .B(_06410_),
    .Y(_06412_));
 sky130_as_sc_hs__and2_2 _37142_ (.A(_06411_),
    .B(_06412_),
    .Y(_06413_));
 sky130_as_sc_hs__nand3_2 _37144_ (.A(_06411_),
    .B(_06412_),
    .C(_06414_),
    .Y(_06415_));
 sky130_as_sc_hs__or2_2 _37145_ (.A(_06413_),
    .B(_06414_),
    .Y(_06416_));
 sky130_as_sc_hs__and2_2 _37146_ (.A(_06415_),
    .B(_06416_),
    .Y(_06417_));
 sky130_as_sc_hs__or2_2 _37148_ (.A(_06417_),
    .B(_06418_),
    .Y(_06419_));
 sky130_as_sc_hs__or2_2 _37152_ (.A(_06421_),
    .B(_06422_),
    .Y(_06423_));
 sky130_as_sc_hs__nand3_2 _37154_ (.A(net142),
    .B(_06423_),
    .C(_06424_),
    .Y(_06425_));
 sky130_as_sc_hs__and2_2 _37155_ (.A(_05946_),
    .B(_06132_),
    .Y(_06426_));
 sky130_as_sc_hs__nor2_2 _37156_ (.A(_05947_),
    .B(_06426_),
    .Y(_06427_));
 sky130_as_sc_hs__or2_2 _37157_ (.A(_05940_),
    .B(_06427_),
    .Y(_06428_));
 sky130_as_sc_hs__nand3_2 _37166_ (.A(_05946_),
    .B(_06435_),
    .C(_06436_),
    .Y(_06437_));
 sky130_as_sc_hs__and2_2 _37169_ (.A(_06438_),
    .B(_06439_),
    .Y(_06440_));
 sky130_as_sc_hs__and2_2 _37173_ (.A(_06442_),
    .B(_06443_),
    .Y(_06444_));
 sky130_as_sc_hs__or2_2 _37178_ (.A(net82),
    .B(_06448_),
    .Y(_06449_));
 sky130_as_sc_hs__and2_2 _37179_ (.A(_06445_),
    .B(_06449_),
    .Y(_06450_));
 sky130_as_sc_hs__nand3_2 _37181_ (.A(_05941_),
    .B(_06437_),
    .C(_06441_),
    .Y(_06452_));
 sky130_as_sc_hs__nand3_2 _37182_ (.A(_05935_),
    .B(_06451_),
    .C(_06452_),
    .Y(_06453_));
 sky130_as_sc_hs__and2_2 _37185_ (.A(_06454_),
    .B(_06455_),
    .Y(_06456_));
 sky130_as_sc_hs__or2_2 _37190_ (.A(net82),
    .B(_06460_),
    .Y(_06461_));
 sky130_as_sc_hs__or2_2 _37192_ (.A(_05940_),
    .B(_06462_),
    .Y(_06463_));
 sky130_as_sc_hs__and2_2 _37193_ (.A(_05950_),
    .B(_06075_),
    .Y(_06464_));
 sky130_as_sc_hs__and2_2 _37194_ (.A(_05951_),
    .B(_06035_),
    .Y(_06465_));
 sky130_as_sc_hs__or2_2 _37195_ (.A(_06464_),
    .B(_06465_),
    .Y(_06466_));
 sky130_as_sc_hs__and2_2 _37198_ (.A(_06467_),
    .B(_06468_),
    .Y(_06469_));
 sky130_as_sc_hs__or2_2 _37199_ (.A(net82),
    .B(_06469_),
    .Y(_06470_));
 sky130_as_sc_hs__and2_2 _37203_ (.A(_06463_),
    .B(_06473_),
    .Y(_06474_));
 sky130_as_sc_hs__and2_2 _37207_ (.A(_05950_),
    .B(_06139_),
    .Y(_06478_));
 sky130_as_sc_hs__and2_2 _37208_ (.A(_05951_),
    .B(_06107_),
    .Y(_06479_));
 sky130_as_sc_hs__or2_2 _37209_ (.A(_06478_),
    .B(_06479_),
    .Y(_06480_));
 sky130_as_sc_hs__and2_2 _37212_ (.A(_06481_),
    .B(_06482_),
    .Y(_06483_));
 sky130_as_sc_hs__or2_2 _37213_ (.A(net82),
    .B(_06483_),
    .Y(_06484_));
 sky130_as_sc_hs__or2_2 _37225_ (.A(_05935_),
    .B(_06495_),
    .Y(_06496_));
 sky130_as_sc_hs__and2_2 _37228_ (.A(_06497_),
    .B(_06498_),
    .Y(_06499_));
 sky130_as_sc_hs__or2_2 _37233_ (.A(net82),
    .B(_06503_),
    .Y(_06504_));
 sky130_as_sc_hs__and2_2 _37234_ (.A(_06500_),
    .B(_06504_),
    .Y(_06505_));
 sky130_as_sc_hs__and2_2 _37238_ (.A(_06507_),
    .B(_06508_),
    .Y(_06509_));
 sky130_as_sc_hs__and2_2 _37242_ (.A(_06511_),
    .B(_06512_),
    .Y(_06513_));
 sky130_as_sc_hs__and2_2 _37244_ (.A(_06510_),
    .B(_06514_),
    .Y(_06515_));
 sky130_as_sc_hs__and2_2 _37246_ (.A(_06506_),
    .B(_06516_),
    .Y(_06517_));
 sky130_as_sc_hs__and2_2 _37248_ (.A(_06496_),
    .B(_06518_),
    .Y(_06519_));
 sky130_as_sc_hs__or2_2 _37249_ (.A(_05929_),
    .B(_06519_),
    .Y(_06520_));
 sky130_as_sc_hs__and2_2 _37250_ (.A(_06477_),
    .B(_06520_),
    .Y(_06521_));
 sky130_as_sc_hs__and2_2 _37251_ (.A(_05968_),
    .B(_06521_),
    .Y(_06522_));
 sky130_as_sc_hs__nor2_2 _37252_ (.A(_19987_),
    .B(_23605_),
    .Y(_06523_));
 sky130_as_sc_hs__nor2_2 _37253_ (.A(_05836_),
    .B(_06153_),
    .Y(_06524_));
 sky130_as_sc_hs__and2_2 _37254_ (.A(_05836_),
    .B(_06153_),
    .Y(_06525_));
 sky130_as_sc_hs__or2_2 _37255_ (.A(_06524_),
    .B(_06525_),
    .Y(_06526_));
 sky130_as_sc_hs__and2_2 _37256_ (.A(\tholin_riscv.instr[5] ),
    .B(\tholin_riscv.Bimm[10] ),
    .Y(_06527_));
 sky130_as_sc_hs__or2_2 _37260_ (.A(_06526_),
    .B(_06529_),
    .Y(_06531_));
 sky130_as_sc_hs__nand3_2 _37261_ (.A(net119),
    .B(_06530_),
    .C(_06531_),
    .Y(_06532_));
 sky130_as_sc_hs__and2_2 _37262_ (.A(_04514_),
    .B(_05398_),
    .Y(_06533_));
 sky130_as_sc_hs__and2_2 _37263_ (.A(_05397_),
    .B(_05504_),
    .Y(_06534_));
 sky130_as_sc_hs__or2_2 _37264_ (.A(_06533_),
    .B(_06534_),
    .Y(_06535_));
 sky130_as_sc_hs__nand3_2 _37266_ (.A(net139),
    .B(_06535_),
    .C(_06536_),
    .Y(_06537_));
 sky130_as_sc_hs__and2_2 _37267_ (.A(_23603_),
    .B(_05967_),
    .Y(_06538_));
 sky130_as_sc_hs__or2_2 _37269_ (.A(_05834_),
    .B(_06539_),
    .Y(_06540_));
 sky130_as_sc_hs__and2_2 _37270_ (.A(_06158_),
    .B(_06540_),
    .Y(_06541_));
 sky130_as_sc_hs__or2_2 _37271_ (.A(_05835_),
    .B(_06541_),
    .Y(_06542_));
 sky130_as_sc_hs__and2_2 _37273_ (.A(net411),
    .B(_19487_),
    .Y(_06544_));
 sky130_as_sc_hs__inv_2 _37274_ (.Y(_06545_),
    .A(_06544_));
 sky130_as_sc_hs__and2_2 _37275_ (.A(_23598_),
    .B(_06544_),
    .Y(_06546_));
 sky130_as_sc_hs__and2_2 _37277_ (.A(_21655_),
    .B(_06544_),
    .Y(_06548_));
 sky130_as_sc_hs__and2_2 _37280_ (.A(_06543_),
    .B(_06550_),
    .Y(_06551_));
 sky130_as_sc_hs__and2_2 _37281_ (.A(\tholin_riscv.div_res[0] ),
    .B(net415),
    .Y(_06552_));
 sky130_as_sc_hs__or2_2 _37282_ (.A(\tholin_riscv.div_res[1] ),
    .B(_06552_),
    .Y(_06553_));
 sky130_as_sc_hs__and2_2 _37283_ (.A(\tholin_riscv.div_res[1] ),
    .B(_06552_),
    .Y(_06554_));
 sky130_as_sc_hs__and2_2 _37284_ (.A(_23603_),
    .B(_06165_),
    .Y(_06555_));
 sky130_as_sc_hs__or2_2 _37286_ (.A(_06554_),
    .B(_06556_),
    .Y(_06557_));
 sky130_as_sc_hs__and2_2 _37287_ (.A(_05834_),
    .B(_06160_),
    .Y(_06558_));
 sky130_as_sc_hs__and2_2 _37288_ (.A(\tholin_riscv.div_shifter[32] ),
    .B(_21655_),
    .Y(_06559_));
 sky130_as_sc_hs__or2_2 _37290_ (.A(\tholin_riscv.div_shifter[33] ),
    .B(_06559_),
    .Y(_06561_));
 sky130_as_sc_hs__and2_2 _37291_ (.A(_05512_),
    .B(_06165_),
    .Y(_06562_));
 sky130_as_sc_hs__nand3_2 _37292_ (.A(_06560_),
    .B(_06561_),
    .C(net109),
    .Y(_06563_));
 sky130_as_sc_hs__and2_2 _37293_ (.A(_23599_),
    .B(_06165_),
    .Y(_06564_));
 sky130_as_sc_hs__and2_2 _37295_ (.A(_21656_),
    .B(_06165_),
    .Y(_06566_));
 sky130_as_sc_hs__and2_2 _37297_ (.A(_06565_),
    .B(_06567_),
    .Y(_06568_));
 sky130_as_sc_hs__nand3_2 _37298_ (.A(net413),
    .B(_06563_),
    .C(_06568_),
    .Y(_06569_));
 sky130_as_sc_hs__nor2_2 _37299_ (.A(_06558_),
    .B(_06569_),
    .Y(_06570_));
 sky130_as_sc_hs__and2_2 _37300_ (.A(_06542_),
    .B(_06570_),
    .Y(_06571_));
 sky130_as_sc_hs__and2_2 _37301_ (.A(_06557_),
    .B(_06571_),
    .Y(_06572_));
 sky130_as_sc_hs__nand3_2 _37302_ (.A(_06532_),
    .B(_06537_),
    .C(_06572_),
    .Y(_06573_));
 sky130_as_sc_hs__nor2_2 _37303_ (.A(_06522_),
    .B(_06573_),
    .Y(_06574_));
 sky130_as_sc_hs__nand3_2 _37304_ (.A(_06425_),
    .B(_06434_),
    .C(_06574_),
    .Y(_06575_));
 sky130_as_sc_hs__nand3_2 _37307_ (.A(_21546_),
    .B(_06575_),
    .C(_06577_),
    .Y(_06578_));
 sky130_as_sc_hs__and2_2 _37317_ (.A(net123),
    .B(_23636_),
    .Y(_06587_));
 sky130_as_sc_hs__and2_2 _37318_ (.A(_24216_),
    .B(net422),
    .Y(_06588_));
 sky130_as_sc_hs__or2_2 _37319_ (.A(_06587_),
    .B(_06588_),
    .Y(_06589_));
 sky130_as_sc_hs__and2_2 _37321_ (.A(_06589_),
    .B(_06590_),
    .Y(_06591_));
 sky130_as_sc_hs__and2_2 _37322_ (.A(net483),
    .B(net432),
    .Y(_06592_));
 sky130_as_sc_hs__or2_2 _37324_ (.A(_06591_),
    .B(_06592_),
    .Y(_06594_));
 sky130_as_sc_hs__and2_2 _37325_ (.A(_06593_),
    .B(_06594_),
    .Y(_06595_));
 sky130_as_sc_hs__or2_2 _37328_ (.A(_06595_),
    .B(_06596_),
    .Y(_06598_));
 sky130_as_sc_hs__or2_2 _37330_ (.A(_06196_),
    .B(_06599_),
    .Y(_06600_));
 sky130_as_sc_hs__and2_2 _37332_ (.A(_06600_),
    .B(_06601_),
    .Y(_06602_));
 sky130_as_sc_hs__and2_2 _37333_ (.A(_23702_),
    .B(net428),
    .Y(_06603_));
 sky130_as_sc_hs__or2_2 _37335_ (.A(_06602_),
    .B(_06603_),
    .Y(_06605_));
 sky130_as_sc_hs__and2_2 _37336_ (.A(_06604_),
    .B(_06605_),
    .Y(_06606_));
 sky130_as_sc_hs__and2_2 _37340_ (.A(_23712_),
    .B(net129),
    .Y(_06610_));
 sky130_as_sc_hs__or2_2 _37342_ (.A(_06609_),
    .B(_06610_),
    .Y(_06612_));
 sky130_as_sc_hs__or2_2 _37344_ (.A(_06212_),
    .B(_06613_),
    .Y(_06614_));
 sky130_as_sc_hs__and2_2 _37346_ (.A(_06614_),
    .B(_06615_),
    .Y(_06616_));
 sky130_as_sc_hs__or2_2 _37348_ (.A(_06608_),
    .B(_06616_),
    .Y(_06618_));
 sky130_as_sc_hs__and2_2 _37349_ (.A(_06617_),
    .B(_06618_),
    .Y(_06619_));
 sky130_as_sc_hs__or2_2 _37351_ (.A(_06607_),
    .B(_06619_),
    .Y(_06621_));
 sky130_as_sc_hs__and2_2 _37352_ (.A(_06620_),
    .B(_06621_),
    .Y(_06622_));
 sky130_as_sc_hs__or2_2 _37355_ (.A(_06622_),
    .B(_06623_),
    .Y(_06625_));
 sky130_as_sc_hs__and2_2 _37356_ (.A(_06624_),
    .B(_06625_),
    .Y(_06626_));
 sky130_as_sc_hs__or2_2 _37358_ (.A(_06606_),
    .B(_06626_),
    .Y(_06628_));
 sky130_as_sc_hs__and2_2 _37359_ (.A(_06627_),
    .B(_06628_),
    .Y(_06629_));
 sky130_as_sc_hs__or2_2 _37361_ (.A(_06586_),
    .B(_06629_),
    .Y(_06631_));
 sky130_as_sc_hs__and2_2 _37362_ (.A(_06630_),
    .B(_06631_),
    .Y(_06632_));
 sky130_as_sc_hs__or2_2 _37364_ (.A(_06585_),
    .B(_06632_),
    .Y(_06634_));
 sky130_as_sc_hs__and2_2 _37365_ (.A(_06633_),
    .B(_06634_),
    .Y(_06635_));
 sky130_as_sc_hs__and2_2 _37368_ (.A(_24814_),
    .B(net420),
    .Y(_06638_));
 sky130_as_sc_hs__and2_2 _37369_ (.A(net86),
    .B(net437),
    .Y(_06639_));
 sky130_as_sc_hs__or2_2 _37370_ (.A(_06638_),
    .B(_06639_),
    .Y(_06640_));
 sky130_as_sc_hs__and2_2 _37372_ (.A(_06640_),
    .B(_06641_),
    .Y(_06642_));
 sky130_as_sc_hs__and2_2 _37373_ (.A(_24808_),
    .B(net75),
    .Y(_06643_));
 sky130_as_sc_hs__or2_2 _37375_ (.A(_06642_),
    .B(_06643_),
    .Y(_06645_));
 sky130_as_sc_hs__and2_2 _37376_ (.A(_06644_),
    .B(_06645_),
    .Y(_06646_));
 sky130_as_sc_hs__and2_2 _37377_ (.A(_24768_),
    .B(net424),
    .Y(_06647_));
 sky130_as_sc_hs__nand3_2 _37378_ (.A(_23689_),
    .B(_23690_),
    .C(_24774_),
    .Y(_06648_));
 sky130_as_sc_hs__or2_2 _37381_ (.A(_06648_),
    .B(_06649_),
    .Y(_06651_));
 sky130_as_sc_hs__and2_2 _37382_ (.A(_06650_),
    .B(_06651_),
    .Y(_06652_));
 sky130_as_sc_hs__or2_2 _37384_ (.A(_06647_),
    .B(_06652_),
    .Y(_06654_));
 sky130_as_sc_hs__and2_2 _37385_ (.A(_06653_),
    .B(_06654_),
    .Y(_06655_));
 sky130_as_sc_hs__or2_2 _37388_ (.A(_06655_),
    .B(_06656_),
    .Y(_06658_));
 sky130_as_sc_hs__and2_2 _37389_ (.A(_06657_),
    .B(_06658_),
    .Y(_06659_));
 sky130_as_sc_hs__or2_2 _37391_ (.A(_06646_),
    .B(_06659_),
    .Y(_06661_));
 sky130_as_sc_hs__and2_2 _37392_ (.A(_06660_),
    .B(_06661_),
    .Y(_06662_));
 sky130_as_sc_hs__and2_2 _37395_ (.A(net445),
    .B(net84),
    .Y(_06665_));
 sky130_as_sc_hs__and2_2 _37396_ (.A(_24501_),
    .B(net435),
    .Y(_06666_));
 sky130_as_sc_hs__or2_2 _37397_ (.A(_06665_),
    .B(_06666_),
    .Y(_06667_));
 sky130_as_sc_hs__and2_2 _37399_ (.A(_06667_),
    .B(_06668_),
    .Y(_06669_));
 sky130_as_sc_hs__and2_2 _37400_ (.A(_24729_),
    .B(net430),
    .Y(_06670_));
 sky130_as_sc_hs__or2_2 _37402_ (.A(_06669_),
    .B(_06670_),
    .Y(_06672_));
 sky130_as_sc_hs__and2_2 _37403_ (.A(_06671_),
    .B(_06672_),
    .Y(_06673_));
 sky130_as_sc_hs__or2_2 _37405_ (.A(_06664_),
    .B(_06673_),
    .Y(_06675_));
 sky130_as_sc_hs__and2_2 _37406_ (.A(_06674_),
    .B(_06675_),
    .Y(_06676_));
 sky130_as_sc_hs__or2_2 _37408_ (.A(_06663_),
    .B(_06676_),
    .Y(_06678_));
 sky130_as_sc_hs__and2_2 _37409_ (.A(_06677_),
    .B(_06678_),
    .Y(_06679_));
 sky130_as_sc_hs__or2_2 _37412_ (.A(_06679_),
    .B(_06680_),
    .Y(_06682_));
 sky130_as_sc_hs__and2_2 _37413_ (.A(_06681_),
    .B(_06682_),
    .Y(_06683_));
 sky130_as_sc_hs__or2_2 _37415_ (.A(_06662_),
    .B(_06683_),
    .Y(_06685_));
 sky130_as_sc_hs__and2_2 _37416_ (.A(_06684_),
    .B(_06685_),
    .Y(_06686_));
 sky130_as_sc_hs__or2_2 _37418_ (.A(_06637_),
    .B(_06686_),
    .Y(_06688_));
 sky130_as_sc_hs__and2_2 _37419_ (.A(_06687_),
    .B(_06688_),
    .Y(_06689_));
 sky130_as_sc_hs__or2_2 _37421_ (.A(_06636_),
    .B(_06689_),
    .Y(_06691_));
 sky130_as_sc_hs__and2_2 _37422_ (.A(_06690_),
    .B(_06691_),
    .Y(_06692_));
 sky130_as_sc_hs__and2_2 _37425_ (.A(net479),
    .B(net449),
    .Y(_06695_));
 sky130_as_sc_hs__and2_2 _37426_ (.A(_24229_),
    .B(net426),
    .Y(_06696_));
 sky130_as_sc_hs__or2_2 _37427_ (.A(_06695_),
    .B(_06696_),
    .Y(_06697_));
 sky130_as_sc_hs__and2_2 _37429_ (.A(_06697_),
    .B(_06698_),
    .Y(_06699_));
 sky130_as_sc_hs__and2_2 _37430_ (.A(net475),
    .B(net451),
    .Y(_06700_));
 sky130_as_sc_hs__or2_2 _37432_ (.A(_06699_),
    .B(_06700_),
    .Y(_06702_));
 sky130_as_sc_hs__and2_2 _37433_ (.A(_06701_),
    .B(_06702_),
    .Y(_06703_));
 sky130_as_sc_hs__and2_2 _37434_ (.A(net477),
    .B(_24527_),
    .Y(_06704_));
 sky130_as_sc_hs__and2_2 _37435_ (.A(net89),
    .B(net439),
    .Y(_06705_));
 sky130_as_sc_hs__or2_2 _37436_ (.A(_06704_),
    .B(_06705_),
    .Y(_06706_));
 sky130_as_sc_hs__and2_2 _37438_ (.A(_06706_),
    .B(_06707_),
    .Y(_06708_));
 sky130_as_sc_hs__and2_2 _37439_ (.A(_23680_),
    .B(net88),
    .Y(_06709_));
 sky130_as_sc_hs__or2_2 _37441_ (.A(_06708_),
    .B(_06709_),
    .Y(_06711_));
 sky130_as_sc_hs__and2_2 _37442_ (.A(_06710_),
    .B(_06711_),
    .Y(_06712_));
 sky130_as_sc_hs__or2_2 _37445_ (.A(_06712_),
    .B(_06713_),
    .Y(_06715_));
 sky130_as_sc_hs__and2_2 _37446_ (.A(_06714_),
    .B(_06715_),
    .Y(_06716_));
 sky130_as_sc_hs__or2_2 _37448_ (.A(_06703_),
    .B(_06716_),
    .Y(_06718_));
 sky130_as_sc_hs__and2_2 _37449_ (.A(_06717_),
    .B(_06718_),
    .Y(_06719_));
 sky130_as_sc_hs__or2_2 _37451_ (.A(_06694_),
    .B(_06719_),
    .Y(_06721_));
 sky130_as_sc_hs__and2_2 _37452_ (.A(_06720_),
    .B(_06721_),
    .Y(_06722_));
 sky130_as_sc_hs__or2_2 _37454_ (.A(_06693_),
    .B(_06722_),
    .Y(_06724_));
 sky130_as_sc_hs__and2_2 _37455_ (.A(_06723_),
    .B(_06724_),
    .Y(_06725_));
 sky130_as_sc_hs__and2_2 _37458_ (.A(net464),
    .B(net443),
    .Y(_06728_));
 sky130_as_sc_hs__and2_2 _37459_ (.A(_23674_),
    .B(net462),
    .Y(_06729_));
 sky130_as_sc_hs__or2_2 _37460_ (.A(_06728_),
    .B(_06729_),
    .Y(_06730_));
 sky130_as_sc_hs__and2_2 _37462_ (.A(_06730_),
    .B(_06731_),
    .Y(_06732_));
 sky130_as_sc_hs__and2_2 _37463_ (.A(_23629_),
    .B(net461),
    .Y(_06733_));
 sky130_as_sc_hs__or2_2 _37465_ (.A(_06732_),
    .B(_06733_),
    .Y(_06735_));
 sky130_as_sc_hs__and2_2 _37466_ (.A(_06734_),
    .B(_06735_),
    .Y(_06736_));
 sky130_as_sc_hs__or2_2 _37468_ (.A(_06727_),
    .B(_06736_),
    .Y(_06738_));
 sky130_as_sc_hs__and2_2 _37469_ (.A(_06737_),
    .B(_06738_),
    .Y(_06739_));
 sky130_as_sc_hs__or2_2 _37471_ (.A(_06726_),
    .B(_06739_),
    .Y(_06741_));
 sky130_as_sc_hs__and2_2 _37472_ (.A(_06740_),
    .B(_06741_),
    .Y(_06742_));
 sky130_as_sc_hs__and2_2 _37473_ (.A(net470),
    .B(net78),
    .Y(_06743_));
 sky130_as_sc_hs__and2_2 _37474_ (.A(net467),
    .B(net452),
    .Y(_06744_));
 sky130_as_sc_hs__and2_2 _37475_ (.A(net469),
    .B(net446),
    .Y(_06745_));
 sky130_as_sc_hs__or2_2 _37476_ (.A(_06744_),
    .B(_06745_),
    .Y(_06746_));
 sky130_as_sc_hs__and2_2 _37478_ (.A(_06746_),
    .B(_06747_),
    .Y(_06748_));
 sky130_as_sc_hs__or2_2 _37480_ (.A(_06743_),
    .B(_06748_),
    .Y(_06750_));
 sky130_as_sc_hs__and2_2 _37481_ (.A(_06749_),
    .B(_06750_),
    .Y(_06751_));
 sky130_as_sc_hs__and2_2 _37482_ (.A(net456),
    .B(_24545_),
    .Y(_06752_));
 sky130_as_sc_hs__nand3_2 _37483_ (.A(_23598_),
    .B(_24053_),
    .C(_02549_),
    .Y(_06753_));
 sky130_as_sc_hs__nand3_2 _37484_ (.A(_24256_),
    .B(_25033_),
    .C(_25034_),
    .Y(_06754_));
 sky130_as_sc_hs__or2_2 _37486_ (.A(_06753_),
    .B(_06754_),
    .Y(_06756_));
 sky130_as_sc_hs__and2_2 _37487_ (.A(_06755_),
    .B(_06756_),
    .Y(_06757_));
 sky130_as_sc_hs__or2_2 _37489_ (.A(_06752_),
    .B(_06757_),
    .Y(_06759_));
 sky130_as_sc_hs__and2_2 _37490_ (.A(_06758_),
    .B(_06759_),
    .Y(_06760_));
 sky130_as_sc_hs__or2_2 _37493_ (.A(_06760_),
    .B(_06761_),
    .Y(_06763_));
 sky130_as_sc_hs__and2_2 _37494_ (.A(_06762_),
    .B(_06763_),
    .Y(_06764_));
 sky130_as_sc_hs__or2_2 _37496_ (.A(_06751_),
    .B(_06764_),
    .Y(_06766_));
 sky130_as_sc_hs__and2_2 _37497_ (.A(_06765_),
    .B(_06766_),
    .Y(_06767_));
 sky130_as_sc_hs__or2_2 _37500_ (.A(_06767_),
    .B(_06768_),
    .Y(_06770_));
 sky130_as_sc_hs__and2_2 _37501_ (.A(_06769_),
    .B(_06770_),
    .Y(_06771_));
 sky130_as_sc_hs__or2_2 _37503_ (.A(_06742_),
    .B(_06771_),
    .Y(_06773_));
 sky130_as_sc_hs__and2_2 _37504_ (.A(_06772_),
    .B(_06773_),
    .Y(_06774_));
 sky130_as_sc_hs__or2_2 _37507_ (.A(_06774_),
    .B(_06775_),
    .Y(_06777_));
 sky130_as_sc_hs__and2_2 _37508_ (.A(_06776_),
    .B(_06777_),
    .Y(_06778_));
 sky130_as_sc_hs__or2_2 _37510_ (.A(_06725_),
    .B(_06778_),
    .Y(_06780_));
 sky130_as_sc_hs__and2_2 _37511_ (.A(_06779_),
    .B(_06780_),
    .Y(_06781_));
 sky130_as_sc_hs__or2_2 _37514_ (.A(_06781_),
    .B(_06782_),
    .Y(_06784_));
 sky130_as_sc_hs__and2_2 _37515_ (.A(_06783_),
    .B(_06784_),
    .Y(_06785_));
 sky130_as_sc_hs__or2_2 _37517_ (.A(_06692_),
    .B(_06785_),
    .Y(_06787_));
 sky130_as_sc_hs__and2_2 _37518_ (.A(_06786_),
    .B(_06787_),
    .Y(_06788_));
 sky130_as_sc_hs__or2_2 _37521_ (.A(_06788_),
    .B(_06789_),
    .Y(_06791_));
 sky130_as_sc_hs__and2_2 _37522_ (.A(_06790_),
    .B(_06791_),
    .Y(_06792_));
 sky130_as_sc_hs__or2_2 _37524_ (.A(_06635_),
    .B(_06792_),
    .Y(_06794_));
 sky130_as_sc_hs__and2_2 _37525_ (.A(_06793_),
    .B(_06794_),
    .Y(_06795_));
 sky130_as_sc_hs__or2_2 _37528_ (.A(_06795_),
    .B(_06796_),
    .Y(_06798_));
 sky130_as_sc_hs__and2_2 _37529_ (.A(_06797_),
    .B(_06798_),
    .Y(_06799_));
 sky130_as_sc_hs__or2_2 _37531_ (.A(_06584_),
    .B(_06799_),
    .Y(_06801_));
 sky130_as_sc_hs__and2_2 _37532_ (.A(_06800_),
    .B(_06801_),
    .Y(_06802_));
 sky130_as_sc_hs__or2_2 _37535_ (.A(_06802_),
    .B(_06803_),
    .Y(_06805_));
 sky130_as_sc_hs__and2_2 _37536_ (.A(_06804_),
    .B(_06805_),
    .Y(_06806_));
 sky130_as_sc_hs__or2_2 _37538_ (.A(_06583_),
    .B(_06806_),
    .Y(_06808_));
 sky130_as_sc_hs__and2_2 _37539_ (.A(_06807_),
    .B(_06808_),
    .Y(_06809_));
 sky130_as_sc_hs__or2_2 _37542_ (.A(_06809_),
    .B(_06810_),
    .Y(_06812_));
 sky130_as_sc_hs__and2_2 _37543_ (.A(_06811_),
    .B(_06812_),
    .Y(_06813_));
 sky130_as_sc_hs__and2_2 _37546_ (.A(_05364_),
    .B(_06417_),
    .Y(_06816_));
 sky130_as_sc_hs__or2_2 _37550_ (.A(_06813_),
    .B(_06818_),
    .Y(_06820_));
 sky130_as_sc_hs__and2_2 _37554_ (.A(_05506_),
    .B(_06823_),
    .Y(_06824_));
 sky130_as_sc_hs__or2_2 _37555_ (.A(_06821_),
    .B(_06824_),
    .Y(_06825_));
 sky130_as_sc_hs__nand3_2 _37557_ (.A(net142),
    .B(_06825_),
    .C(_06826_),
    .Y(_06827_));
 sky130_as_sc_hs__and2_2 _37558_ (.A(_05946_),
    .B(_06041_),
    .Y(_06828_));
 sky130_as_sc_hs__and2_2 _37559_ (.A(net82),
    .B(_06077_),
    .Y(_06829_));
 sky130_as_sc_hs__nor2_2 _37560_ (.A(_06828_),
    .B(_06829_),
    .Y(_06830_));
 sky130_as_sc_hs__or2_2 _37567_ (.A(_05935_),
    .B(_06836_),
    .Y(_06837_));
 sky130_as_sc_hs__or2_2 _37569_ (.A(net82),
    .B(_05985_),
    .Y(_06839_));
 sky130_as_sc_hs__or2_2 _37570_ (.A(net82),
    .B(_05995_),
    .Y(_06840_));
 sky130_as_sc_hs__and2_2 _37572_ (.A(_06840_),
    .B(_06841_),
    .Y(_06842_));
 sky130_as_sc_hs__nand3_2 _37574_ (.A(_05941_),
    .B(_06838_),
    .C(_06839_),
    .Y(_06844_));
 sky130_as_sc_hs__nand3_2 _37575_ (.A(_05935_),
    .B(_06843_),
    .C(_06844_),
    .Y(_06845_));
 sky130_as_sc_hs__and2_2 _37581_ (.A(_06849_),
    .B(_06850_),
    .Y(_06851_));
 sky130_as_sc_hs__or2_2 _37582_ (.A(_05935_),
    .B(_06851_),
    .Y(_06852_));
 sky130_as_sc_hs__and2_2 _37593_ (.A(_06852_),
    .B(_06862_),
    .Y(_06863_));
 sky130_as_sc_hs__nand3_2 _37594_ (.A(_05929_),
    .B(_06837_),
    .C(_06845_),
    .Y(_06864_));
 sky130_as_sc_hs__or2_2 _37595_ (.A(_05929_),
    .B(_06863_),
    .Y(_06865_));
 sky130_as_sc_hs__and2_2 _37596_ (.A(_06864_),
    .B(_06865_),
    .Y(_06866_));
 sky130_as_sc_hs__or2_2 _37598_ (.A(_05824_),
    .B(_05849_),
    .Y(_06868_));
 sky130_as_sc_hs__nand3_2 _37599_ (.A(_05850_),
    .B(_06527_),
    .C(_06868_),
    .Y(_06869_));
 sky130_as_sc_hs__nor2_2 _37600_ (.A(_05834_),
    .B(_06524_),
    .Y(_06870_));
 sky130_as_sc_hs__or2_2 _37601_ (.A(_05824_),
    .B(_06870_),
    .Y(_06871_));
 sky130_as_sc_hs__or2_2 _37604_ (.A(_06527_),
    .B(_06873_),
    .Y(_06874_));
 sky130_as_sc_hs__and2_2 _37606_ (.A(net119),
    .B(_06875_),
    .Y(_06876_));
 sky130_as_sc_hs__or2_2 _37607_ (.A(_05822_),
    .B(_06539_),
    .Y(_06877_));
 sky130_as_sc_hs__and2_2 _37608_ (.A(_06158_),
    .B(_06877_),
    .Y(_06878_));
 sky130_as_sc_hs__or2_2 _37609_ (.A(_05823_),
    .B(_06878_),
    .Y(_06879_));
 sky130_as_sc_hs__or2_2 _37610_ (.A(\tholin_riscv.div_res[1] ),
    .B(\tholin_riscv.div_res[0] ),
    .Y(_06880_));
 sky130_as_sc_hs__and2_2 _37611_ (.A(net415),
    .B(_06880_),
    .Y(_06881_));
 sky130_as_sc_hs__or2_2 _37613_ (.A(\tholin_riscv.div_res[2] ),
    .B(_06881_),
    .Y(_06883_));
 sky130_as_sc_hs__nand3_2 _37614_ (.A(net111),
    .B(_06882_),
    .C(_06883_),
    .Y(_06884_));
 sky130_as_sc_hs__and2_2 _37615_ (.A(_05822_),
    .B(_06160_),
    .Y(_06885_));
 sky130_as_sc_hs__or2_2 _37616_ (.A(\tholin_riscv.div_shifter[33] ),
    .B(\tholin_riscv.div_shifter[32] ),
    .Y(_06886_));
 sky130_as_sc_hs__and2_2 _37617_ (.A(_21655_),
    .B(_06886_),
    .Y(_06887_));
 sky130_as_sc_hs__or2_2 _37619_ (.A(\tholin_riscv.div_shifter[34] ),
    .B(_06887_),
    .Y(_06889_));
 sky130_as_sc_hs__nand3_2 _37620_ (.A(net109),
    .B(_06888_),
    .C(_06889_),
    .Y(_06890_));
 sky130_as_sc_hs__and2_2 _37623_ (.A(_06891_),
    .B(_06892_),
    .Y(_06893_));
 sky130_as_sc_hs__nand3_2 _37624_ (.A(net413),
    .B(_06890_),
    .C(_06893_),
    .Y(_06894_));
 sky130_as_sc_hs__nor2_2 _37625_ (.A(_06885_),
    .B(_06894_),
    .Y(_06895_));
 sky130_as_sc_hs__nand3_2 _37626_ (.A(_06879_),
    .B(_06884_),
    .C(_06895_),
    .Y(_06896_));
 sky130_as_sc_hs__nor2_2 _37627_ (.A(_06876_),
    .B(_06896_),
    .Y(_06897_));
 sky130_as_sc_hs__and2_2 _37628_ (.A(_06867_),
    .B(_06897_),
    .Y(_06898_));
 sky130_as_sc_hs__and2_2 _37629_ (.A(_04511_),
    .B(_04514_),
    .Y(_06899_));
 sky130_as_sc_hs__or2_2 _37630_ (.A(_04515_),
    .B(_06899_),
    .Y(_06900_));
 sky130_as_sc_hs__or2_2 _37631_ (.A(_05399_),
    .B(_05505_),
    .Y(_06901_));
 sky130_as_sc_hs__or2_2 _37633_ (.A(_06900_),
    .B(_06901_),
    .Y(_06903_));
 sky130_as_sc_hs__nand3_2 _37634_ (.A(net139),
    .B(_06902_),
    .C(_06903_),
    .Y(_06904_));
 sky130_as_sc_hs__and2_2 _37642_ (.A(_06904_),
    .B(_06911_),
    .Y(_06912_));
 sky130_as_sc_hs__nand3_2 _37643_ (.A(_06827_),
    .B(_06898_),
    .C(_06912_),
    .Y(_06913_));
 sky130_as_sc_hs__and2_2 _37644_ (.A(_19472_),
    .B(_21572_),
    .Y(_06914_));
 sky130_as_sc_hs__nand3_2 _37647_ (.A(_21569_),
    .B(_06915_),
    .C(_06916_),
    .Y(_06917_));
 sky130_as_sc_hs__nand3_2 _37648_ (.A(_21546_),
    .B(_06913_),
    .C(_06917_),
    .Y(_06918_));
 sky130_as_sc_hs__and2_2 _37659_ (.A(_23636_),
    .B(_25874_),
    .Y(_06928_));
 sky130_as_sc_hs__and2_2 _37660_ (.A(_24229_),
    .B(net422),
    .Y(_06929_));
 sky130_as_sc_hs__or2_2 _37661_ (.A(_06928_),
    .B(_06929_),
    .Y(_06930_));
 sky130_as_sc_hs__and2_2 _37663_ (.A(_06930_),
    .B(_06931_),
    .Y(_06932_));
 sky130_as_sc_hs__and2_2 _37664_ (.A(net483),
    .B(net430),
    .Y(_06933_));
 sky130_as_sc_hs__or2_2 _37666_ (.A(_06932_),
    .B(_06933_),
    .Y(_06935_));
 sky130_as_sc_hs__and2_2 _37667_ (.A(_06934_),
    .B(_06935_),
    .Y(_06936_));
 sky130_as_sc_hs__or2_2 _37670_ (.A(_06936_),
    .B(_06937_),
    .Y(_06939_));
 sky130_as_sc_hs__or2_2 _37672_ (.A(_06597_),
    .B(_06940_),
    .Y(_06941_));
 sky130_as_sc_hs__and2_2 _37674_ (.A(_06941_),
    .B(_06942_),
    .Y(_06943_));
 sky130_as_sc_hs__and2_2 _37675_ (.A(net121),
    .B(_23702_),
    .Y(_06944_));
 sky130_as_sc_hs__or2_2 _37677_ (.A(_06943_),
    .B(_06944_),
    .Y(_06946_));
 sky130_as_sc_hs__and2_2 _37678_ (.A(_06945_),
    .B(_06946_),
    .Y(_06947_));
 sky130_as_sc_hs__and2_2 _37682_ (.A(_24216_),
    .B(net129),
    .Y(_06951_));
 sky130_as_sc_hs__or2_2 _37684_ (.A(_06950_),
    .B(_06951_),
    .Y(_06953_));
 sky130_as_sc_hs__and2_2 _37685_ (.A(_06952_),
    .B(_06953_),
    .Y(_06954_));
 sky130_as_sc_hs__or2_2 _37687_ (.A(_06949_),
    .B(_06954_),
    .Y(_06956_));
 sky130_as_sc_hs__and2_2 _37688_ (.A(_06955_),
    .B(_06956_),
    .Y(_06957_));
 sky130_as_sc_hs__or2_2 _37690_ (.A(_06948_),
    .B(_06957_),
    .Y(_06959_));
 sky130_as_sc_hs__and2_2 _37691_ (.A(_06958_),
    .B(_06959_),
    .Y(_06960_));
 sky130_as_sc_hs__or2_2 _37694_ (.A(_06960_),
    .B(_06961_),
    .Y(_06963_));
 sky130_as_sc_hs__and2_2 _37695_ (.A(_06962_),
    .B(_06963_),
    .Y(_06964_));
 sky130_as_sc_hs__or2_2 _37697_ (.A(_06947_),
    .B(_06964_),
    .Y(_06966_));
 sky130_as_sc_hs__and2_2 _37698_ (.A(_06965_),
    .B(_06966_),
    .Y(_06967_));
 sky130_as_sc_hs__or2_2 _37700_ (.A(_06927_),
    .B(_06967_),
    .Y(_06969_));
 sky130_as_sc_hs__and2_2 _37701_ (.A(_06968_),
    .B(_06969_),
    .Y(_06970_));
 sky130_as_sc_hs__or2_2 _37703_ (.A(_06926_),
    .B(_06970_),
    .Y(_06972_));
 sky130_as_sc_hs__and2_2 _37704_ (.A(_06971_),
    .B(_06972_),
    .Y(_06973_));
 sky130_as_sc_hs__and2_2 _37707_ (.A(_24814_),
    .B(net75),
    .Y(_06976_));
 sky130_as_sc_hs__and2_2 _37708_ (.A(net452),
    .B(net437),
    .Y(_06977_));
 sky130_as_sc_hs__and2_2 _37709_ (.A(_06976_),
    .B(_06977_),
    .Y(_06978_));
 sky130_as_sc_hs__or2_2 _37710_ (.A(_06976_),
    .B(_06977_),
    .Y(_06979_));
 sky130_as_sc_hs__nor2b_2 _37711_ (.A(_06978_),
    .Y(_06980_),
    .B(_06979_));
 sky130_as_sc_hs__and2_2 _37712_ (.A(net123),
    .B(_24774_),
    .Y(_06981_));
 sky130_as_sc_hs__and2_2 _37713_ (.A(net85),
    .B(net441),
    .Y(_06982_));
 sky130_as_sc_hs__or2_2 _37714_ (.A(_06981_),
    .B(_06982_),
    .Y(_06983_));
 sky130_as_sc_hs__and2_2 _37716_ (.A(_06983_),
    .B(_06984_),
    .Y(_06985_));
 sky130_as_sc_hs__and2_2 _37717_ (.A(_24768_),
    .B(net420),
    .Y(_06986_));
 sky130_as_sc_hs__or2_2 _37719_ (.A(_06985_),
    .B(_06986_),
    .Y(_06988_));
 sky130_as_sc_hs__and2_2 _37720_ (.A(_06987_),
    .B(_06988_),
    .Y(_06989_));
 sky130_as_sc_hs__or2_2 _37723_ (.A(_06989_),
    .B(_06990_),
    .Y(_06992_));
 sky130_as_sc_hs__and2_2 _37724_ (.A(_06991_),
    .B(_06992_),
    .Y(_06993_));
 sky130_as_sc_hs__or2_2 _37726_ (.A(_06980_),
    .B(_06993_),
    .Y(_06995_));
 sky130_as_sc_hs__and2_2 _37727_ (.A(_06994_),
    .B(_06995_),
    .Y(_06996_));
 sky130_as_sc_hs__and2_2 _37730_ (.A(net444),
    .B(net432),
    .Y(_06999_));
 sky130_as_sc_hs__and2_2 _37731_ (.A(_24545_),
    .B(net435),
    .Y(_07000_));
 sky130_as_sc_hs__or2_2 _37732_ (.A(_06999_),
    .B(_07000_),
    .Y(_07001_));
 sky130_as_sc_hs__and2_2 _37734_ (.A(_07001_),
    .B(_07002_),
    .Y(_07003_));
 sky130_as_sc_hs__and2_2 _37735_ (.A(_24729_),
    .B(net428),
    .Y(_07004_));
 sky130_as_sc_hs__or2_2 _37737_ (.A(_07003_),
    .B(_07004_),
    .Y(_07006_));
 sky130_as_sc_hs__and2_2 _37738_ (.A(_07005_),
    .B(_07006_),
    .Y(_07007_));
 sky130_as_sc_hs__or2_2 _37740_ (.A(_06998_),
    .B(_07007_),
    .Y(_07009_));
 sky130_as_sc_hs__and2_2 _37741_ (.A(_07008_),
    .B(_07009_),
    .Y(_07010_));
 sky130_as_sc_hs__or2_2 _37743_ (.A(_06997_),
    .B(_07010_),
    .Y(_07012_));
 sky130_as_sc_hs__and2_2 _37744_ (.A(_07011_),
    .B(_07012_),
    .Y(_07013_));
 sky130_as_sc_hs__or2_2 _37747_ (.A(_07013_),
    .B(_07014_),
    .Y(_07016_));
 sky130_as_sc_hs__and2_2 _37748_ (.A(_07015_),
    .B(_07016_),
    .Y(_07017_));
 sky130_as_sc_hs__or2_2 _37750_ (.A(_06996_),
    .B(_07017_),
    .Y(_07019_));
 sky130_as_sc_hs__and2_2 _37751_ (.A(_07018_),
    .B(_07019_),
    .Y(_07020_));
 sky130_as_sc_hs__or2_2 _37753_ (.A(_06975_),
    .B(_07020_),
    .Y(_07022_));
 sky130_as_sc_hs__and2_2 _37754_ (.A(_07021_),
    .B(_07022_),
    .Y(_07023_));
 sky130_as_sc_hs__or2_2 _37756_ (.A(_06974_),
    .B(_07023_),
    .Y(_07025_));
 sky130_as_sc_hs__and2_2 _37757_ (.A(_07024_),
    .B(_07025_),
    .Y(_07026_));
 sky130_as_sc_hs__and2_2 _37760_ (.A(_23657_),
    .B(net449),
    .Y(_07029_));
 sky130_as_sc_hs__and2_2 _37761_ (.A(_24256_),
    .B(net426),
    .Y(_07030_));
 sky130_as_sc_hs__or2_2 _37762_ (.A(_07029_),
    .B(_07030_),
    .Y(_07031_));
 sky130_as_sc_hs__and2_2 _37764_ (.A(_07031_),
    .B(_07032_),
    .Y(_07033_));
 sky130_as_sc_hs__and2_2 _37765_ (.A(net451),
    .B(net84),
    .Y(_07034_));
 sky130_as_sc_hs__or2_2 _37767_ (.A(_07033_),
    .B(_07034_),
    .Y(_07036_));
 sky130_as_sc_hs__and2_2 _37768_ (.A(_07035_),
    .B(_07036_),
    .Y(_07037_));
 sky130_as_sc_hs__and2_2 _37769_ (.A(_24527_),
    .B(net438),
    .Y(_07038_));
 sky130_as_sc_hs__and2_2 _37770_ (.A(net472),
    .B(net89),
    .Y(_07039_));
 sky130_as_sc_hs__or2_2 _37771_ (.A(_07038_),
    .B(_07039_),
    .Y(_07040_));
 sky130_as_sc_hs__and2_2 _37773_ (.A(_07040_),
    .B(_07041_),
    .Y(_07042_));
 sky130_as_sc_hs__and2_2 _37774_ (.A(net479),
    .B(net88),
    .Y(_07043_));
 sky130_as_sc_hs__or2_2 _37776_ (.A(_07042_),
    .B(_07043_),
    .Y(_07045_));
 sky130_as_sc_hs__and2_2 _37777_ (.A(_07044_),
    .B(_07045_),
    .Y(_07046_));
 sky130_as_sc_hs__or2_2 _37780_ (.A(_07046_),
    .B(_07047_),
    .Y(_07049_));
 sky130_as_sc_hs__and2_2 _37781_ (.A(_07048_),
    .B(_07049_),
    .Y(_07050_));
 sky130_as_sc_hs__or2_2 _37783_ (.A(_07037_),
    .B(_07050_),
    .Y(_07052_));
 sky130_as_sc_hs__and2_2 _37784_ (.A(_07051_),
    .B(_07052_),
    .Y(_07053_));
 sky130_as_sc_hs__or2_2 _37786_ (.A(_07028_),
    .B(_07053_),
    .Y(_07055_));
 sky130_as_sc_hs__and2_2 _37787_ (.A(_07054_),
    .B(_07055_),
    .Y(_07056_));
 sky130_as_sc_hs__or2_2 _37789_ (.A(_07027_),
    .B(_07056_),
    .Y(_07058_));
 sky130_as_sc_hs__and2_2 _37790_ (.A(_07057_),
    .B(_07058_),
    .Y(_07059_));
 sky130_as_sc_hs__and2_2 _37793_ (.A(_23674_),
    .B(net465),
    .Y(_07062_));
 sky130_as_sc_hs__and2_2 _37794_ (.A(net480),
    .B(net463),
    .Y(_07063_));
 sky130_as_sc_hs__or2_2 _37795_ (.A(_07062_),
    .B(_07063_),
    .Y(_07064_));
 sky130_as_sc_hs__and2_2 _37797_ (.A(_07064_),
    .B(_07065_),
    .Y(_07066_));
 sky130_as_sc_hs__and2_2 _37798_ (.A(net476),
    .B(net460),
    .Y(_07067_));
 sky130_as_sc_hs__or2_2 _37800_ (.A(_07066_),
    .B(_07067_),
    .Y(_07069_));
 sky130_as_sc_hs__and2_2 _37801_ (.A(_07068_),
    .B(_07069_),
    .Y(_07070_));
 sky130_as_sc_hs__or2_2 _37803_ (.A(_07061_),
    .B(_07070_),
    .Y(_07072_));
 sky130_as_sc_hs__and2_2 _37804_ (.A(_07071_),
    .B(_07072_),
    .Y(_07073_));
 sky130_as_sc_hs__or2_2 _37806_ (.A(_07060_),
    .B(_07073_),
    .Y(_07075_));
 sky130_as_sc_hs__and2_2 _37807_ (.A(_07074_),
    .B(_07075_),
    .Y(_07076_));
 sky130_as_sc_hs__and2_2 _37808_ (.A(net467),
    .B(net446),
    .Y(_07077_));
 sky130_as_sc_hs__and2_2 _37809_ (.A(net469),
    .B(net78),
    .Y(_07078_));
 sky130_as_sc_hs__or2_2 _37810_ (.A(_07077_),
    .B(_07078_),
    .Y(_07079_));
 sky130_as_sc_hs__and2_2 _37812_ (.A(_07079_),
    .B(_07080_),
    .Y(_07081_));
 sky130_as_sc_hs__and2_2 _37813_ (.A(net470),
    .B(net442),
    .Y(_07082_));
 sky130_as_sc_hs__or2_2 _37815_ (.A(_07081_),
    .B(_07082_),
    .Y(_07084_));
 sky130_as_sc_hs__and2_2 _37816_ (.A(_07083_),
    .B(_07084_),
    .Y(_07085_));
 sky130_as_sc_hs__and2_2 _37817_ (.A(net456),
    .B(net454),
    .Y(_07086_));
 sky130_as_sc_hs__nand3_2 _37818_ (.A(_23598_),
    .B(_23712_),
    .C(_02549_),
    .Y(_07087_));
 sky130_as_sc_hs__nand3_2 _37819_ (.A(_24501_),
    .B(_25033_),
    .C(_25034_),
    .Y(_07088_));
 sky130_as_sc_hs__or2_2 _37821_ (.A(_07087_),
    .B(_07088_),
    .Y(_07090_));
 sky130_as_sc_hs__and2_2 _37822_ (.A(_07089_),
    .B(_07090_),
    .Y(_07091_));
 sky130_as_sc_hs__or2_2 _37824_ (.A(_07086_),
    .B(_07091_),
    .Y(_07093_));
 sky130_as_sc_hs__and2_2 _37825_ (.A(_07092_),
    .B(_07093_),
    .Y(_07094_));
 sky130_as_sc_hs__or2_2 _37828_ (.A(_07094_),
    .B(_07095_),
    .Y(_07097_));
 sky130_as_sc_hs__and2_2 _37829_ (.A(_07096_),
    .B(_07097_),
    .Y(_07098_));
 sky130_as_sc_hs__or2_2 _37831_ (.A(_07085_),
    .B(_07098_),
    .Y(_07100_));
 sky130_as_sc_hs__and2_2 _37832_ (.A(_07099_),
    .B(_07100_),
    .Y(_07101_));
 sky130_as_sc_hs__or2_2 _37835_ (.A(_07101_),
    .B(_07102_),
    .Y(_07104_));
 sky130_as_sc_hs__and2_2 _37836_ (.A(_07103_),
    .B(_07104_),
    .Y(_07105_));
 sky130_as_sc_hs__or2_2 _37838_ (.A(_07076_),
    .B(_07105_),
    .Y(_07107_));
 sky130_as_sc_hs__and2_2 _37839_ (.A(_07106_),
    .B(_07107_),
    .Y(_07108_));
 sky130_as_sc_hs__or2_2 _37842_ (.A(_07108_),
    .B(_07109_),
    .Y(_07111_));
 sky130_as_sc_hs__and2_2 _37843_ (.A(_07110_),
    .B(_07111_),
    .Y(_07112_));
 sky130_as_sc_hs__or2_2 _37845_ (.A(_07059_),
    .B(_07112_),
    .Y(_07114_));
 sky130_as_sc_hs__and2_2 _37846_ (.A(_07113_),
    .B(_07114_),
    .Y(_07115_));
 sky130_as_sc_hs__or2_2 _37849_ (.A(_07115_),
    .B(_07116_),
    .Y(_07118_));
 sky130_as_sc_hs__and2_2 _37850_ (.A(_07117_),
    .B(_07118_),
    .Y(_07119_));
 sky130_as_sc_hs__or2_2 _37852_ (.A(_07026_),
    .B(_07119_),
    .Y(_07121_));
 sky130_as_sc_hs__and2_2 _37853_ (.A(_07120_),
    .B(_07121_),
    .Y(_07122_));
 sky130_as_sc_hs__or2_2 _37856_ (.A(_07122_),
    .B(_07123_),
    .Y(_07125_));
 sky130_as_sc_hs__and2_2 _37857_ (.A(_07124_),
    .B(_07125_),
    .Y(_07126_));
 sky130_as_sc_hs__or2_2 _37859_ (.A(_06973_),
    .B(_07126_),
    .Y(_07128_));
 sky130_as_sc_hs__and2_2 _37860_ (.A(_07127_),
    .B(_07128_),
    .Y(_07129_));
 sky130_as_sc_hs__or2_2 _37863_ (.A(_07129_),
    .B(_07130_),
    .Y(_07132_));
 sky130_as_sc_hs__and2_2 _37864_ (.A(_07131_),
    .B(_07132_),
    .Y(_07133_));
 sky130_as_sc_hs__or2_2 _37866_ (.A(_06925_),
    .B(_07133_),
    .Y(_07135_));
 sky130_as_sc_hs__and2_2 _37867_ (.A(_07134_),
    .B(_07135_),
    .Y(_07136_));
 sky130_as_sc_hs__or2_2 _37870_ (.A(_07136_),
    .B(_07137_),
    .Y(_07139_));
 sky130_as_sc_hs__and2_2 _37871_ (.A(_07138_),
    .B(_07139_),
    .Y(_07140_));
 sky130_as_sc_hs__or2_2 _37873_ (.A(_06924_),
    .B(_07140_),
    .Y(_07142_));
 sky130_as_sc_hs__and2_2 _37874_ (.A(_07141_),
    .B(_07142_),
    .Y(_07143_));
 sky130_as_sc_hs__or2_2 _37876_ (.A(_06923_),
    .B(_07143_),
    .Y(_07145_));
 sky130_as_sc_hs__and2_2 _37877_ (.A(_07144_),
    .B(_07145_),
    .Y(_07146_));
 sky130_as_sc_hs__or2_2 _37879_ (.A(_07146_),
    .B(_07147_),
    .Y(_07148_));
 sky130_as_sc_hs__nor2b_2 _37882_ (.A(_06822_),
    .Y(_07151_),
    .B(_06821_));
 sky130_as_sc_hs__or2_2 _37886_ (.A(_07150_),
    .B(_07153_),
    .Y(_07155_));
 sky130_as_sc_hs__nand3_2 _37887_ (.A(net142),
    .B(_07154_),
    .C(_07155_),
    .Y(_07156_));
 sky130_as_sc_hs__nor2_2 _37888_ (.A(_04515_),
    .B(_04517_),
    .Y(_07157_));
 sky130_as_sc_hs__or2_2 _37889_ (.A(_04518_),
    .B(_07157_),
    .Y(_07158_));
 sky130_as_sc_hs__or2_2 _37890_ (.A(_05400_),
    .B(_05505_),
    .Y(_07159_));
 sky130_as_sc_hs__or2_2 _37892_ (.A(_07158_),
    .B(_07159_),
    .Y(_07161_));
 sky130_as_sc_hs__nand3_2 _37893_ (.A(net139),
    .B(_07160_),
    .C(_07161_),
    .Y(_07162_));
 sky130_as_sc_hs__or2_2 _37894_ (.A(_05810_),
    .B(_05851_),
    .Y(_07163_));
 sky130_as_sc_hs__nand3_2 _37895_ (.A(_05852_),
    .B(_06527_),
    .C(_07163_),
    .Y(_07164_));
 sky130_as_sc_hs__nor2_2 _37896_ (.A(_05823_),
    .B(_06870_),
    .Y(_07165_));
 sky130_as_sc_hs__nor2_2 _37897_ (.A(_05822_),
    .B(_07165_),
    .Y(_07166_));
 sky130_as_sc_hs__or2_2 _37898_ (.A(_05810_),
    .B(_07166_),
    .Y(_07167_));
 sky130_as_sc_hs__or2_2 _37901_ (.A(_06527_),
    .B(_07169_),
    .Y(_07170_));
 sky130_as_sc_hs__and2_2 _37903_ (.A(net119),
    .B(_07171_),
    .Y(_07172_));
 sky130_as_sc_hs__or2_2 _37907_ (.A(\tholin_riscv.div_res[2] ),
    .B(_06880_),
    .Y(_07176_));
 sky130_as_sc_hs__and2_2 _37908_ (.A(net415),
    .B(_07176_),
    .Y(_07177_));
 sky130_as_sc_hs__or2_2 _37910_ (.A(\tholin_riscv.div_res[3] ),
    .B(_07177_),
    .Y(_07179_));
 sky130_as_sc_hs__nand3_2 _37911_ (.A(net111),
    .B(_07178_),
    .C(_07179_),
    .Y(_07180_));
 sky130_as_sc_hs__nor2_2 _37912_ (.A(_05807_),
    .B(_06161_),
    .Y(_07181_));
 sky130_as_sc_hs__or2_2 _37913_ (.A(\tholin_riscv.div_shifter[34] ),
    .B(_06886_),
    .Y(_07182_));
 sky130_as_sc_hs__and2_2 _37914_ (.A(_21655_),
    .B(_07182_),
    .Y(_07183_));
 sky130_as_sc_hs__or2_2 _37916_ (.A(\tholin_riscv.div_shifter[35] ),
    .B(_07183_),
    .Y(_07185_));
 sky130_as_sc_hs__nand3_2 _37917_ (.A(net109),
    .B(_07184_),
    .C(_07185_),
    .Y(_07186_));
 sky130_as_sc_hs__and2_2 _37920_ (.A(_07187_),
    .B(_07188_),
    .Y(_07189_));
 sky130_as_sc_hs__nand3_2 _37921_ (.A(net413),
    .B(_07186_),
    .C(_07189_),
    .Y(_07190_));
 sky130_as_sc_hs__nor2_2 _37922_ (.A(_07181_),
    .B(_07190_),
    .Y(_07191_));
 sky130_as_sc_hs__nand3_2 _37923_ (.A(_07175_),
    .B(_07180_),
    .C(_07191_),
    .Y(_07192_));
 sky130_as_sc_hs__nor2_2 _37924_ (.A(_07172_),
    .B(_07192_),
    .Y(_07193_));
 sky130_as_sc_hs__and2_2 _37925_ (.A(_05946_),
    .B(_06466_),
    .Y(_07194_));
 sky130_as_sc_hs__and2_2 _37926_ (.A(_05945_),
    .B(_06503_),
    .Y(_07195_));
 sky130_as_sc_hs__nor2_2 _37927_ (.A(_07194_),
    .B(_07195_),
    .Y(_07196_));
 sky130_as_sc_hs__or2_2 _37934_ (.A(_05935_),
    .B(_07202_),
    .Y(_07203_));
 sky130_as_sc_hs__or2_2 _37936_ (.A(net82),
    .B(_06440_),
    .Y(_07205_));
 sky130_as_sc_hs__or2_2 _37937_ (.A(net82),
    .B(_06444_),
    .Y(_07206_));
 sky130_as_sc_hs__and2_2 _37939_ (.A(_07206_),
    .B(_07207_),
    .Y(_07208_));
 sky130_as_sc_hs__nand3_2 _37941_ (.A(_05941_),
    .B(_07204_),
    .C(_07205_),
    .Y(_07210_));
 sky130_as_sc_hs__nand3_2 _37942_ (.A(_05935_),
    .B(_07209_),
    .C(_07210_),
    .Y(_07211_));
 sky130_as_sc_hs__and2_2 _37944_ (.A(_05945_),
    .B(_06491_),
    .Y(_07213_));
 sky130_as_sc_hs__and2_2 _37945_ (.A(_05946_),
    .B(_06480_),
    .Y(_07214_));
 sky130_as_sc_hs__nor2_2 _37946_ (.A(_07213_),
    .B(_07214_),
    .Y(_07215_));
 sky130_as_sc_hs__and2_2 _37948_ (.A(_07212_),
    .B(_07216_),
    .Y(_07217_));
 sky130_as_sc_hs__or2_2 _37949_ (.A(_05935_),
    .B(_07217_),
    .Y(_07218_));
 sky130_as_sc_hs__and2_2 _37960_ (.A(_07218_),
    .B(_07228_),
    .Y(_07229_));
 sky130_as_sc_hs__nand3_2 _37961_ (.A(_05929_),
    .B(_07203_),
    .C(_07211_),
    .Y(_07230_));
 sky130_as_sc_hs__or2_2 _37962_ (.A(_05929_),
    .B(_07229_),
    .Y(_07231_));
 sky130_as_sc_hs__and2_2 _37963_ (.A(_07230_),
    .B(_07231_),
    .Y(_07232_));
 sky130_as_sc_hs__and2_2 _37972_ (.A(_07193_),
    .B(_07233_),
    .Y(_07241_));
 sky130_as_sc_hs__and2_2 _37973_ (.A(_07240_),
    .B(_07241_),
    .Y(_07242_));
 sky130_as_sc_hs__nand3_2 _37974_ (.A(_07156_),
    .B(_07162_),
    .C(_07242_),
    .Y(_07243_));
 sky130_as_sc_hs__and2_2 _37975_ (.A(\tholin_riscv.PC[3] ),
    .B(\tholin_riscv.PC[2] ),
    .Y(_07244_));
 sky130_as_sc_hs__nor2_2 _37976_ (.A(\tholin_riscv.PC[3] ),
    .B(\tholin_riscv.PC[2] ),
    .Y(_07245_));
 sky130_as_sc_hs__nor2_2 _37977_ (.A(_07244_),
    .B(_07245_),
    .Y(_07246_));
 sky130_as_sc_hs__inv_2 _37978_ (.Y(_07247_),
    .A(_07246_));
 sky130_as_sc_hs__nand3_2 _37981_ (.A(_21569_),
    .B(_07248_),
    .C(_07249_),
    .Y(_07250_));
 sky130_as_sc_hs__nand3_2 _37982_ (.A(_21546_),
    .B(_07243_),
    .C(_07250_),
    .Y(_07251_));
 sky130_as_sc_hs__and2_2 _37993_ (.A(_23636_),
    .B(net420),
    .Y(_07261_));
 sky130_as_sc_hs__and2_2 _37994_ (.A(_24256_),
    .B(net422),
    .Y(_07262_));
 sky130_as_sc_hs__or2_2 _37995_ (.A(_07261_),
    .B(_07262_),
    .Y(_07263_));
 sky130_as_sc_hs__and2_2 _37997_ (.A(_07263_),
    .B(_07264_),
    .Y(_07265_));
 sky130_as_sc_hs__and2_2 _37998_ (.A(net482),
    .B(net428),
    .Y(_07266_));
 sky130_as_sc_hs__or2_2 _38000_ (.A(_07265_),
    .B(_07266_),
    .Y(_07268_));
 sky130_as_sc_hs__and2_2 _38001_ (.A(_07267_),
    .B(_07268_),
    .Y(_07269_));
 sky130_as_sc_hs__or2_2 _38004_ (.A(_07269_),
    .B(_07270_),
    .Y(_07272_));
 sky130_as_sc_hs__or2_2 _38006_ (.A(_06938_),
    .B(_07273_),
    .Y(_07274_));
 sky130_as_sc_hs__and2_2 _38008_ (.A(_07274_),
    .B(_07275_),
    .Y(_07276_));
 sky130_as_sc_hs__and2_2 _38009_ (.A(net123),
    .B(_23702_),
    .Y(_07277_));
 sky130_as_sc_hs__or2_2 _38011_ (.A(_07276_),
    .B(_07277_),
    .Y(_07279_));
 sky130_as_sc_hs__and2_2 _38012_ (.A(_07278_),
    .B(_07279_),
    .Y(_07280_));
 sky130_as_sc_hs__and2_2 _38014_ (.A(_24229_),
    .B(net129),
    .Y(_07282_));
 sky130_as_sc_hs__or2_2 _38016_ (.A(_06978_),
    .B(_07282_),
    .Y(_07284_));
 sky130_as_sc_hs__and2_2 _38017_ (.A(_07283_),
    .B(_07284_),
    .Y(_07285_));
 sky130_as_sc_hs__or2_2 _38019_ (.A(_07281_),
    .B(_07285_),
    .Y(_07287_));
 sky130_as_sc_hs__or2_2 _38021_ (.A(_06952_),
    .B(_07288_),
    .Y(_07289_));
 sky130_as_sc_hs__and2_2 _38023_ (.A(_07289_),
    .B(_07290_),
    .Y(_07291_));
 sky130_as_sc_hs__or2_2 _38026_ (.A(_07291_),
    .B(_07292_),
    .Y(_07294_));
 sky130_as_sc_hs__and2_2 _38027_ (.A(_07293_),
    .B(_07294_),
    .Y(_07295_));
 sky130_as_sc_hs__or2_2 _38029_ (.A(_07280_),
    .B(_07295_),
    .Y(_07297_));
 sky130_as_sc_hs__and2_2 _38030_ (.A(_07296_),
    .B(_07297_),
    .Y(_07298_));
 sky130_as_sc_hs__or2_2 _38032_ (.A(_07260_),
    .B(_07298_),
    .Y(_07300_));
 sky130_as_sc_hs__and2_2 _38033_ (.A(_07299_),
    .B(_07300_),
    .Y(_07301_));
 sky130_as_sc_hs__or2_2 _38035_ (.A(_07259_),
    .B(_07301_),
    .Y(_07303_));
 sky130_as_sc_hs__and2_2 _38036_ (.A(_07302_),
    .B(_07303_),
    .Y(_07304_));
 sky130_as_sc_hs__and2_2 _38039_ (.A(_24774_),
    .B(net424),
    .Y(_07307_));
 sky130_as_sc_hs__and2_2 _38040_ (.A(net452),
    .B(net441),
    .Y(_07308_));
 sky130_as_sc_hs__or2_2 _38041_ (.A(_07307_),
    .B(_07308_),
    .Y(_07309_));
 sky130_as_sc_hs__and2_2 _38043_ (.A(_07309_),
    .B(_07310_),
    .Y(_07311_));
 sky130_as_sc_hs__and2_2 _38044_ (.A(_24768_),
    .B(net75),
    .Y(_07312_));
 sky130_as_sc_hs__or2_2 _38046_ (.A(_07311_),
    .B(_07312_),
    .Y(_07314_));
 sky130_as_sc_hs__and2_2 _38047_ (.A(_07313_),
    .B(_07314_),
    .Y(_07315_));
 sky130_as_sc_hs__or2_2 _38050_ (.A(_07315_),
    .B(_07316_),
    .Y(_07318_));
 sky130_as_sc_hs__and2_2 _38051_ (.A(_07317_),
    .B(_07318_),
    .Y(_07319_));
 sky130_as_sc_hs__and2_2 _38052_ (.A(net447),
    .B(net436),
    .Y(_07320_));
 sky130_as_sc_hs__or2_2 _38054_ (.A(_07319_),
    .B(_07320_),
    .Y(_07322_));
 sky130_as_sc_hs__and2_2 _38055_ (.A(_07321_),
    .B(_07322_),
    .Y(_07323_));
 sky130_as_sc_hs__and2_2 _38058_ (.A(net444),
    .B(net429),
    .Y(_07326_));
 sky130_as_sc_hs__and2_2 _38059_ (.A(net454),
    .B(net434),
    .Y(_07327_));
 sky130_as_sc_hs__or2_2 _38060_ (.A(_07326_),
    .B(_07327_),
    .Y(_07328_));
 sky130_as_sc_hs__and2_2 _38062_ (.A(_07328_),
    .B(_07329_),
    .Y(_07330_));
 sky130_as_sc_hs__and2_2 _38063_ (.A(net120),
    .B(_24729_),
    .Y(_07331_));
 sky130_as_sc_hs__or2_2 _38065_ (.A(_07330_),
    .B(_07331_),
    .Y(_07333_));
 sky130_as_sc_hs__and2_2 _38066_ (.A(_07332_),
    .B(_07333_),
    .Y(_07334_));
 sky130_as_sc_hs__or2_2 _38068_ (.A(_07325_),
    .B(_07334_),
    .Y(_07336_));
 sky130_as_sc_hs__and2_2 _38069_ (.A(_07335_),
    .B(_07336_),
    .Y(_07337_));
 sky130_as_sc_hs__or2_2 _38071_ (.A(_07324_),
    .B(_07337_),
    .Y(_07339_));
 sky130_as_sc_hs__and2_2 _38072_ (.A(_07338_),
    .B(_07339_),
    .Y(_07340_));
 sky130_as_sc_hs__or2_2 _38075_ (.A(_07340_),
    .B(_07341_),
    .Y(_07343_));
 sky130_as_sc_hs__and2_2 _38076_ (.A(_07342_),
    .B(_07343_),
    .Y(_07344_));
 sky130_as_sc_hs__or2_2 _38078_ (.A(_07323_),
    .B(_07344_),
    .Y(_07346_));
 sky130_as_sc_hs__and2_2 _38079_ (.A(_07345_),
    .B(_07346_),
    .Y(_07347_));
 sky130_as_sc_hs__or2_2 _38081_ (.A(_07306_),
    .B(_07347_),
    .Y(_07349_));
 sky130_as_sc_hs__and2_2 _38082_ (.A(_07348_),
    .B(_07349_),
    .Y(_07350_));
 sky130_as_sc_hs__or2_2 _38084_ (.A(_07305_),
    .B(_07350_),
    .Y(_07352_));
 sky130_as_sc_hs__and2_2 _38085_ (.A(_07351_),
    .B(_07352_),
    .Y(_07353_));
 sky130_as_sc_hs__and2_2 _38088_ (.A(net449),
    .B(net83),
    .Y(_07356_));
 sky130_as_sc_hs__and2_2 _38089_ (.A(_24501_),
    .B(net426),
    .Y(_07357_));
 sky130_as_sc_hs__or2_2 _38090_ (.A(_07356_),
    .B(_07357_),
    .Y(_07358_));
 sky130_as_sc_hs__and2_2 _38092_ (.A(_07358_),
    .B(_07359_),
    .Y(_07360_));
 sky130_as_sc_hs__and2_2 _38093_ (.A(net451),
    .B(net431),
    .Y(_07361_));
 sky130_as_sc_hs__or2_2 _38095_ (.A(_07360_),
    .B(_07361_),
    .Y(_07363_));
 sky130_as_sc_hs__and2_2 _38096_ (.A(_07362_),
    .B(_07363_),
    .Y(_07364_));
 sky130_as_sc_hs__and2_2 _38097_ (.A(net472),
    .B(_24527_),
    .Y(_07365_));
 sky130_as_sc_hs__and2_2 _38098_ (.A(net478),
    .B(net89),
    .Y(_07366_));
 sky130_as_sc_hs__or2_2 _38099_ (.A(_07365_),
    .B(_07366_),
    .Y(_07367_));
 sky130_as_sc_hs__and2_2 _38101_ (.A(_07367_),
    .B(_07368_),
    .Y(_07369_));
 sky130_as_sc_hs__and2_2 _38102_ (.A(net474),
    .B(net88),
    .Y(_07370_));
 sky130_as_sc_hs__or2_2 _38104_ (.A(_07369_),
    .B(_07370_),
    .Y(_07372_));
 sky130_as_sc_hs__and2_2 _38105_ (.A(_07371_),
    .B(_07372_),
    .Y(_07373_));
 sky130_as_sc_hs__or2_2 _38108_ (.A(_07373_),
    .B(_07374_),
    .Y(_07376_));
 sky130_as_sc_hs__and2_2 _38109_ (.A(_07375_),
    .B(_07376_),
    .Y(_07377_));
 sky130_as_sc_hs__or2_2 _38111_ (.A(_07364_),
    .B(_07377_),
    .Y(_07379_));
 sky130_as_sc_hs__and2_2 _38112_ (.A(_07378_),
    .B(_07379_),
    .Y(_07380_));
 sky130_as_sc_hs__or2_2 _38114_ (.A(_07355_),
    .B(_07380_),
    .Y(_07382_));
 sky130_as_sc_hs__and2_2 _38115_ (.A(_07381_),
    .B(_07382_),
    .Y(_07383_));
 sky130_as_sc_hs__or2_2 _38117_ (.A(_07354_),
    .B(_07383_),
    .Y(_07385_));
 sky130_as_sc_hs__and2_2 _38118_ (.A(_07384_),
    .B(_07385_),
    .Y(_07386_));
 sky130_as_sc_hs__and2_2 _38121_ (.A(net480),
    .B(net465),
    .Y(_07389_));
 sky130_as_sc_hs__and2_2 _38122_ (.A(net476),
    .B(net463),
    .Y(_07390_));
 sky130_as_sc_hs__or2_2 _38123_ (.A(_07389_),
    .B(_07390_),
    .Y(_07391_));
 sky130_as_sc_hs__and2_2 _38125_ (.A(_07391_),
    .B(_07392_),
    .Y(_07393_));
 sky130_as_sc_hs__and2_2 _38126_ (.A(net460),
    .B(net438),
    .Y(_07394_));
 sky130_as_sc_hs__or2_2 _38128_ (.A(_07393_),
    .B(_07394_),
    .Y(_07396_));
 sky130_as_sc_hs__and2_2 _38129_ (.A(_07395_),
    .B(_07396_),
    .Y(_07397_));
 sky130_as_sc_hs__or2_2 _38131_ (.A(_07388_),
    .B(_07397_),
    .Y(_07399_));
 sky130_as_sc_hs__and2_2 _38132_ (.A(_07398_),
    .B(_07399_),
    .Y(_07400_));
 sky130_as_sc_hs__or2_2 _38134_ (.A(_07387_),
    .B(_07400_),
    .Y(_07402_));
 sky130_as_sc_hs__and2_2 _38135_ (.A(_07401_),
    .B(_07402_),
    .Y(_07403_));
 sky130_as_sc_hs__and2_2 _38136_ (.A(net467),
    .B(net78),
    .Y(_07404_));
 sky130_as_sc_hs__and2_2 _38137_ (.A(net469),
    .B(net442),
    .Y(_07405_));
 sky130_as_sc_hs__or2_2 _38138_ (.A(_07404_),
    .B(_07405_),
    .Y(_07406_));
 sky130_as_sc_hs__and2_2 _38140_ (.A(_07406_),
    .B(_07407_),
    .Y(_07408_));
 sky130_as_sc_hs__and2_2 _38141_ (.A(_23674_),
    .B(net471),
    .Y(_07409_));
 sky130_as_sc_hs__or2_2 _38143_ (.A(_07408_),
    .B(_07409_),
    .Y(_07411_));
 sky130_as_sc_hs__and2_2 _38144_ (.A(_07410_),
    .B(_07411_),
    .Y(_07412_));
 sky130_as_sc_hs__and2_2 _38145_ (.A(net456),
    .B(net85),
    .Y(_07413_));
 sky130_as_sc_hs__or2_2 _38149_ (.A(_07414_),
    .B(_07415_),
    .Y(_07417_));
 sky130_as_sc_hs__and2_2 _38150_ (.A(_07416_),
    .B(_07417_),
    .Y(_07418_));
 sky130_as_sc_hs__or2_2 _38152_ (.A(_07413_),
    .B(_07418_),
    .Y(_07420_));
 sky130_as_sc_hs__and2_2 _38153_ (.A(_07419_),
    .B(_07420_),
    .Y(_07421_));
 sky130_as_sc_hs__or2_2 _38156_ (.A(_07421_),
    .B(_07422_),
    .Y(_07424_));
 sky130_as_sc_hs__and2_2 _38157_ (.A(_07423_),
    .B(_07424_),
    .Y(_07425_));
 sky130_as_sc_hs__or2_2 _38159_ (.A(_07412_),
    .B(_07425_),
    .Y(_07427_));
 sky130_as_sc_hs__and2_2 _38160_ (.A(_07426_),
    .B(_07427_),
    .Y(_07428_));
 sky130_as_sc_hs__or2_2 _38163_ (.A(_07428_),
    .B(_07429_),
    .Y(_07431_));
 sky130_as_sc_hs__and2_2 _38164_ (.A(_07430_),
    .B(_07431_),
    .Y(_07432_));
 sky130_as_sc_hs__or2_2 _38166_ (.A(_07403_),
    .B(_07432_),
    .Y(_07434_));
 sky130_as_sc_hs__and2_2 _38167_ (.A(_07433_),
    .B(_07434_),
    .Y(_07435_));
 sky130_as_sc_hs__or2_2 _38170_ (.A(_07435_),
    .B(_07436_),
    .Y(_07438_));
 sky130_as_sc_hs__and2_2 _38171_ (.A(_07437_),
    .B(_07438_),
    .Y(_07439_));
 sky130_as_sc_hs__or2_2 _38173_ (.A(_07386_),
    .B(_07439_),
    .Y(_07441_));
 sky130_as_sc_hs__and2_2 _38174_ (.A(_07440_),
    .B(_07441_),
    .Y(_07442_));
 sky130_as_sc_hs__or2_2 _38177_ (.A(_07442_),
    .B(_07443_),
    .Y(_07445_));
 sky130_as_sc_hs__and2_2 _38178_ (.A(_07444_),
    .B(_07445_),
    .Y(_07446_));
 sky130_as_sc_hs__or2_2 _38180_ (.A(_07353_),
    .B(_07446_),
    .Y(_07448_));
 sky130_as_sc_hs__and2_2 _38181_ (.A(_07447_),
    .B(_07448_),
    .Y(_07449_));
 sky130_as_sc_hs__or2_2 _38184_ (.A(_07449_),
    .B(_07450_),
    .Y(_07452_));
 sky130_as_sc_hs__and2_2 _38185_ (.A(_07451_),
    .B(_07452_),
    .Y(_07453_));
 sky130_as_sc_hs__or2_2 _38187_ (.A(_07304_),
    .B(_07453_),
    .Y(_07455_));
 sky130_as_sc_hs__and2_2 _38188_ (.A(_07454_),
    .B(_07455_),
    .Y(_07456_));
 sky130_as_sc_hs__or2_2 _38191_ (.A(_07456_),
    .B(_07457_),
    .Y(_07459_));
 sky130_as_sc_hs__and2_2 _38192_ (.A(_07458_),
    .B(_07459_),
    .Y(_07460_));
 sky130_as_sc_hs__or2_2 _38194_ (.A(_07258_),
    .B(_07460_),
    .Y(_07462_));
 sky130_as_sc_hs__and2_2 _38195_ (.A(_07461_),
    .B(_07462_),
    .Y(_07463_));
 sky130_as_sc_hs__or2_2 _38198_ (.A(_07463_),
    .B(_07464_),
    .Y(_07466_));
 sky130_as_sc_hs__and2_2 _38199_ (.A(_07465_),
    .B(_07466_),
    .Y(_07467_));
 sky130_as_sc_hs__nand3_2 _38200_ (.A(_07257_),
    .B(_07465_),
    .C(_07466_),
    .Y(_07468_));
 sky130_as_sc_hs__or2_2 _38201_ (.A(_07257_),
    .B(_07467_),
    .Y(_07469_));
 sky130_as_sc_hs__and2_2 _38202_ (.A(_07468_),
    .B(_07469_),
    .Y(_07470_));
 sky130_as_sc_hs__nand3_2 _38204_ (.A(_07468_),
    .B(_07469_),
    .C(_07471_),
    .Y(_07472_));
 sky130_as_sc_hs__or2_2 _38205_ (.A(_07470_),
    .B(_07471_),
    .Y(_07473_));
 sky130_as_sc_hs__and2_2 _38206_ (.A(_07472_),
    .B(_07473_),
    .Y(_07474_));
 sky130_as_sc_hs__and2_2 _38207_ (.A(_06813_),
    .B(_07146_),
    .Y(_07475_));
 sky130_as_sc_hs__nand2b_2 _38208_ (.B(_07475_),
    .Y(_07476_),
    .A(_06815_));
 sky130_as_sc_hs__and2_2 _38211_ (.A(_07476_),
    .B(_07478_),
    .Y(_07479_));
 sky130_as_sc_hs__and2_2 _38212_ (.A(_06816_),
    .B(_07475_),
    .Y(_07480_));
 sky130_as_sc_hs__and2_2 _38215_ (.A(_07474_),
    .B(_07482_),
    .Y(_07483_));
 sky130_as_sc_hs__nor2_2 _38217_ (.A(_07474_),
    .B(_07482_),
    .Y(_07485_));
 sky130_as_sc_hs__or2_2 _38218_ (.A(_07483_),
    .B(_07485_),
    .Y(_07486_));
 sky130_as_sc_hs__nand3_2 _38219_ (.A(_05501_),
    .B(_07150_),
    .C(_07151_),
    .Y(_07487_));
 sky130_as_sc_hs__or2_2 _38222_ (.A(_07486_),
    .B(_07488_),
    .Y(_07490_));
 sky130_as_sc_hs__nand3_2 _38223_ (.A(net142),
    .B(_07489_),
    .C(_07490_),
    .Y(_07491_));
 sky130_as_sc_hs__nor2_2 _38224_ (.A(_04518_),
    .B(_04520_),
    .Y(_07492_));
 sky130_as_sc_hs__nor2_2 _38225_ (.A(_04521_),
    .B(_07492_),
    .Y(_07493_));
 sky130_as_sc_hs__nor2_2 _38226_ (.A(_05401_),
    .B(_05505_),
    .Y(_07494_));
 sky130_as_sc_hs__or2_2 _38228_ (.A(_07493_),
    .B(_07494_),
    .Y(_07496_));
 sky130_as_sc_hs__nand3_2 _38229_ (.A(net139),
    .B(_07495_),
    .C(_07496_),
    .Y(_07497_));
 sky130_as_sc_hs__or2_2 _38230_ (.A(_05795_),
    .B(_05853_),
    .Y(_07498_));
 sky130_as_sc_hs__or2_2 _38231_ (.A(_05808_),
    .B(_07166_),
    .Y(_07499_));
 sky130_as_sc_hs__and2_2 _38232_ (.A(_05807_),
    .B(_07499_),
    .Y(_07500_));
 sky130_as_sc_hs__or2_2 _38233_ (.A(_05795_),
    .B(_07500_),
    .Y(_07501_));
 sky130_as_sc_hs__nand3_2 _38239_ (.A(net119),
    .B(_07504_),
    .C(_07506_),
    .Y(_07507_));
 sky130_as_sc_hs__or2_2 _38240_ (.A(_05941_),
    .B(_06031_),
    .Y(_07508_));
 sky130_as_sc_hs__nand3_2 _38242_ (.A(_05935_),
    .B(_07508_),
    .C(_07509_),
    .Y(_07510_));
 sky130_as_sc_hs__or2_2 _38246_ (.A(_05935_),
    .B(_07513_),
    .Y(_07514_));
 sky130_as_sc_hs__and2_2 _38249_ (.A(_07515_),
    .B(_07516_),
    .Y(_07517_));
 sky130_as_sc_hs__or2_2 _38251_ (.A(_05935_),
    .B(_07235_),
    .Y(_07519_));
 sky130_as_sc_hs__and2_2 _38252_ (.A(_07518_),
    .B(_07519_),
    .Y(_07520_));
 sky130_as_sc_hs__nand3_2 _38253_ (.A(_05929_),
    .B(_07510_),
    .C(_07514_),
    .Y(_07521_));
 sky130_as_sc_hs__and2_2 _38261_ (.A(net140),
    .B(_07528_),
    .Y(_07529_));
 sky130_as_sc_hs__or2_2 _38265_ (.A(\tholin_riscv.div_res[3] ),
    .B(_07176_),
    .Y(_07533_));
 sky130_as_sc_hs__and2_2 _38266_ (.A(net415),
    .B(_07533_),
    .Y(_07534_));
 sky130_as_sc_hs__or2_2 _38268_ (.A(\tholin_riscv.div_res[4] ),
    .B(_07534_),
    .Y(_07536_));
 sky130_as_sc_hs__nand3_2 _38269_ (.A(net111),
    .B(_07535_),
    .C(_07536_),
    .Y(_07537_));
 sky130_as_sc_hs__nor2_2 _38270_ (.A(_05792_),
    .B(_06161_),
    .Y(_07538_));
 sky130_as_sc_hs__or2_2 _38271_ (.A(\tholin_riscv.div_shifter[35] ),
    .B(_07182_),
    .Y(_07539_));
 sky130_as_sc_hs__and2_2 _38272_ (.A(_21655_),
    .B(_07539_),
    .Y(_07540_));
 sky130_as_sc_hs__or2_2 _38274_ (.A(\tholin_riscv.div_shifter[36] ),
    .B(_07540_),
    .Y(_07542_));
 sky130_as_sc_hs__nand3_2 _38275_ (.A(net109),
    .B(_07541_),
    .C(_07542_),
    .Y(_07543_));
 sky130_as_sc_hs__and2_2 _38278_ (.A(_07544_),
    .B(_07545_),
    .Y(_07546_));
 sky130_as_sc_hs__nand3_2 _38279_ (.A(net412),
    .B(_07543_),
    .C(_07546_),
    .Y(_07547_));
 sky130_as_sc_hs__nor2_2 _38280_ (.A(_07538_),
    .B(_07547_),
    .Y(_07548_));
 sky130_as_sc_hs__nand3_2 _38281_ (.A(_07532_),
    .B(_07537_),
    .C(_07548_),
    .Y(_07549_));
 sky130_as_sc_hs__nor2_2 _38282_ (.A(_07529_),
    .B(_07549_),
    .Y(_07550_));
 sky130_as_sc_hs__and2_2 _38283_ (.A(_07524_),
    .B(_07550_),
    .Y(_07551_));
 sky130_as_sc_hs__and2_2 _38284_ (.A(_07507_),
    .B(_07551_),
    .Y(_07552_));
 sky130_as_sc_hs__nand3_2 _38285_ (.A(_07491_),
    .B(_07497_),
    .C(_07552_),
    .Y(_07553_));
 sky130_as_sc_hs__and2_2 _38286_ (.A(\tholin_riscv.PC[4] ),
    .B(_07244_),
    .Y(_07554_));
 sky130_as_sc_hs__nor2_2 _38287_ (.A(\tholin_riscv.PC[4] ),
    .B(_07244_),
    .Y(_07555_));
 sky130_as_sc_hs__nor2_2 _38288_ (.A(_07554_),
    .B(_07555_),
    .Y(_07556_));
 sky130_as_sc_hs__inv_2 _38289_ (.Y(_07557_),
    .A(_07556_));
 sky130_as_sc_hs__nand3_2 _38292_ (.A(_21569_),
    .B(_07558_),
    .C(_07559_),
    .Y(_07560_));
 sky130_as_sc_hs__nand3_2 _38293_ (.A(_21546_),
    .B(_07553_),
    .C(_07560_),
    .Y(_07561_));
 sky130_as_sc_hs__and2_2 _38302_ (.A(_23636_),
    .B(net75),
    .Y(_07569_));
 sky130_as_sc_hs__and2_2 _38303_ (.A(_24501_),
    .B(net422),
    .Y(_07570_));
 sky130_as_sc_hs__or2_2 _38304_ (.A(_07569_),
    .B(_07570_),
    .Y(_07571_));
 sky130_as_sc_hs__and2_2 _38306_ (.A(_07571_),
    .B(_07572_),
    .Y(_07573_));
 sky130_as_sc_hs__and2_2 _38307_ (.A(net482),
    .B(net121),
    .Y(_07574_));
 sky130_as_sc_hs__or2_2 _38309_ (.A(_07573_),
    .B(_07574_),
    .Y(_07576_));
 sky130_as_sc_hs__and2_2 _38310_ (.A(_07575_),
    .B(_07576_),
    .Y(_07577_));
 sky130_as_sc_hs__or2_2 _38313_ (.A(_07577_),
    .B(_07578_),
    .Y(_07580_));
 sky130_as_sc_hs__or2_2 _38315_ (.A(_07271_),
    .B(_07581_),
    .Y(_07582_));
 sky130_as_sc_hs__and2_2 _38317_ (.A(_07582_),
    .B(_07583_),
    .Y(_07584_));
 sky130_as_sc_hs__and2_2 _38318_ (.A(_23702_),
    .B(net424),
    .Y(_07585_));
 sky130_as_sc_hs__or2_2 _38320_ (.A(_07584_),
    .B(_07585_),
    .Y(_07587_));
 sky130_as_sc_hs__and2_2 _38321_ (.A(_07586_),
    .B(_07587_),
    .Y(_07588_));
 sky130_as_sc_hs__and2_2 _38323_ (.A(_24256_),
    .B(net129),
    .Y(_07590_));
 sky130_as_sc_hs__or2_2 _38325_ (.A(_07589_),
    .B(_07590_),
    .Y(_07592_));
 sky130_as_sc_hs__or2_2 _38327_ (.A(_07283_),
    .B(_07593_),
    .Y(_07594_));
 sky130_as_sc_hs__and2_2 _38329_ (.A(_07594_),
    .B(_07595_),
    .Y(_07596_));
 sky130_as_sc_hs__or2_2 _38332_ (.A(_07596_),
    .B(_07597_),
    .Y(_07599_));
 sky130_as_sc_hs__and2_2 _38333_ (.A(_07598_),
    .B(_07599_),
    .Y(_07600_));
 sky130_as_sc_hs__or2_2 _38335_ (.A(_07588_),
    .B(_07600_),
    .Y(_07602_));
 sky130_as_sc_hs__and2_2 _38336_ (.A(_07601_),
    .B(_07602_),
    .Y(_07603_));
 sky130_as_sc_hs__or2_2 _38338_ (.A(_07568_),
    .B(_07603_),
    .Y(_07605_));
 sky130_as_sc_hs__and2_2 _38339_ (.A(_07604_),
    .B(_07605_),
    .Y(_07606_));
 sky130_as_sc_hs__or2_2 _38341_ (.A(_07567_),
    .B(_07606_),
    .Y(_07608_));
 sky130_as_sc_hs__and2_2 _38342_ (.A(_07607_),
    .B(_07608_),
    .Y(_07609_));
 sky130_as_sc_hs__and2_2 _38345_ (.A(_24774_),
    .B(net420),
    .Y(_07612_));
 sky130_as_sc_hs__and2_2 _38346_ (.A(net446),
    .B(net441),
    .Y(_07613_));
 sky130_as_sc_hs__or2_2 _38348_ (.A(_07612_),
    .B(_07613_),
    .Y(_07615_));
 sky130_as_sc_hs__and2_2 _38349_ (.A(_07614_),
    .B(_07615_),
    .Y(_07616_));
 sky130_as_sc_hs__or2_2 _38352_ (.A(_07616_),
    .B(_07617_),
    .Y(_07619_));
 sky130_as_sc_hs__and2_2 _38353_ (.A(_07618_),
    .B(_07619_),
    .Y(_07620_));
 sky130_as_sc_hs__and2_2 _38354_ (.A(net79),
    .B(net436),
    .Y(_07621_));
 sky130_as_sc_hs__or2_2 _38356_ (.A(_07620_),
    .B(_07621_),
    .Y(_07623_));
 sky130_as_sc_hs__and2_2 _38357_ (.A(_07622_),
    .B(_07623_),
    .Y(_07624_));
 sky130_as_sc_hs__and2_2 _38360_ (.A(net444),
    .B(net427),
    .Y(_07627_));
 sky130_as_sc_hs__and2_2 _38361_ (.A(net85),
    .B(net434),
    .Y(_07628_));
 sky130_as_sc_hs__or2_2 _38362_ (.A(_07627_),
    .B(_07628_),
    .Y(_07629_));
 sky130_as_sc_hs__and2_2 _38364_ (.A(_07629_),
    .B(_07630_),
    .Y(_07631_));
 sky130_as_sc_hs__and2_2 _38365_ (.A(net123),
    .B(_24729_),
    .Y(_07632_));
 sky130_as_sc_hs__or2_2 _38367_ (.A(_07631_),
    .B(_07632_),
    .Y(_07634_));
 sky130_as_sc_hs__and2_2 _38368_ (.A(_07633_),
    .B(_07634_),
    .Y(_07635_));
 sky130_as_sc_hs__or2_2 _38370_ (.A(_07626_),
    .B(_07635_),
    .Y(_07637_));
 sky130_as_sc_hs__and2_2 _38371_ (.A(_07636_),
    .B(_07637_),
    .Y(_07638_));
 sky130_as_sc_hs__or2_2 _38373_ (.A(_07625_),
    .B(_07638_),
    .Y(_07640_));
 sky130_as_sc_hs__and2_2 _38374_ (.A(_07639_),
    .B(_07640_),
    .Y(_07641_));
 sky130_as_sc_hs__or2_2 _38377_ (.A(_07641_),
    .B(_07642_),
    .Y(_07644_));
 sky130_as_sc_hs__and2_2 _38378_ (.A(_07643_),
    .B(_07644_),
    .Y(_07645_));
 sky130_as_sc_hs__or2_2 _38380_ (.A(_07624_),
    .B(_07645_),
    .Y(_07647_));
 sky130_as_sc_hs__and2_2 _38381_ (.A(_07646_),
    .B(_07647_),
    .Y(_07648_));
 sky130_as_sc_hs__or2_2 _38383_ (.A(_07611_),
    .B(_07648_),
    .Y(_07650_));
 sky130_as_sc_hs__and2_2 _38384_ (.A(_07649_),
    .B(_07650_),
    .Y(_07651_));
 sky130_as_sc_hs__or2_2 _38386_ (.A(_07610_),
    .B(_07651_),
    .Y(_07653_));
 sky130_as_sc_hs__and2_2 _38387_ (.A(_07652_),
    .B(_07653_),
    .Y(_07654_));
 sky130_as_sc_hs__and2_2 _38390_ (.A(net449),
    .B(net431),
    .Y(_07657_));
 sky130_as_sc_hs__and2_2 _38391_ (.A(_24545_),
    .B(net426),
    .Y(_07658_));
 sky130_as_sc_hs__or2_2 _38392_ (.A(_07657_),
    .B(_07658_),
    .Y(_07659_));
 sky130_as_sc_hs__and2_2 _38394_ (.A(_07659_),
    .B(_07660_),
    .Y(_07661_));
 sky130_as_sc_hs__and2_2 _38395_ (.A(net451),
    .B(net429),
    .Y(_07662_));
 sky130_as_sc_hs__or2_2 _38397_ (.A(_07661_),
    .B(_07662_),
    .Y(_07664_));
 sky130_as_sc_hs__and2_2 _38398_ (.A(_07663_),
    .B(_07664_),
    .Y(_07665_));
 sky130_as_sc_hs__and2_2 _38399_ (.A(net479),
    .B(_24527_),
    .Y(_07666_));
 sky130_as_sc_hs__and2_2 _38400_ (.A(net474),
    .B(net89),
    .Y(_07667_));
 sky130_as_sc_hs__or2_2 _38401_ (.A(_07666_),
    .B(_07667_),
    .Y(_07668_));
 sky130_as_sc_hs__and2_2 _38403_ (.A(_07668_),
    .B(_07669_),
    .Y(_07670_));
 sky130_as_sc_hs__and2_2 _38404_ (.A(net88),
    .B(net84),
    .Y(_07671_));
 sky130_as_sc_hs__or2_2 _38406_ (.A(_07670_),
    .B(_07671_),
    .Y(_07673_));
 sky130_as_sc_hs__and2_2 _38407_ (.A(_07672_),
    .B(_07673_),
    .Y(_07674_));
 sky130_as_sc_hs__or2_2 _38410_ (.A(_07674_),
    .B(_07675_),
    .Y(_07677_));
 sky130_as_sc_hs__and2_2 _38411_ (.A(_07676_),
    .B(_07677_),
    .Y(_07678_));
 sky130_as_sc_hs__or2_2 _38413_ (.A(_07665_),
    .B(_07678_),
    .Y(_07680_));
 sky130_as_sc_hs__and2_2 _38414_ (.A(_07679_),
    .B(_07680_),
    .Y(_07681_));
 sky130_as_sc_hs__or2_2 _38416_ (.A(_07656_),
    .B(_07681_),
    .Y(_07683_));
 sky130_as_sc_hs__and2_2 _38417_ (.A(_07682_),
    .B(_07683_),
    .Y(_07684_));
 sky130_as_sc_hs__or2_2 _38419_ (.A(_07655_),
    .B(_07684_),
    .Y(_07686_));
 sky130_as_sc_hs__and2_2 _38420_ (.A(_07685_),
    .B(_07686_),
    .Y(_07687_));
 sky130_as_sc_hs__and2_2 _38423_ (.A(net476),
    .B(net465),
    .Y(_07690_));
 sky130_as_sc_hs__and2_2 _38424_ (.A(net463),
    .B(net438),
    .Y(_07691_));
 sky130_as_sc_hs__or2_2 _38425_ (.A(_07690_),
    .B(_07691_),
    .Y(_07692_));
 sky130_as_sc_hs__and2_2 _38427_ (.A(_07692_),
    .B(_07693_),
    .Y(_07694_));
 sky130_as_sc_hs__and2_2 _38428_ (.A(net472),
    .B(net460),
    .Y(_07695_));
 sky130_as_sc_hs__or2_2 _38430_ (.A(_07694_),
    .B(_07695_),
    .Y(_07697_));
 sky130_as_sc_hs__and2_2 _38431_ (.A(_07696_),
    .B(_07697_),
    .Y(_07698_));
 sky130_as_sc_hs__or2_2 _38433_ (.A(_07689_),
    .B(_07698_),
    .Y(_07700_));
 sky130_as_sc_hs__and2_2 _38434_ (.A(_07699_),
    .B(_07700_),
    .Y(_07701_));
 sky130_as_sc_hs__or2_2 _38436_ (.A(_07688_),
    .B(_07701_),
    .Y(_07703_));
 sky130_as_sc_hs__and2_2 _38437_ (.A(_07702_),
    .B(_07703_),
    .Y(_07704_));
 sky130_as_sc_hs__and2_2 _38438_ (.A(net467),
    .B(net442),
    .Y(_07705_));
 sky130_as_sc_hs__and2_2 _38439_ (.A(_23674_),
    .B(net469),
    .Y(_07706_));
 sky130_as_sc_hs__or2_2 _38440_ (.A(_07705_),
    .B(_07706_),
    .Y(_07707_));
 sky130_as_sc_hs__and2_2 _38442_ (.A(_07707_),
    .B(_07708_),
    .Y(_07709_));
 sky130_as_sc_hs__and2_2 _38443_ (.A(net480),
    .B(net471),
    .Y(_07710_));
 sky130_as_sc_hs__or2_2 _38445_ (.A(_07709_),
    .B(_07710_),
    .Y(_07712_));
 sky130_as_sc_hs__and2_2 _38446_ (.A(_07711_),
    .B(_07712_),
    .Y(_07713_));
 sky130_as_sc_hs__and2_2 _38447_ (.A(net456),
    .B(net452),
    .Y(_07714_));
 sky130_as_sc_hs__or2_2 _38451_ (.A(_07715_),
    .B(_07716_),
    .Y(_07718_));
 sky130_as_sc_hs__and2_2 _38452_ (.A(_07717_),
    .B(_07718_),
    .Y(_07719_));
 sky130_as_sc_hs__or2_2 _38454_ (.A(_07714_),
    .B(_07719_),
    .Y(_07721_));
 sky130_as_sc_hs__and2_2 _38455_ (.A(_07720_),
    .B(_07721_),
    .Y(_07722_));
 sky130_as_sc_hs__or2_2 _38458_ (.A(_07722_),
    .B(_07723_),
    .Y(_07725_));
 sky130_as_sc_hs__and2_2 _38459_ (.A(_07724_),
    .B(_07725_),
    .Y(_07726_));
 sky130_as_sc_hs__or2_2 _38461_ (.A(_07713_),
    .B(_07726_),
    .Y(_07728_));
 sky130_as_sc_hs__and2_2 _38462_ (.A(_07727_),
    .B(_07728_),
    .Y(_07729_));
 sky130_as_sc_hs__or2_2 _38465_ (.A(_07729_),
    .B(_07730_),
    .Y(_07732_));
 sky130_as_sc_hs__and2_2 _38466_ (.A(_07731_),
    .B(_07732_),
    .Y(_07733_));
 sky130_as_sc_hs__or2_2 _38468_ (.A(_07704_),
    .B(_07733_),
    .Y(_07735_));
 sky130_as_sc_hs__and2_2 _38469_ (.A(_07734_),
    .B(_07735_),
    .Y(_07736_));
 sky130_as_sc_hs__or2_2 _38472_ (.A(_07736_),
    .B(_07737_),
    .Y(_07739_));
 sky130_as_sc_hs__and2_2 _38473_ (.A(_07738_),
    .B(_07739_),
    .Y(_07740_));
 sky130_as_sc_hs__or2_2 _38475_ (.A(_07687_),
    .B(_07740_),
    .Y(_07742_));
 sky130_as_sc_hs__and2_2 _38476_ (.A(_07741_),
    .B(_07742_),
    .Y(_07743_));
 sky130_as_sc_hs__or2_2 _38479_ (.A(_07743_),
    .B(_07744_),
    .Y(_07746_));
 sky130_as_sc_hs__and2_2 _38480_ (.A(_07745_),
    .B(_07746_),
    .Y(_07747_));
 sky130_as_sc_hs__or2_2 _38482_ (.A(_07654_),
    .B(_07747_),
    .Y(_07749_));
 sky130_as_sc_hs__and2_2 _38483_ (.A(_07748_),
    .B(_07749_),
    .Y(_07750_));
 sky130_as_sc_hs__or2_2 _38486_ (.A(_07750_),
    .B(_07751_),
    .Y(_07753_));
 sky130_as_sc_hs__and2_2 _38487_ (.A(_07752_),
    .B(_07753_),
    .Y(_07754_));
 sky130_as_sc_hs__or2_2 _38489_ (.A(_07609_),
    .B(_07754_),
    .Y(_07756_));
 sky130_as_sc_hs__and2_2 _38490_ (.A(_07755_),
    .B(_07756_),
    .Y(_07757_));
 sky130_as_sc_hs__or2_2 _38493_ (.A(_07757_),
    .B(_07758_),
    .Y(_07760_));
 sky130_as_sc_hs__and2_2 _38494_ (.A(_07759_),
    .B(_07760_),
    .Y(_07761_));
 sky130_as_sc_hs__or2_2 _38496_ (.A(_07566_),
    .B(_07761_),
    .Y(_07763_));
 sky130_as_sc_hs__and2_2 _38497_ (.A(_07762_),
    .B(_07763_),
    .Y(_07764_));
 sky130_as_sc_hs__or2_2 _38500_ (.A(_07764_),
    .B(_07765_),
    .Y(_07767_));
 sky130_as_sc_hs__and2_2 _38501_ (.A(_07766_),
    .B(_07767_),
    .Y(_07768_));
 sky130_as_sc_hs__or2_2 _38503_ (.A(_07565_),
    .B(_07768_),
    .Y(_07770_));
 sky130_as_sc_hs__and2_2 _38504_ (.A(_07769_),
    .B(_07770_),
    .Y(_07771_));
 sky130_as_sc_hs__nand3_2 _38506_ (.A(_07769_),
    .B(_07770_),
    .C(_07772_),
    .Y(_07773_));
 sky130_as_sc_hs__or2_2 _38507_ (.A(_07771_),
    .B(_07772_),
    .Y(_07774_));
 sky130_as_sc_hs__and2_2 _38508_ (.A(_07773_),
    .B(_07774_),
    .Y(_07775_));
 sky130_as_sc_hs__or2_2 _38510_ (.A(_07775_),
    .B(_07776_),
    .Y(_07777_));
 sky130_as_sc_hs__or2_2 _38514_ (.A(_07779_),
    .B(_07780_),
    .Y(_07781_));
 sky130_as_sc_hs__nand3_2 _38516_ (.A(net142),
    .B(_07781_),
    .C(_07782_),
    .Y(_07783_));
 sky130_as_sc_hs__and2_2 _38517_ (.A(_04522_),
    .B(_05405_),
    .Y(_07784_));
 sky130_as_sc_hs__or2_2 _38518_ (.A(_04523_),
    .B(_07784_),
    .Y(_07785_));
 sky130_as_sc_hs__or2_2 _38521_ (.A(_07785_),
    .B(_07786_),
    .Y(_07788_));
 sky130_as_sc_hs__nand3_2 _38522_ (.A(net139),
    .B(_07787_),
    .C(_07788_),
    .Y(_07789_));
 sky130_as_sc_hs__or2_2 _38524_ (.A(_05793_),
    .B(_07500_),
    .Y(_07791_));
 sky130_as_sc_hs__or2_2 _38527_ (.A(_05779_),
    .B(_07792_),
    .Y(_07794_));
 sky130_as_sc_hs__nand3_2 _38532_ (.A(net119),
    .B(_07796_),
    .C(_07798_),
    .Y(_07799_));
 sky130_as_sc_hs__or2_2 _38533_ (.A(_05941_),
    .B(_06462_),
    .Y(_07800_));
 sky130_as_sc_hs__nand3_2 _38535_ (.A(_05935_),
    .B(_07800_),
    .C(_07801_),
    .Y(_07802_));
 sky130_as_sc_hs__or2_2 _38539_ (.A(_05935_),
    .B(_07805_),
    .Y(_07806_));
 sky130_as_sc_hs__and2_2 _38542_ (.A(_07807_),
    .B(_07808_),
    .Y(_07809_));
 sky130_as_sc_hs__or2_2 _38544_ (.A(_05935_),
    .B(_06906_),
    .Y(_07811_));
 sky130_as_sc_hs__and2_2 _38545_ (.A(_07810_),
    .B(_07811_),
    .Y(_07812_));
 sky130_as_sc_hs__nand3_2 _38546_ (.A(_05929_),
    .B(_07802_),
    .C(_07806_),
    .Y(_07813_));
 sky130_as_sc_hs__and2_2 _38554_ (.A(net140),
    .B(_07820_),
    .Y(_07821_));
 sky130_as_sc_hs__or2_2 _38555_ (.A(\tholin_riscv.div_res[4] ),
    .B(_07533_),
    .Y(_07822_));
 sky130_as_sc_hs__and2_2 _38556_ (.A(net415),
    .B(_07822_),
    .Y(_07823_));
 sky130_as_sc_hs__or2_2 _38557_ (.A(\tholin_riscv.div_res[5] ),
    .B(_07823_),
    .Y(_07824_));
 sky130_as_sc_hs__nand3_2 _38559_ (.A(net111),
    .B(_07824_),
    .C(_07825_),
    .Y(_07826_));
 sky130_as_sc_hs__nor2_2 _38563_ (.A(_05777_),
    .B(_06161_),
    .Y(_07830_));
 sky130_as_sc_hs__or2_2 _38564_ (.A(\tholin_riscv.div_shifter[36] ),
    .B(_07539_),
    .Y(_07831_));
 sky130_as_sc_hs__and2_2 _38565_ (.A(_21655_),
    .B(_07831_),
    .Y(_07832_));
 sky130_as_sc_hs__or2_2 _38567_ (.A(\tholin_riscv.div_shifter[37] ),
    .B(_07832_),
    .Y(_07834_));
 sky130_as_sc_hs__nand3_2 _38568_ (.A(net109),
    .B(_07833_),
    .C(_07834_),
    .Y(_07835_));
 sky130_as_sc_hs__and2_2 _38571_ (.A(_07836_),
    .B(_07837_),
    .Y(_07838_));
 sky130_as_sc_hs__nand3_2 _38572_ (.A(net413),
    .B(_07835_),
    .C(_07838_),
    .Y(_07839_));
 sky130_as_sc_hs__nor2_2 _38573_ (.A(_07830_),
    .B(_07839_),
    .Y(_07840_));
 sky130_as_sc_hs__nand3_2 _38574_ (.A(_07826_),
    .B(_07829_),
    .C(_07840_),
    .Y(_07841_));
 sky130_as_sc_hs__nor2_2 _38575_ (.A(_07821_),
    .B(_07841_),
    .Y(_07842_));
 sky130_as_sc_hs__and2_2 _38576_ (.A(_07816_),
    .B(_07842_),
    .Y(_07843_));
 sky130_as_sc_hs__and2_2 _38577_ (.A(_07799_),
    .B(_07843_),
    .Y(_07844_));
 sky130_as_sc_hs__nand3_2 _38578_ (.A(_07783_),
    .B(_07789_),
    .C(_07844_),
    .Y(_07845_));
 sky130_as_sc_hs__and2_2 _38579_ (.A(\tholin_riscv.PC[5] ),
    .B(_07554_),
    .Y(_07846_));
 sky130_as_sc_hs__nor2_2 _38580_ (.A(\tholin_riscv.PC[5] ),
    .B(_07554_),
    .Y(_07847_));
 sky130_as_sc_hs__nor2_2 _38581_ (.A(_07846_),
    .B(_07847_),
    .Y(_07848_));
 sky130_as_sc_hs__nand3_2 _38584_ (.A(_21569_),
    .B(_07849_),
    .C(_07850_),
    .Y(_07851_));
 sky130_as_sc_hs__nand3_2 _38585_ (.A(_21546_),
    .B(_07845_),
    .C(_07851_),
    .Y(_07852_));
 sky130_as_sc_hs__and2_2 _38595_ (.A(_24545_),
    .B(net422),
    .Y(_07861_));
 sky130_as_sc_hs__and2_2 _38596_ (.A(net122),
    .B(_23624_),
    .Y(_07862_));
 sky130_as_sc_hs__or2_2 _38597_ (.A(_07861_),
    .B(_07862_),
    .Y(_07863_));
 sky130_as_sc_hs__inv_2 _38599_ (.Y(_07865_),
    .A(_07864_));
 sky130_as_sc_hs__and2_2 _38600_ (.A(_07863_),
    .B(_07864_),
    .Y(_07866_));
 sky130_as_sc_hs__or2_2 _38603_ (.A(_07866_),
    .B(_07867_),
    .Y(_07869_));
 sky130_as_sc_hs__or2_2 _38605_ (.A(_07579_),
    .B(_07870_),
    .Y(_07871_));
 sky130_as_sc_hs__and2_2 _38607_ (.A(_07871_),
    .B(_07872_),
    .Y(_07873_));
 sky130_as_sc_hs__and2_2 _38608_ (.A(_23702_),
    .B(net420),
    .Y(_07874_));
 sky130_as_sc_hs__or2_2 _38610_ (.A(_07873_),
    .B(_07874_),
    .Y(_07876_));
 sky130_as_sc_hs__and2_2 _38611_ (.A(_07875_),
    .B(_07876_),
    .Y(_07877_));
 sky130_as_sc_hs__and2_2 _38613_ (.A(_24501_),
    .B(net129),
    .Y(_07879_));
 sky130_as_sc_hs__or2_2 _38615_ (.A(_07878_),
    .B(_07879_),
    .Y(_07881_));
 sky130_as_sc_hs__and2_2 _38616_ (.A(_07880_),
    .B(_07881_),
    .Y(_07882_));
 sky130_as_sc_hs__or2_2 _38619_ (.A(_07882_),
    .B(_07883_),
    .Y(_07885_));
 sky130_as_sc_hs__and2_2 _38620_ (.A(_07884_),
    .B(_07885_),
    .Y(_07886_));
 sky130_as_sc_hs__or2_2 _38622_ (.A(_07877_),
    .B(_07886_),
    .Y(_07888_));
 sky130_as_sc_hs__and2_2 _38623_ (.A(_07887_),
    .B(_07888_),
    .Y(_07889_));
 sky130_as_sc_hs__or2_2 _38625_ (.A(_07860_),
    .B(_07889_),
    .Y(_07891_));
 sky130_as_sc_hs__and2_2 _38626_ (.A(_07890_),
    .B(_07891_),
    .Y(_07892_));
 sky130_as_sc_hs__or2_2 _38628_ (.A(_07859_),
    .B(_07892_),
    .Y(_07894_));
 sky130_as_sc_hs__and2_2 _38629_ (.A(_07893_),
    .B(_07894_),
    .Y(_07895_));
 sky130_as_sc_hs__and2_2 _38632_ (.A(_24774_),
    .B(net75),
    .Y(_07898_));
 sky130_as_sc_hs__and2_2 _38633_ (.A(net78),
    .B(net441),
    .Y(_07899_));
 sky130_as_sc_hs__or2_2 _38634_ (.A(_07898_),
    .B(_07899_),
    .Y(_07900_));
 sky130_as_sc_hs__or2_2 _38637_ (.A(_07614_),
    .B(_07902_),
    .Y(_07903_));
 sky130_as_sc_hs__and2_2 _38639_ (.A(_07903_),
    .B(_07904_),
    .Y(_07905_));
 sky130_as_sc_hs__and2_2 _38640_ (.A(net442),
    .B(net436),
    .Y(_07906_));
 sky130_as_sc_hs__or2_2 _38642_ (.A(_07905_),
    .B(_07906_),
    .Y(_07908_));
 sky130_as_sc_hs__and2_2 _38643_ (.A(_07907_),
    .B(_07908_),
    .Y(_07909_));
 sky130_as_sc_hs__or2_2 _38649_ (.A(_07912_),
    .B(_07913_),
    .Y(_07915_));
 sky130_as_sc_hs__and2_2 _38650_ (.A(_07914_),
    .B(_07915_),
    .Y(_07916_));
 sky130_as_sc_hs__and2_2 _38651_ (.A(_24729_),
    .B(net424),
    .Y(_07917_));
 sky130_as_sc_hs__or2_2 _38653_ (.A(_07916_),
    .B(_07917_),
    .Y(_07919_));
 sky130_as_sc_hs__and2_2 _38654_ (.A(_07918_),
    .B(_07919_),
    .Y(_07920_));
 sky130_as_sc_hs__or2_2 _38656_ (.A(_07911_),
    .B(_07920_),
    .Y(_07922_));
 sky130_as_sc_hs__and2_2 _38657_ (.A(_07921_),
    .B(_07922_),
    .Y(_07923_));
 sky130_as_sc_hs__or2_2 _38659_ (.A(_07910_),
    .B(_07923_),
    .Y(_07925_));
 sky130_as_sc_hs__and2_2 _38660_ (.A(_07924_),
    .B(_07925_),
    .Y(_07926_));
 sky130_as_sc_hs__or2_2 _38663_ (.A(_07926_),
    .B(_07927_),
    .Y(_07929_));
 sky130_as_sc_hs__and2_2 _38664_ (.A(_07928_),
    .B(_07929_),
    .Y(_07930_));
 sky130_as_sc_hs__or2_2 _38666_ (.A(_07909_),
    .B(_07930_),
    .Y(_07932_));
 sky130_as_sc_hs__and2_2 _38667_ (.A(_07931_),
    .B(_07932_),
    .Y(_07933_));
 sky130_as_sc_hs__or2_2 _38669_ (.A(_07897_),
    .B(_07933_),
    .Y(_07935_));
 sky130_as_sc_hs__and2_2 _38670_ (.A(_07934_),
    .B(_07935_),
    .Y(_07936_));
 sky130_as_sc_hs__or2_2 _38672_ (.A(_07896_),
    .B(_07936_),
    .Y(_07938_));
 sky130_as_sc_hs__and2_2 _38673_ (.A(_07937_),
    .B(_07938_),
    .Y(_07939_));
 sky130_as_sc_hs__and2_2 _38676_ (.A(net449),
    .B(net429),
    .Y(_07942_));
 sky130_as_sc_hs__and2_2 _38677_ (.A(net454),
    .B(net426),
    .Y(_07943_));
 sky130_as_sc_hs__or2_2 _38678_ (.A(_07942_),
    .B(_07943_),
    .Y(_07944_));
 sky130_as_sc_hs__and2_2 _38680_ (.A(_07944_),
    .B(_07945_),
    .Y(_07946_));
 sky130_as_sc_hs__and2_2 _38681_ (.A(net451),
    .B(net427),
    .Y(_07947_));
 sky130_as_sc_hs__or2_2 _38683_ (.A(_07946_),
    .B(_07947_),
    .Y(_07949_));
 sky130_as_sc_hs__and2_2 _38684_ (.A(_07948_),
    .B(_07949_),
    .Y(_07950_));
 sky130_as_sc_hs__and2_2 _38685_ (.A(net474),
    .B(_24527_),
    .Y(_07951_));
 sky130_as_sc_hs__and2_2 _38686_ (.A(net89),
    .B(net83),
    .Y(_07952_));
 sky130_as_sc_hs__or2_2 _38687_ (.A(_07951_),
    .B(_07952_),
    .Y(_07953_));
 sky130_as_sc_hs__and2_2 _38689_ (.A(_07953_),
    .B(_07954_),
    .Y(_07955_));
 sky130_as_sc_hs__and2_2 _38690_ (.A(net88),
    .B(net431),
    .Y(_07956_));
 sky130_as_sc_hs__or2_2 _38692_ (.A(_07955_),
    .B(_07956_),
    .Y(_07958_));
 sky130_as_sc_hs__and2_2 _38693_ (.A(_07957_),
    .B(_07958_),
    .Y(_07959_));
 sky130_as_sc_hs__or2_2 _38696_ (.A(_07959_),
    .B(_07960_),
    .Y(_07962_));
 sky130_as_sc_hs__and2_2 _38697_ (.A(_07961_),
    .B(_07962_),
    .Y(_07963_));
 sky130_as_sc_hs__or2_2 _38699_ (.A(_07950_),
    .B(_07963_),
    .Y(_07965_));
 sky130_as_sc_hs__and2_2 _38700_ (.A(_07964_),
    .B(_07965_),
    .Y(_07966_));
 sky130_as_sc_hs__or2_2 _38702_ (.A(_07941_),
    .B(_07966_),
    .Y(_07968_));
 sky130_as_sc_hs__and2_2 _38703_ (.A(_07967_),
    .B(_07968_),
    .Y(_07969_));
 sky130_as_sc_hs__or2_2 _38705_ (.A(_07940_),
    .B(_07969_),
    .Y(_07971_));
 sky130_as_sc_hs__and2_2 _38706_ (.A(_07970_),
    .B(_07971_),
    .Y(_07972_));
 sky130_as_sc_hs__and2_2 _38709_ (.A(net465),
    .B(net438),
    .Y(_07975_));
 sky130_as_sc_hs__and2_2 _38710_ (.A(net472),
    .B(net463),
    .Y(_07976_));
 sky130_as_sc_hs__or2_2 _38711_ (.A(_07975_),
    .B(_07976_),
    .Y(_07977_));
 sky130_as_sc_hs__and2_2 _38713_ (.A(_07977_),
    .B(_07978_),
    .Y(_07979_));
 sky130_as_sc_hs__and2_2 _38714_ (.A(net478),
    .B(net460),
    .Y(_07980_));
 sky130_as_sc_hs__or2_2 _38716_ (.A(_07979_),
    .B(_07980_),
    .Y(_07982_));
 sky130_as_sc_hs__and2_2 _38717_ (.A(_07981_),
    .B(_07982_),
    .Y(_07983_));
 sky130_as_sc_hs__or2_2 _38719_ (.A(_07974_),
    .B(_07983_),
    .Y(_07985_));
 sky130_as_sc_hs__and2_2 _38720_ (.A(_07984_),
    .B(_07985_),
    .Y(_07986_));
 sky130_as_sc_hs__or2_2 _38722_ (.A(_07973_),
    .B(_07986_),
    .Y(_07988_));
 sky130_as_sc_hs__and2_2 _38723_ (.A(_07987_),
    .B(_07988_),
    .Y(_07989_));
 sky130_as_sc_hs__and2_2 _38724_ (.A(_23674_),
    .B(net466),
    .Y(_07990_));
 sky130_as_sc_hs__and2_2 _38725_ (.A(net480),
    .B(net468),
    .Y(_07991_));
 sky130_as_sc_hs__or2_2 _38726_ (.A(_07990_),
    .B(_07991_),
    .Y(_07992_));
 sky130_as_sc_hs__and2_2 _38728_ (.A(_07992_),
    .B(_07993_),
    .Y(_07994_));
 sky130_as_sc_hs__and2_2 _38729_ (.A(net476),
    .B(net471),
    .Y(_07995_));
 sky130_as_sc_hs__or2_2 _38731_ (.A(_07994_),
    .B(_07995_),
    .Y(_07997_));
 sky130_as_sc_hs__and2_2 _38732_ (.A(_07996_),
    .B(_07997_),
    .Y(_07998_));
 sky130_as_sc_hs__and2_2 _38733_ (.A(net457),
    .B(net446),
    .Y(_07999_));
 sky130_as_sc_hs__or2_2 _38737_ (.A(_08000_),
    .B(_08001_),
    .Y(_08003_));
 sky130_as_sc_hs__and2_2 _38738_ (.A(_08002_),
    .B(_08003_),
    .Y(_08004_));
 sky130_as_sc_hs__or2_2 _38740_ (.A(_07999_),
    .B(_08004_),
    .Y(_08006_));
 sky130_as_sc_hs__and2_2 _38741_ (.A(_08005_),
    .B(_08006_),
    .Y(_08007_));
 sky130_as_sc_hs__or2_2 _38744_ (.A(_08007_),
    .B(_08008_),
    .Y(_08010_));
 sky130_as_sc_hs__and2_2 _38745_ (.A(_08009_),
    .B(_08010_),
    .Y(_08011_));
 sky130_as_sc_hs__or2_2 _38747_ (.A(_07998_),
    .B(_08011_),
    .Y(_08013_));
 sky130_as_sc_hs__and2_2 _38748_ (.A(_08012_),
    .B(_08013_),
    .Y(_08014_));
 sky130_as_sc_hs__or2_2 _38751_ (.A(_08014_),
    .B(_08015_),
    .Y(_08017_));
 sky130_as_sc_hs__and2_2 _38752_ (.A(_08016_),
    .B(_08017_),
    .Y(_08018_));
 sky130_as_sc_hs__or2_2 _38754_ (.A(_07989_),
    .B(_08018_),
    .Y(_08020_));
 sky130_as_sc_hs__and2_2 _38755_ (.A(_08019_),
    .B(_08020_),
    .Y(_08021_));
 sky130_as_sc_hs__or2_2 _38758_ (.A(_08021_),
    .B(_08022_),
    .Y(_08024_));
 sky130_as_sc_hs__and2_2 _38759_ (.A(_08023_),
    .B(_08024_),
    .Y(_08025_));
 sky130_as_sc_hs__or2_2 _38761_ (.A(_07972_),
    .B(_08025_),
    .Y(_08027_));
 sky130_as_sc_hs__and2_2 _38762_ (.A(_08026_),
    .B(_08027_),
    .Y(_08028_));
 sky130_as_sc_hs__or2_2 _38765_ (.A(_08028_),
    .B(_08029_),
    .Y(_08031_));
 sky130_as_sc_hs__and2_2 _38766_ (.A(_08030_),
    .B(_08031_),
    .Y(_08032_));
 sky130_as_sc_hs__or2_2 _38768_ (.A(_07939_),
    .B(_08032_),
    .Y(_08034_));
 sky130_as_sc_hs__and2_2 _38769_ (.A(_08033_),
    .B(_08034_),
    .Y(_08035_));
 sky130_as_sc_hs__or2_2 _38772_ (.A(_08035_),
    .B(_08036_),
    .Y(_08038_));
 sky130_as_sc_hs__and2_2 _38773_ (.A(_08037_),
    .B(_08038_),
    .Y(_08039_));
 sky130_as_sc_hs__or2_2 _38775_ (.A(_07895_),
    .B(_08039_),
    .Y(_08041_));
 sky130_as_sc_hs__and2_2 _38776_ (.A(_08040_),
    .B(_08041_),
    .Y(_08042_));
 sky130_as_sc_hs__or2_2 _38779_ (.A(_08042_),
    .B(_08043_),
    .Y(_08045_));
 sky130_as_sc_hs__and2_2 _38780_ (.A(_08044_),
    .B(_08045_),
    .Y(_08046_));
 sky130_as_sc_hs__or2_2 _38782_ (.A(_07858_),
    .B(_08046_),
    .Y(_08048_));
 sky130_as_sc_hs__and2_2 _38783_ (.A(_08047_),
    .B(_08048_),
    .Y(_08049_));
 sky130_as_sc_hs__or2_2 _38786_ (.A(_08049_),
    .B(_08050_),
    .Y(_08052_));
 sky130_as_sc_hs__and2_2 _38787_ (.A(_08051_),
    .B(_08052_),
    .Y(_08053_));
 sky130_as_sc_hs__or2_2 _38789_ (.A(_07857_),
    .B(_08053_),
    .Y(_08055_));
 sky130_as_sc_hs__and2_2 _38790_ (.A(_08054_),
    .B(_08055_),
    .Y(_08056_));
 sky130_as_sc_hs__or2_2 _38793_ (.A(_08056_),
    .B(_08057_),
    .Y(_08059_));
 sky130_as_sc_hs__and2_2 _38794_ (.A(_08058_),
    .B(_08059_),
    .Y(_08060_));
 sky130_as_sc_hs__inv_2 _38797_ (.Y(_08063_),
    .A(_08062_));
 sky130_as_sc_hs__and2_2 _38798_ (.A(_07474_),
    .B(_07775_),
    .Y(_08064_));
 sky130_as_sc_hs__or2_2 _38802_ (.A(_08060_),
    .B(_08066_),
    .Y(_08068_));
 sky130_as_sc_hs__or2_2 _38805_ (.A(_07487_),
    .B(_08070_),
    .Y(_08071_));
 sky130_as_sc_hs__or2_2 _38807_ (.A(_08069_),
    .B(_08072_),
    .Y(_08073_));
 sky130_as_sc_hs__nand3_2 _38809_ (.A(net142),
    .B(_08073_),
    .C(_08074_),
    .Y(_08075_));
 sky130_as_sc_hs__or2_2 _38810_ (.A(_05406_),
    .B(_05505_),
    .Y(_08076_));
 sky130_as_sc_hs__or2_2 _38811_ (.A(_05396_),
    .B(_08076_),
    .Y(_08077_));
 sky130_as_sc_hs__nand3_2 _38813_ (.A(net139),
    .B(_08077_),
    .C(_08078_),
    .Y(_08079_));
 sky130_as_sc_hs__or2_2 _38816_ (.A(_05768_),
    .B(_08081_),
    .Y(_08082_));
 sky130_as_sc_hs__and2_2 _38818_ (.A(_08082_),
    .B(_08083_),
    .Y(_08084_));
 sky130_as_sc_hs__or2_2 _38820_ (.A(_05768_),
    .B(_05858_),
    .Y(_08086_));
 sky130_as_sc_hs__nand3_2 _38823_ (.A(net118),
    .B(_08085_),
    .C(_08088_),
    .Y(_08089_));
 sky130_as_sc_hs__or2_2 _38824_ (.A(_05940_),
    .B(_06842_),
    .Y(_08090_));
 sky130_as_sc_hs__or2_2 _38825_ (.A(_05941_),
    .B(_06834_),
    .Y(_08091_));
 sky130_as_sc_hs__nand3_2 _38826_ (.A(_05935_),
    .B(_08090_),
    .C(_08091_),
    .Y(_08092_));
 sky130_as_sc_hs__and2_2 _38829_ (.A(_08093_),
    .B(_08094_),
    .Y(_08095_));
 sky130_as_sc_hs__or2_2 _38830_ (.A(_05935_),
    .B(_08095_),
    .Y(_08096_));
 sky130_as_sc_hs__or2_2 _38835_ (.A(_05935_),
    .B(_06429_),
    .Y(_08101_));
 sky130_as_sc_hs__and2_2 _38836_ (.A(_08100_),
    .B(_08101_),
    .Y(_08102_));
 sky130_as_sc_hs__nand3_2 _38837_ (.A(_05929_),
    .B(_08092_),
    .C(_08096_),
    .Y(_08103_));
 sky130_as_sc_hs__and2_2 _38845_ (.A(net140),
    .B(_08110_),
    .Y(_08111_));
 sky130_as_sc_hs__or2_2 _38846_ (.A(\tholin_riscv.div_res[5] ),
    .B(_07822_),
    .Y(_08112_));
 sky130_as_sc_hs__and2_2 _38847_ (.A(net415),
    .B(_08112_),
    .Y(_08113_));
 sky130_as_sc_hs__or2_2 _38848_ (.A(\tholin_riscv.div_res[6] ),
    .B(_08113_),
    .Y(_08114_));
 sky130_as_sc_hs__nand3_2 _38850_ (.A(net111),
    .B(_08114_),
    .C(_08115_),
    .Y(_08116_));
 sky130_as_sc_hs__nor2_2 _38854_ (.A(_05766_),
    .B(_06161_),
    .Y(_08120_));
 sky130_as_sc_hs__or2_2 _38855_ (.A(\tholin_riscv.div_shifter[37] ),
    .B(_07831_),
    .Y(_08121_));
 sky130_as_sc_hs__and2_2 _38856_ (.A(_21655_),
    .B(_08121_),
    .Y(_08122_));
 sky130_as_sc_hs__or2_2 _38858_ (.A(\tholin_riscv.div_shifter[38] ),
    .B(_08122_),
    .Y(_08124_));
 sky130_as_sc_hs__nand3_2 _38859_ (.A(net109),
    .B(_08123_),
    .C(_08124_),
    .Y(_08125_));
 sky130_as_sc_hs__and2_2 _38862_ (.A(_08126_),
    .B(_08127_),
    .Y(_08128_));
 sky130_as_sc_hs__nand3_2 _38863_ (.A(net412),
    .B(_08125_),
    .C(_08128_),
    .Y(_08129_));
 sky130_as_sc_hs__nor2_2 _38864_ (.A(_08120_),
    .B(_08129_),
    .Y(_08130_));
 sky130_as_sc_hs__nand3_2 _38865_ (.A(_08116_),
    .B(_08119_),
    .C(_08130_),
    .Y(_08131_));
 sky130_as_sc_hs__nor2_2 _38866_ (.A(_08111_),
    .B(_08131_),
    .Y(_08132_));
 sky130_as_sc_hs__and2_2 _38867_ (.A(_08106_),
    .B(_08132_),
    .Y(_08133_));
 sky130_as_sc_hs__and2_2 _38868_ (.A(_08089_),
    .B(_08133_),
    .Y(_08134_));
 sky130_as_sc_hs__nand3_2 _38869_ (.A(_08075_),
    .B(_08079_),
    .C(_08134_),
    .Y(_08135_));
 sky130_as_sc_hs__and2_2 _38870_ (.A(\tholin_riscv.PC[6] ),
    .B(_07846_),
    .Y(_08136_));
 sky130_as_sc_hs__nor2_2 _38871_ (.A(\tholin_riscv.PC[6] ),
    .B(_07846_),
    .Y(_08137_));
 sky130_as_sc_hs__nor2_2 _38872_ (.A(_08136_),
    .B(_08137_),
    .Y(_08138_));
 sky130_as_sc_hs__inv_2 _38873_ (.Y(_08139_),
    .A(_08138_));
 sky130_as_sc_hs__nand3_2 _38876_ (.A(_21569_),
    .B(_08140_),
    .C(_08141_),
    .Y(_08142_));
 sky130_as_sc_hs__nand3_2 _38877_ (.A(_21546_),
    .B(_08135_),
    .C(_08142_),
    .Y(_08143_));
 sky130_as_sc_hs__and2_2 _38888_ (.A(_23702_),
    .B(net75),
    .Y(_08153_));
 sky130_as_sc_hs__and2_2 _38889_ (.A(net454),
    .B(net422),
    .Y(_08154_));
 sky130_as_sc_hs__and2_2 _38890_ (.A(_23624_),
    .B(net424),
    .Y(_08155_));
 sky130_as_sc_hs__and2_2 _38891_ (.A(_08154_),
    .B(_08155_),
    .Y(_08156_));
 sky130_as_sc_hs__nor2_2 _38892_ (.A(_08154_),
    .B(_08155_),
    .Y(_08157_));
 sky130_as_sc_hs__nor2_2 _38893_ (.A(_08156_),
    .B(_08157_),
    .Y(_08158_));
 sky130_as_sc_hs__or2_2 _38895_ (.A(_08158_),
    .B(_08159_),
    .Y(_08160_));
 sky130_as_sc_hs__and2_2 _38897_ (.A(_08160_),
    .B(_08161_),
    .Y(_08162_));
 sky130_as_sc_hs__or2_2 _38899_ (.A(_08153_),
    .B(_08162_),
    .Y(_08164_));
 sky130_as_sc_hs__and2_2 _38900_ (.A(_08163_),
    .B(_08164_),
    .Y(_08165_));
 sky130_as_sc_hs__and2_2 _38902_ (.A(_24545_),
    .B(net129),
    .Y(_08167_));
 sky130_as_sc_hs__or2_2 _38904_ (.A(_08166_),
    .B(_08167_),
    .Y(_08169_));
 sky130_as_sc_hs__or2_2 _38906_ (.A(_07880_),
    .B(_08170_),
    .Y(_08171_));
 sky130_as_sc_hs__and2_2 _38908_ (.A(_08171_),
    .B(_08172_),
    .Y(_08173_));
 sky130_as_sc_hs__or2_2 _38910_ (.A(_08165_),
    .B(_08173_),
    .Y(_08175_));
 sky130_as_sc_hs__and2_2 _38911_ (.A(_08174_),
    .B(_08175_),
    .Y(_08176_));
 sky130_as_sc_hs__or2_2 _38913_ (.A(_08152_),
    .B(_08176_),
    .Y(_08178_));
 sky130_as_sc_hs__and2_2 _38914_ (.A(_08177_),
    .B(_08178_),
    .Y(_08179_));
 sky130_as_sc_hs__or2_2 _38916_ (.A(_08151_),
    .B(_08179_),
    .Y(_08181_));
 sky130_as_sc_hs__and2_2 _38917_ (.A(_08180_),
    .B(_08181_),
    .Y(_08182_));
 sky130_as_sc_hs__nand3_2 _38922_ (.A(net442),
    .B(_07898_),
    .C(_07899_),
    .Y(_08187_));
 sky130_as_sc_hs__and2_2 _38923_ (.A(_08186_),
    .B(_08187_),
    .Y(_08188_));
 sky130_as_sc_hs__and2_2 _38924_ (.A(_23674_),
    .B(net437),
    .Y(_08189_));
 sky130_as_sc_hs__or2_2 _38926_ (.A(_08188_),
    .B(_08189_),
    .Y(_08191_));
 sky130_as_sc_hs__and2_2 _38927_ (.A(_08190_),
    .B(_08191_),
    .Y(_08192_));
 sky130_as_sc_hs__and2_2 _38930_ (.A(net122),
    .B(net444),
    .Y(_08195_));
 sky130_as_sc_hs__and2_2 _38931_ (.A(net446),
    .B(net435),
    .Y(_08196_));
 sky130_as_sc_hs__or2_2 _38932_ (.A(_08195_),
    .B(_08196_),
    .Y(_08197_));
 sky130_as_sc_hs__and2_2 _38934_ (.A(_08197_),
    .B(_08198_),
    .Y(_08199_));
 sky130_as_sc_hs__and2_2 _38935_ (.A(_24729_),
    .B(_02481_),
    .Y(_08200_));
 sky130_as_sc_hs__or2_2 _38937_ (.A(_08199_),
    .B(_08200_),
    .Y(_08202_));
 sky130_as_sc_hs__and2_2 _38938_ (.A(_08201_),
    .B(_08202_),
    .Y(_08203_));
 sky130_as_sc_hs__or2_2 _38940_ (.A(_08194_),
    .B(_08203_),
    .Y(_08205_));
 sky130_as_sc_hs__and2_2 _38941_ (.A(_08204_),
    .B(_08205_),
    .Y(_08206_));
 sky130_as_sc_hs__or2_2 _38943_ (.A(_08193_),
    .B(_08206_),
    .Y(_08208_));
 sky130_as_sc_hs__and2_2 _38944_ (.A(_08207_),
    .B(_08208_),
    .Y(_08209_));
 sky130_as_sc_hs__or2_2 _38947_ (.A(_08209_),
    .B(_08210_),
    .Y(_08212_));
 sky130_as_sc_hs__and2_2 _38948_ (.A(_08211_),
    .B(_08212_),
    .Y(_08213_));
 sky130_as_sc_hs__or2_2 _38950_ (.A(_08192_),
    .B(_08213_),
    .Y(_08215_));
 sky130_as_sc_hs__and2_2 _38951_ (.A(_08214_),
    .B(_08215_),
    .Y(_08216_));
 sky130_as_sc_hs__or2_2 _38953_ (.A(_08184_),
    .B(_08216_),
    .Y(_08218_));
 sky130_as_sc_hs__and2_2 _38954_ (.A(_08217_),
    .B(_08218_),
    .Y(_08219_));
 sky130_as_sc_hs__or2_2 _38956_ (.A(_08183_),
    .B(_08219_),
    .Y(_08221_));
 sky130_as_sc_hs__and2_2 _38957_ (.A(_08220_),
    .B(_08221_),
    .Y(_08222_));
 sky130_as_sc_hs__and2_2 _38960_ (.A(net449),
    .B(net427),
    .Y(_08225_));
 sky130_as_sc_hs__and2_2 _38961_ (.A(net85),
    .B(net425),
    .Y(_08226_));
 sky130_as_sc_hs__or2_2 _38962_ (.A(_08225_),
    .B(_08226_),
    .Y(_08227_));
 sky130_as_sc_hs__and2_2 _38964_ (.A(_08227_),
    .B(_08228_),
    .Y(_08229_));
 sky130_as_sc_hs__and2_2 _38965_ (.A(net120),
    .B(net451),
    .Y(_08230_));
 sky130_as_sc_hs__or2_2 _38967_ (.A(_08229_),
    .B(_08230_),
    .Y(_08232_));
 sky130_as_sc_hs__and2_2 _38968_ (.A(_08231_),
    .B(_08232_),
    .Y(_08233_));
 sky130_as_sc_hs__and2_2 _38969_ (.A(_24527_),
    .B(net83),
    .Y(_08234_));
 sky130_as_sc_hs__and2_2 _38970_ (.A(net89),
    .B(net431),
    .Y(_08235_));
 sky130_as_sc_hs__or2_2 _38971_ (.A(_08234_),
    .B(_08235_),
    .Y(_08236_));
 sky130_as_sc_hs__and2_2 _38973_ (.A(_08236_),
    .B(_08237_),
    .Y(_08238_));
 sky130_as_sc_hs__and2_2 _38974_ (.A(net88),
    .B(net429),
    .Y(_08239_));
 sky130_as_sc_hs__or2_2 _38976_ (.A(_08238_),
    .B(_08239_),
    .Y(_08241_));
 sky130_as_sc_hs__and2_2 _38977_ (.A(_08240_),
    .B(_08241_),
    .Y(_08242_));
 sky130_as_sc_hs__or2_2 _38980_ (.A(_08242_),
    .B(_08243_),
    .Y(_08245_));
 sky130_as_sc_hs__and2_2 _38981_ (.A(_08244_),
    .B(_08245_),
    .Y(_08246_));
 sky130_as_sc_hs__or2_2 _38983_ (.A(_08233_),
    .B(_08246_),
    .Y(_08248_));
 sky130_as_sc_hs__and2_2 _38984_ (.A(_08247_),
    .B(_08248_),
    .Y(_08249_));
 sky130_as_sc_hs__or2_2 _38986_ (.A(_08224_),
    .B(_08249_),
    .Y(_08251_));
 sky130_as_sc_hs__and2_2 _38987_ (.A(_08250_),
    .B(_08251_),
    .Y(_08252_));
 sky130_as_sc_hs__or2_2 _38989_ (.A(_08223_),
    .B(_08252_),
    .Y(_08254_));
 sky130_as_sc_hs__and2_2 _38990_ (.A(_08253_),
    .B(_08254_),
    .Y(_08255_));
 sky130_as_sc_hs__and2_2 _38993_ (.A(net472),
    .B(net465),
    .Y(_08258_));
 sky130_as_sc_hs__and2_2 _38994_ (.A(net478),
    .B(net463),
    .Y(_08259_));
 sky130_as_sc_hs__or2_2 _38995_ (.A(_08258_),
    .B(_08259_),
    .Y(_08260_));
 sky130_as_sc_hs__and2_2 _38997_ (.A(_08260_),
    .B(_08261_),
    .Y(_08262_));
 sky130_as_sc_hs__and2_2 _38998_ (.A(net474),
    .B(net460),
    .Y(_08263_));
 sky130_as_sc_hs__or2_2 _39000_ (.A(_08262_),
    .B(_08263_),
    .Y(_08265_));
 sky130_as_sc_hs__and2_2 _39001_ (.A(_08264_),
    .B(_08265_),
    .Y(_08266_));
 sky130_as_sc_hs__or2_2 _39003_ (.A(_08257_),
    .B(_08266_),
    .Y(_08268_));
 sky130_as_sc_hs__and2_2 _39004_ (.A(_08267_),
    .B(_08268_),
    .Y(_08269_));
 sky130_as_sc_hs__or2_2 _39006_ (.A(_08256_),
    .B(_08269_),
    .Y(_08271_));
 sky130_as_sc_hs__and2_2 _39007_ (.A(_08270_),
    .B(_08271_),
    .Y(_08272_));
 sky130_as_sc_hs__and2_2 _39008_ (.A(net480),
    .B(net466),
    .Y(_08273_));
 sky130_as_sc_hs__and2_2 _39009_ (.A(net476),
    .B(net468),
    .Y(_08274_));
 sky130_as_sc_hs__or2_2 _39010_ (.A(_08273_),
    .B(_08274_),
    .Y(_08275_));
 sky130_as_sc_hs__and2_2 _39012_ (.A(_08275_),
    .B(_08276_),
    .Y(_08277_));
 sky130_as_sc_hs__and2_2 _39013_ (.A(net471),
    .B(net438),
    .Y(_08278_));
 sky130_as_sc_hs__or2_2 _39015_ (.A(_08277_),
    .B(_08278_),
    .Y(_08280_));
 sky130_as_sc_hs__and2_2 _39016_ (.A(_08279_),
    .B(_08280_),
    .Y(_08281_));
 sky130_as_sc_hs__and2_2 _39017_ (.A(net457),
    .B(net78),
    .Y(_08282_));
 sky130_as_sc_hs__or2_2 _39021_ (.A(_08283_),
    .B(_08284_),
    .Y(_08286_));
 sky130_as_sc_hs__and2_2 _39022_ (.A(_08285_),
    .B(_08286_),
    .Y(_08287_));
 sky130_as_sc_hs__or2_2 _39024_ (.A(_08282_),
    .B(_08287_),
    .Y(_08289_));
 sky130_as_sc_hs__and2_2 _39025_ (.A(_08288_),
    .B(_08289_),
    .Y(_08290_));
 sky130_as_sc_hs__or2_2 _39028_ (.A(_08290_),
    .B(_08291_),
    .Y(_08293_));
 sky130_as_sc_hs__and2_2 _39029_ (.A(_08292_),
    .B(_08293_),
    .Y(_08294_));
 sky130_as_sc_hs__or2_2 _39031_ (.A(_08281_),
    .B(_08294_),
    .Y(_08296_));
 sky130_as_sc_hs__and2_2 _39032_ (.A(_08295_),
    .B(_08296_),
    .Y(_08297_));
 sky130_as_sc_hs__or2_2 _39035_ (.A(_08297_),
    .B(_08298_),
    .Y(_08300_));
 sky130_as_sc_hs__and2_2 _39036_ (.A(_08299_),
    .B(_08300_),
    .Y(_08301_));
 sky130_as_sc_hs__or2_2 _39038_ (.A(_08272_),
    .B(_08301_),
    .Y(_08303_));
 sky130_as_sc_hs__and2_2 _39039_ (.A(_08302_),
    .B(_08303_),
    .Y(_08304_));
 sky130_as_sc_hs__or2_2 _39042_ (.A(_08304_),
    .B(_08305_),
    .Y(_08307_));
 sky130_as_sc_hs__and2_2 _39043_ (.A(_08306_),
    .B(_08307_),
    .Y(_08308_));
 sky130_as_sc_hs__or2_2 _39045_ (.A(_08255_),
    .B(_08308_),
    .Y(_08310_));
 sky130_as_sc_hs__and2_2 _39046_ (.A(_08309_),
    .B(_08310_),
    .Y(_08311_));
 sky130_as_sc_hs__or2_2 _39049_ (.A(_08311_),
    .B(_08312_),
    .Y(_08314_));
 sky130_as_sc_hs__and2_2 _39050_ (.A(_08313_),
    .B(_08314_),
    .Y(_08315_));
 sky130_as_sc_hs__or2_2 _39052_ (.A(_08222_),
    .B(_08315_),
    .Y(_08317_));
 sky130_as_sc_hs__and2_2 _39053_ (.A(_08316_),
    .B(_08317_),
    .Y(_08318_));
 sky130_as_sc_hs__or2_2 _39056_ (.A(_08318_),
    .B(_08319_),
    .Y(_08321_));
 sky130_as_sc_hs__and2_2 _39057_ (.A(_08320_),
    .B(_08321_),
    .Y(_08322_));
 sky130_as_sc_hs__or2_2 _39059_ (.A(_08182_),
    .B(_08322_),
    .Y(_08324_));
 sky130_as_sc_hs__and2_2 _39060_ (.A(_08323_),
    .B(_08324_),
    .Y(_08325_));
 sky130_as_sc_hs__or2_2 _39063_ (.A(_08325_),
    .B(_08326_),
    .Y(_08328_));
 sky130_as_sc_hs__and2_2 _39064_ (.A(_08327_),
    .B(_08328_),
    .Y(_08329_));
 sky130_as_sc_hs__or2_2 _39066_ (.A(_08150_),
    .B(_08329_),
    .Y(_08331_));
 sky130_as_sc_hs__and2_2 _39067_ (.A(_08330_),
    .B(_08331_),
    .Y(_08332_));
 sky130_as_sc_hs__or2_2 _39070_ (.A(_08332_),
    .B(_08333_),
    .Y(_08335_));
 sky130_as_sc_hs__and2_2 _39071_ (.A(_08334_),
    .B(_08335_),
    .Y(_08336_));
 sky130_as_sc_hs__or2_2 _39073_ (.A(_08149_),
    .B(_08336_),
    .Y(_08338_));
 sky130_as_sc_hs__and2_2 _39074_ (.A(_08337_),
    .B(_08338_),
    .Y(_08339_));
 sky130_as_sc_hs__or2_2 _39076_ (.A(_08148_),
    .B(_08339_),
    .Y(_08341_));
 sky130_as_sc_hs__and2_2 _39077_ (.A(_08340_),
    .B(_08341_),
    .Y(_08342_));
 sky130_as_sc_hs__and2_2 _39078_ (.A(_08058_),
    .B(_08067_),
    .Y(_08343_));
 sky130_as_sc_hs__or2_2 _39080_ (.A(_08342_),
    .B(_08343_),
    .Y(_08345_));
 sky130_as_sc_hs__and2_2 _39081_ (.A(_08344_),
    .B(_08345_),
    .Y(_08346_));
 sky130_as_sc_hs__nand3_2 _39082_ (.A(_07150_),
    .B(_07151_),
    .C(_08069_),
    .Y(_08347_));
 sky130_as_sc_hs__nor2_2 _39083_ (.A(_08070_),
    .B(_08347_),
    .Y(_08348_));
 sky130_as_sc_hs__or2_2 _39087_ (.A(_08346_),
    .B(_08350_),
    .Y(_08352_));
 sky130_as_sc_hs__nand3_2 _39088_ (.A(net142),
    .B(_08351_),
    .C(_08352_),
    .Y(_08353_));
 sky130_as_sc_hs__or2_2 _39089_ (.A(_05407_),
    .B(_05505_),
    .Y(_08354_));
 sky130_as_sc_hs__or2_2 _39091_ (.A(_05394_),
    .B(_08354_),
    .Y(_08356_));
 sky130_as_sc_hs__nand3_2 _39092_ (.A(net139),
    .B(_08355_),
    .C(_08356_),
    .Y(_08357_));
 sky130_as_sc_hs__or2_2 _39095_ (.A(_05757_),
    .B(_08359_),
    .Y(_08360_));
 sky130_as_sc_hs__and2_2 _39097_ (.A(_08360_),
    .B(_08361_),
    .Y(_08362_));
 sky130_as_sc_hs__or2_2 _39099_ (.A(_05757_),
    .B(_05860_),
    .Y(_08364_));
 sky130_as_sc_hs__nand3_2 _39102_ (.A(net118),
    .B(_08363_),
    .C(_08366_),
    .Y(_08367_));
 sky130_as_sc_hs__or2_2 _39108_ (.A(_05940_),
    .B(_07208_),
    .Y(_08373_));
 sky130_as_sc_hs__or2_2 _39109_ (.A(_05941_),
    .B(_07200_),
    .Y(_08374_));
 sky130_as_sc_hs__nand3_2 _39110_ (.A(_05935_),
    .B(_08373_),
    .C(_08374_),
    .Y(_08375_));
 sky130_as_sc_hs__and2_2 _39113_ (.A(_08376_),
    .B(_08377_),
    .Y(_08378_));
 sky130_as_sc_hs__or2_2 _39114_ (.A(_05935_),
    .B(_08378_),
    .Y(_08379_));
 sky130_as_sc_hs__or2_2 _39119_ (.A(_05935_),
    .B(_05961_),
    .Y(_08384_));
 sky130_as_sc_hs__and2_2 _39120_ (.A(_08383_),
    .B(_08384_),
    .Y(_08385_));
 sky130_as_sc_hs__nand3_2 _39121_ (.A(_05929_),
    .B(_08375_),
    .C(_08379_),
    .Y(_08386_));
 sky130_as_sc_hs__and2_2 _39124_ (.A(_05968_),
    .B(_08388_),
    .Y(_08389_));
 sky130_as_sc_hs__or2_2 _39125_ (.A(\tholin_riscv.div_res[6] ),
    .B(_08112_),
    .Y(_08390_));
 sky130_as_sc_hs__and2_2 _39126_ (.A(net414),
    .B(_08390_),
    .Y(_08391_));
 sky130_as_sc_hs__or2_2 _39127_ (.A(\tholin_riscv.div_res[7] ),
    .B(_08391_),
    .Y(_08392_));
 sky130_as_sc_hs__nand3_2 _39129_ (.A(net110),
    .B(_08392_),
    .C(_08393_),
    .Y(_08394_));
 sky130_as_sc_hs__nor2_2 _39133_ (.A(_05755_),
    .B(_06161_),
    .Y(_08398_));
 sky130_as_sc_hs__or2_2 _39134_ (.A(\tholin_riscv.div_shifter[38] ),
    .B(_08121_),
    .Y(_08399_));
 sky130_as_sc_hs__and2_2 _39135_ (.A(_21655_),
    .B(_08399_),
    .Y(_08400_));
 sky130_as_sc_hs__or2_2 _39137_ (.A(\tholin_riscv.div_shifter[39] ),
    .B(_08400_),
    .Y(_08402_));
 sky130_as_sc_hs__nand3_2 _39138_ (.A(net108),
    .B(_08401_),
    .C(_08402_),
    .Y(_08403_));
 sky130_as_sc_hs__and2_2 _39141_ (.A(_08404_),
    .B(_08405_),
    .Y(_08406_));
 sky130_as_sc_hs__nand3_2 _39142_ (.A(net412),
    .B(_08403_),
    .C(_08406_),
    .Y(_08407_));
 sky130_as_sc_hs__nor2_2 _39143_ (.A(_08398_),
    .B(_08407_),
    .Y(_08408_));
 sky130_as_sc_hs__nand3_2 _39144_ (.A(_08394_),
    .B(_08397_),
    .C(_08408_),
    .Y(_08409_));
 sky130_as_sc_hs__nor2_2 _39145_ (.A(_08389_),
    .B(_08409_),
    .Y(_08410_));
 sky130_as_sc_hs__and2_2 _39146_ (.A(_08372_),
    .B(_08410_),
    .Y(_08411_));
 sky130_as_sc_hs__and2_2 _39147_ (.A(_08367_),
    .B(_08411_),
    .Y(_08412_));
 sky130_as_sc_hs__nand3_2 _39148_ (.A(_08353_),
    .B(_08357_),
    .C(_08412_),
    .Y(_08413_));
 sky130_as_sc_hs__and2_2 _39150_ (.A(\tholin_riscv.PC[7] ),
    .B(_08136_),
    .Y(_08415_));
 sky130_as_sc_hs__nor2_2 _39151_ (.A(\tholin_riscv.PC[7] ),
    .B(_08136_),
    .Y(_08416_));
 sky130_as_sc_hs__nor2_2 _39152_ (.A(_08415_),
    .B(_08416_),
    .Y(_08417_));
 sky130_as_sc_hs__inv_2 _39153_ (.Y(_08418_),
    .A(_08417_));
 sky130_as_sc_hs__nand3_2 _39155_ (.A(_21569_),
    .B(_08414_),
    .C(_08419_),
    .Y(_08420_));
 sky130_as_sc_hs__nand3_2 _39156_ (.A(_21546_),
    .B(_08413_),
    .C(_08420_),
    .Y(_08421_));
 sky130_as_sc_hs__or2_2 _39161_ (.A(_19875_),
    .B(_19876_),
    .Y(_08425_));
 sky130_as_sc_hs__and2_2 _39162_ (.A(\tholin_riscv.load_funct ),
    .B(_08425_),
    .Y(_08426_));
 sky130_as_sc_hs__and2_2 _39164_ (.A(_08426_),
    .B(_08427_),
    .Y(_08428_));
 sky130_as_sc_hs__or2_2 _39165_ (.A(_19819_),
    .B(_08428_),
    .Y(_08429_));
 sky130_as_sc_hs__nand3_2 _39167_ (.A(_07866_),
    .B(_07867_),
    .C(_08158_),
    .Y(_08431_));
 sky130_as_sc_hs__and2_2 _39173_ (.A(net454),
    .B(net129),
    .Y(_08437_));
 sky130_as_sc_hs__or2_2 _39175_ (.A(_08436_),
    .B(_08437_),
    .Y(_08439_));
 sky130_as_sc_hs__or2_2 _39177_ (.A(_08168_),
    .B(_08440_),
    .Y(_08441_));
 sky130_as_sc_hs__and2_2 _39179_ (.A(_08441_),
    .B(_08442_),
    .Y(_08443_));
 sky130_as_sc_hs__and2_2 _39180_ (.A(net85),
    .B(net422),
    .Y(_08444_));
 sky130_as_sc_hs__and2_2 _39181_ (.A(_23624_),
    .B(net420),
    .Y(_08445_));
 sky130_as_sc_hs__and2_2 _39182_ (.A(_08444_),
    .B(_08445_),
    .Y(_08446_));
 sky130_as_sc_hs__or2_2 _39183_ (.A(_08444_),
    .B(_08445_),
    .Y(_08447_));
 sky130_as_sc_hs__nor2b_2 _39184_ (.A(_08446_),
    .Y(_08448_),
    .B(_08447_));
 sky130_as_sc_hs__and2_2 _39185_ (.A(_07865_),
    .B(_08158_),
    .Y(_08449_));
 sky130_as_sc_hs__or2_2 _39186_ (.A(_08156_),
    .B(_08449_),
    .Y(_08450_));
 sky130_as_sc_hs__or2_2 _39187_ (.A(_08448_),
    .B(_08450_),
    .Y(_08451_));
 sky130_as_sc_hs__and2_2 _39189_ (.A(_08451_),
    .B(_08452_),
    .Y(_08453_));
 sky130_as_sc_hs__or2_2 _39191_ (.A(_08443_),
    .B(_08453_),
    .Y(_08455_));
 sky130_as_sc_hs__and2_2 _39192_ (.A(_08454_),
    .B(_08455_),
    .Y(_08456_));
 sky130_as_sc_hs__or2_2 _39194_ (.A(_08435_),
    .B(_08456_),
    .Y(_08458_));
 sky130_as_sc_hs__and2_2 _39195_ (.A(_08457_),
    .B(_08458_),
    .Y(_08459_));
 sky130_as_sc_hs__or2_2 _39197_ (.A(_08434_),
    .B(_08459_),
    .Y(_08461_));
 sky130_as_sc_hs__and2_2 _39198_ (.A(_08460_),
    .B(_08461_),
    .Y(_08462_));
 sky130_as_sc_hs__and2_2 _39201_ (.A(_23674_),
    .B(net440),
    .Y(_08465_));
 sky130_as_sc_hs__and2_2 _39202_ (.A(net480),
    .B(net437),
    .Y(_08466_));
 sky130_as_sc_hs__and2_2 _39203_ (.A(_08465_),
    .B(_08466_),
    .Y(_08467_));
 sky130_as_sc_hs__or2_2 _39204_ (.A(_08465_),
    .B(_08466_),
    .Y(_08468_));
 sky130_as_sc_hs__nor2b_2 _39205_ (.A(_08467_),
    .Y(_08469_),
    .B(_08468_));
 sky130_as_sc_hs__and2_2 _39208_ (.A(net444),
    .B(net423),
    .Y(_08472_));
 sky130_as_sc_hs__and2_2 _39209_ (.A(net79),
    .B(net435),
    .Y(_08473_));
 sky130_as_sc_hs__or2_2 _39210_ (.A(_08472_),
    .B(_08473_),
    .Y(_08474_));
 sky130_as_sc_hs__and2_2 _39212_ (.A(_08474_),
    .B(_08475_),
    .Y(_08476_));
 sky130_as_sc_hs__and2_2 _39213_ (.A(_24729_),
    .B(net75),
    .Y(_08477_));
 sky130_as_sc_hs__or2_2 _39215_ (.A(_08476_),
    .B(_08477_),
    .Y(_08479_));
 sky130_as_sc_hs__and2_2 _39216_ (.A(_08478_),
    .B(_08479_),
    .Y(_08480_));
 sky130_as_sc_hs__or2_2 _39218_ (.A(_08471_),
    .B(_08480_),
    .Y(_08482_));
 sky130_as_sc_hs__and2_2 _39219_ (.A(_08481_),
    .B(_08482_),
    .Y(_08483_));
 sky130_as_sc_hs__or2_2 _39221_ (.A(_08470_),
    .B(_08483_),
    .Y(_08485_));
 sky130_as_sc_hs__and2_2 _39222_ (.A(_08484_),
    .B(_08485_),
    .Y(_08486_));
 sky130_as_sc_hs__or2_2 _39225_ (.A(_08486_),
    .B(_08487_),
    .Y(_08489_));
 sky130_as_sc_hs__and2_2 _39226_ (.A(_08488_),
    .B(_08489_),
    .Y(_08490_));
 sky130_as_sc_hs__or2_2 _39228_ (.A(_08469_),
    .B(_08490_),
    .Y(_08492_));
 sky130_as_sc_hs__and2_2 _39229_ (.A(_08491_),
    .B(_08492_),
    .Y(_08493_));
 sky130_as_sc_hs__or2_2 _39231_ (.A(_08464_),
    .B(_08493_),
    .Y(_08495_));
 sky130_as_sc_hs__and2_2 _39232_ (.A(_08494_),
    .B(_08495_),
    .Y(_08496_));
 sky130_as_sc_hs__or2_2 _39234_ (.A(_08463_),
    .B(_08496_),
    .Y(_08498_));
 sky130_as_sc_hs__and2_2 _39235_ (.A(_08497_),
    .B(_08498_),
    .Y(_08499_));
 sky130_as_sc_hs__and2_2 _39238_ (.A(net120),
    .B(net449),
    .Y(_08502_));
 sky130_as_sc_hs__and2_2 _39239_ (.A(net452),
    .B(net425),
    .Y(_08503_));
 sky130_as_sc_hs__or2_2 _39240_ (.A(_08502_),
    .B(_08503_),
    .Y(_08504_));
 sky130_as_sc_hs__and2_2 _39242_ (.A(_08504_),
    .B(_08505_),
    .Y(_08506_));
 sky130_as_sc_hs__and2_2 _39243_ (.A(net122),
    .B(net451),
    .Y(_08507_));
 sky130_as_sc_hs__or2_2 _39245_ (.A(_08506_),
    .B(_08507_),
    .Y(_08509_));
 sky130_as_sc_hs__and2_2 _39246_ (.A(_08508_),
    .B(_08509_),
    .Y(_08510_));
 sky130_as_sc_hs__and2_2 _39247_ (.A(_24527_),
    .B(net431),
    .Y(_08511_));
 sky130_as_sc_hs__and2_2 _39248_ (.A(net89),
    .B(net429),
    .Y(_08512_));
 sky130_as_sc_hs__or2_2 _39249_ (.A(_08511_),
    .B(_08512_),
    .Y(_08513_));
 sky130_as_sc_hs__and2_2 _39251_ (.A(_08513_),
    .B(_08514_),
    .Y(_08515_));
 sky130_as_sc_hs__and2_2 _39252_ (.A(net88),
    .B(net427),
    .Y(_08516_));
 sky130_as_sc_hs__or2_2 _39254_ (.A(_08515_),
    .B(_08516_),
    .Y(_08518_));
 sky130_as_sc_hs__and2_2 _39255_ (.A(_08517_),
    .B(_08518_),
    .Y(_08519_));
 sky130_as_sc_hs__or2_2 _39258_ (.A(_08519_),
    .B(_08520_),
    .Y(_08522_));
 sky130_as_sc_hs__and2_2 _39259_ (.A(_08521_),
    .B(_08522_),
    .Y(_08523_));
 sky130_as_sc_hs__or2_2 _39261_ (.A(_08510_),
    .B(_08523_),
    .Y(_08525_));
 sky130_as_sc_hs__and2_2 _39262_ (.A(_08524_),
    .B(_08525_),
    .Y(_08526_));
 sky130_as_sc_hs__or2_2 _39264_ (.A(_08501_),
    .B(_08526_),
    .Y(_08528_));
 sky130_as_sc_hs__and2_2 _39265_ (.A(_08527_),
    .B(_08528_),
    .Y(_08529_));
 sky130_as_sc_hs__or2_2 _39267_ (.A(_08500_),
    .B(_08529_),
    .Y(_08531_));
 sky130_as_sc_hs__and2_2 _39268_ (.A(_08530_),
    .B(_08531_),
    .Y(_08532_));
 sky130_as_sc_hs__and2_2 _39271_ (.A(net478),
    .B(net465),
    .Y(_08535_));
 sky130_as_sc_hs__and2_2 _39272_ (.A(net474),
    .B(net463),
    .Y(_08536_));
 sky130_as_sc_hs__or2_2 _39273_ (.A(_08535_),
    .B(_08536_),
    .Y(_08537_));
 sky130_as_sc_hs__and2_2 _39275_ (.A(_08537_),
    .B(_08538_),
    .Y(_08539_));
 sky130_as_sc_hs__and2_2 _39276_ (.A(net460),
    .B(net83),
    .Y(_08540_));
 sky130_as_sc_hs__or2_2 _39278_ (.A(_08539_),
    .B(_08540_),
    .Y(_08542_));
 sky130_as_sc_hs__and2_2 _39279_ (.A(_08541_),
    .B(_08542_),
    .Y(_08543_));
 sky130_as_sc_hs__or2_2 _39281_ (.A(_08534_),
    .B(_08543_),
    .Y(_08545_));
 sky130_as_sc_hs__and2_2 _39282_ (.A(_08544_),
    .B(_08545_),
    .Y(_08546_));
 sky130_as_sc_hs__or2_2 _39284_ (.A(_08533_),
    .B(_08546_),
    .Y(_08548_));
 sky130_as_sc_hs__and2_2 _39285_ (.A(_08547_),
    .B(_08548_),
    .Y(_08549_));
 sky130_as_sc_hs__and2_2 _39286_ (.A(net476),
    .B(net466),
    .Y(_08550_));
 sky130_as_sc_hs__and2_2 _39287_ (.A(net468),
    .B(net438),
    .Y(_08551_));
 sky130_as_sc_hs__or2_2 _39288_ (.A(_08550_),
    .B(_08551_),
    .Y(_08552_));
 sky130_as_sc_hs__and2_2 _39290_ (.A(_08552_),
    .B(_08553_),
    .Y(_08554_));
 sky130_as_sc_hs__and2_2 _39291_ (.A(net472),
    .B(net471),
    .Y(_08555_));
 sky130_as_sc_hs__or2_2 _39293_ (.A(_08554_),
    .B(_08555_),
    .Y(_08557_));
 sky130_as_sc_hs__and2_2 _39294_ (.A(_08556_),
    .B(_08557_),
    .Y(_08558_));
 sky130_as_sc_hs__and2_2 _39295_ (.A(net456),
    .B(net442),
    .Y(_08559_));
 sky130_as_sc_hs__and2_2 _39296_ (.A(_24545_),
    .B(net418),
    .Y(_08560_));
 sky130_as_sc_hs__and2_2 _39297_ (.A(net446),
    .B(_25035_),
    .Y(_08561_));
 sky130_as_sc_hs__or2_2 _39298_ (.A(_08560_),
    .B(_08561_),
    .Y(_08562_));
 sky130_as_sc_hs__and2_2 _39300_ (.A(_08562_),
    .B(_08563_),
    .Y(_08564_));
 sky130_as_sc_hs__or2_2 _39302_ (.A(_08559_),
    .B(_08564_),
    .Y(_08566_));
 sky130_as_sc_hs__and2_2 _39303_ (.A(_08565_),
    .B(_08566_),
    .Y(_08567_));
 sky130_as_sc_hs__or2_2 _39306_ (.A(_08567_),
    .B(_08568_),
    .Y(_08570_));
 sky130_as_sc_hs__and2_2 _39307_ (.A(_08569_),
    .B(_08570_),
    .Y(_08571_));
 sky130_as_sc_hs__or2_2 _39309_ (.A(_08558_),
    .B(_08571_),
    .Y(_08573_));
 sky130_as_sc_hs__and2_2 _39310_ (.A(_08572_),
    .B(_08573_),
    .Y(_08574_));
 sky130_as_sc_hs__or2_2 _39313_ (.A(_08574_),
    .B(_08575_),
    .Y(_08577_));
 sky130_as_sc_hs__and2_2 _39314_ (.A(_08576_),
    .B(_08577_),
    .Y(_08578_));
 sky130_as_sc_hs__or2_2 _39316_ (.A(_08549_),
    .B(_08578_),
    .Y(_08580_));
 sky130_as_sc_hs__and2_2 _39317_ (.A(_08579_),
    .B(_08580_),
    .Y(_08581_));
 sky130_as_sc_hs__or2_2 _39320_ (.A(_08581_),
    .B(_08582_),
    .Y(_08584_));
 sky130_as_sc_hs__and2_2 _39321_ (.A(_08583_),
    .B(_08584_),
    .Y(_08585_));
 sky130_as_sc_hs__or2_2 _39323_ (.A(_08532_),
    .B(_08585_),
    .Y(_08587_));
 sky130_as_sc_hs__and2_2 _39324_ (.A(_08586_),
    .B(_08587_),
    .Y(_08588_));
 sky130_as_sc_hs__or2_2 _39327_ (.A(_08588_),
    .B(_08589_),
    .Y(_08591_));
 sky130_as_sc_hs__and2_2 _39328_ (.A(_08590_),
    .B(_08591_),
    .Y(_08592_));
 sky130_as_sc_hs__or2_2 _39330_ (.A(_08499_),
    .B(_08592_),
    .Y(_08594_));
 sky130_as_sc_hs__and2_2 _39331_ (.A(_08593_),
    .B(_08594_),
    .Y(_08595_));
 sky130_as_sc_hs__or2_2 _39334_ (.A(_08595_),
    .B(_08596_),
    .Y(_08598_));
 sky130_as_sc_hs__and2_2 _39335_ (.A(_08597_),
    .B(_08598_),
    .Y(_08599_));
 sky130_as_sc_hs__or2_2 _39337_ (.A(_08462_),
    .B(_08599_),
    .Y(_08601_));
 sky130_as_sc_hs__and2_2 _39338_ (.A(_08600_),
    .B(_08601_),
    .Y(_08602_));
 sky130_as_sc_hs__or2_2 _39341_ (.A(_08602_),
    .B(_08603_),
    .Y(_08605_));
 sky130_as_sc_hs__and2_2 _39342_ (.A(_08604_),
    .B(_08605_),
    .Y(_08606_));
 sky130_as_sc_hs__or2_2 _39344_ (.A(_08433_),
    .B(_08606_),
    .Y(_08608_));
 sky130_as_sc_hs__and2_2 _39345_ (.A(_08607_),
    .B(_08608_),
    .Y(_08609_));
 sky130_as_sc_hs__or2_2 _39348_ (.A(_08609_),
    .B(_08610_),
    .Y(_08612_));
 sky130_as_sc_hs__and2_2 _39349_ (.A(_08611_),
    .B(_08612_),
    .Y(_08613_));
 sky130_as_sc_hs__or2_2 _39351_ (.A(_08432_),
    .B(_08613_),
    .Y(_08615_));
 sky130_as_sc_hs__and2_2 _39352_ (.A(_08614_),
    .B(_08615_),
    .Y(_08616_));
 sky130_as_sc_hs__or2_2 _39355_ (.A(_08616_),
    .B(_08617_),
    .Y(_08619_));
 sky130_as_sc_hs__and2_2 _39356_ (.A(_08618_),
    .B(_08619_),
    .Y(_08620_));
 sky130_as_sc_hs__and2_2 _39357_ (.A(_08060_),
    .B(_08342_),
    .Y(_08621_));
 sky130_as_sc_hs__and2_2 _39358_ (.A(_08064_),
    .B(_08621_),
    .Y(_08622_));
 sky130_as_sc_hs__and2_2 _39359_ (.A(_07480_),
    .B(_08622_),
    .Y(_08623_));
 sky130_as_sc_hs__nor2b_2 _39361_ (.A(_07479_),
    .Y(_08625_),
    .B(_08622_));
 sky130_as_sc_hs__nand2b_2 _39363_ (.B(_08341_),
    .Y(_08627_),
    .A(_08058_));
 sky130_as_sc_hs__nand3_2 _39364_ (.A(_08340_),
    .B(_08626_),
    .C(_08627_),
    .Y(_08628_));
 sky130_as_sc_hs__nor2_2 _39365_ (.A(_08625_),
    .B(_08628_),
    .Y(_08629_));
 sky130_as_sc_hs__and2_2 _39367_ (.A(_08620_),
    .B(_08630_),
    .Y(_08631_));
 sky130_as_sc_hs__nor2_2 _39369_ (.A(_08620_),
    .B(_08630_),
    .Y(_08633_));
 sky130_as_sc_hs__or2_2 _39370_ (.A(_08631_),
    .B(_08633_),
    .Y(_08634_));
 sky130_as_sc_hs__and2_2 _39371_ (.A(_08346_),
    .B(_08348_),
    .Y(_08635_));
 sky130_as_sc_hs__or2_2 _39372_ (.A(_05505_),
    .B(_08635_),
    .Y(_08636_));
 sky130_as_sc_hs__and2_2 _39373_ (.A(_05506_),
    .B(_08636_),
    .Y(_08637_));
 sky130_as_sc_hs__and2_2 _39374_ (.A(_08634_),
    .B(_08637_),
    .Y(_08638_));
 sky130_as_sc_hs__or2_2 _39375_ (.A(_08634_),
    .B(_08637_),
    .Y(_08639_));
 sky130_as_sc_hs__nor2_2 _39377_ (.A(_08638_),
    .B(_08640_),
    .Y(_08641_));
 sky130_as_sc_hs__or2_2 _39378_ (.A(_05408_),
    .B(_05505_),
    .Y(_08642_));
 sky130_as_sc_hs__or2_2 _39379_ (.A(_05392_),
    .B(_08642_),
    .Y(_08643_));
 sky130_as_sc_hs__nand3_2 _39381_ (.A(net139),
    .B(_08643_),
    .C(_08644_),
    .Y(_08645_));
 sky130_as_sc_hs__or2_2 _39382_ (.A(_05862_),
    .B(_05865_),
    .Y(_08646_));
 sky130_as_sc_hs__or2_2 _39385_ (.A(_05865_),
    .B(_08648_),
    .Y(_08649_));
 sky130_as_sc_hs__and2_2 _39387_ (.A(_08649_),
    .B(_08650_),
    .Y(_08651_));
 sky130_as_sc_hs__nand3_2 _39391_ (.A(net118),
    .B(_08653_),
    .C(_08654_),
    .Y(_08655_));
 sky130_as_sc_hs__or2_2 _39395_ (.A(_05935_),
    .B(_06103_),
    .Y(_08659_));
 sky130_as_sc_hs__nand3_2 _39397_ (.A(_05929_),
    .B(_08659_),
    .C(_08660_),
    .Y(_08661_));
 sky130_as_sc_hs__and2_2 _39400_ (.A(_05968_),
    .B(_08663_),
    .Y(_08664_));
 sky130_as_sc_hs__or2_2 _39401_ (.A(\tholin_riscv.div_res[7] ),
    .B(_08390_),
    .Y(_08665_));
 sky130_as_sc_hs__and2_2 _39402_ (.A(net414),
    .B(_08665_),
    .Y(_08666_));
 sky130_as_sc_hs__or2_2 _39403_ (.A(\tholin_riscv.div_res[8] ),
    .B(_08666_),
    .Y(_08667_));
 sky130_as_sc_hs__nand3_2 _39405_ (.A(net110),
    .B(_08667_),
    .C(_08668_),
    .Y(_08669_));
 sky130_as_sc_hs__nor2_2 _39409_ (.A(_05863_),
    .B(_06161_),
    .Y(_08673_));
 sky130_as_sc_hs__or2_2 _39410_ (.A(\tholin_riscv.div_shifter[39] ),
    .B(_08399_),
    .Y(_08674_));
 sky130_as_sc_hs__and2_2 _39411_ (.A(_21655_),
    .B(_08674_),
    .Y(_08675_));
 sky130_as_sc_hs__or2_2 _39413_ (.A(\tholin_riscv.div_shifter[40] ),
    .B(_08675_),
    .Y(_08677_));
 sky130_as_sc_hs__nand3_2 _39414_ (.A(net108),
    .B(_08676_),
    .C(_08677_),
    .Y(_08678_));
 sky130_as_sc_hs__and2_2 _39417_ (.A(_08679_),
    .B(_08680_),
    .Y(_08681_));
 sky130_as_sc_hs__nand3_2 _39418_ (.A(net412),
    .B(_08678_),
    .C(_08681_),
    .Y(_08682_));
 sky130_as_sc_hs__nor2_2 _39419_ (.A(_08673_),
    .B(_08682_),
    .Y(_08683_));
 sky130_as_sc_hs__nand3_2 _39420_ (.A(_08669_),
    .B(_08672_),
    .C(_08683_),
    .Y(_08684_));
 sky130_as_sc_hs__nor2_2 _39421_ (.A(_08664_),
    .B(_08684_),
    .Y(_08685_));
 sky130_as_sc_hs__and2_2 _39422_ (.A(_08658_),
    .B(_08685_),
    .Y(_08686_));
 sky130_as_sc_hs__nand3_2 _39423_ (.A(_08645_),
    .B(_08655_),
    .C(_08686_),
    .Y(_08687_));
 sky130_as_sc_hs__or2_2 _39424_ (.A(_08641_),
    .B(_08687_),
    .Y(_08688_));
 sky130_as_sc_hs__and2_2 _39426_ (.A(\tholin_riscv.PC[8] ),
    .B(_08415_),
    .Y(_08690_));
 sky130_as_sc_hs__nor2_2 _39427_ (.A(\tholin_riscv.PC[8] ),
    .B(_08415_),
    .Y(_08691_));
 sky130_as_sc_hs__nor2_2 _39428_ (.A(_08690_),
    .B(_08691_),
    .Y(_08692_));
 sky130_as_sc_hs__inv_2 _39429_ (.Y(_08693_),
    .A(_08692_));
 sky130_as_sc_hs__nand3_2 _39431_ (.A(_21569_),
    .B(_08689_),
    .C(_08694_),
    .Y(_08695_));
 sky130_as_sc_hs__nand3_2 _39432_ (.A(_21546_),
    .B(_08688_),
    .C(_08695_),
    .Y(_08696_));
 sky130_as_sc_hs__or2_2 _39437_ (.A(_19827_),
    .B(_08428_),
    .Y(_08700_));
 sky130_as_sc_hs__and2_2 _39442_ (.A(net85),
    .B(net129),
    .Y(_08705_));
 sky130_as_sc_hs__or2_2 _39444_ (.A(_08467_),
    .B(_08705_),
    .Y(_08707_));
 sky130_as_sc_hs__or2_2 _39446_ (.A(_08438_),
    .B(_08708_),
    .Y(_08709_));
 sky130_as_sc_hs__and2_2 _39448_ (.A(_08709_),
    .B(_08710_),
    .Y(_08711_));
 sky130_as_sc_hs__and2_2 _39449_ (.A(net452),
    .B(net422),
    .Y(_08712_));
 sky130_as_sc_hs__and2_2 _39450_ (.A(_23624_),
    .B(net75),
    .Y(_08713_));
 sky130_as_sc_hs__or2_2 _39451_ (.A(_08712_),
    .B(_08713_),
    .Y(_08714_));
 sky130_as_sc_hs__and2_2 _39453_ (.A(_08714_),
    .B(_08715_),
    .Y(_08716_));
 sky130_as_sc_hs__and2_2 _39454_ (.A(_08156_),
    .B(_08448_),
    .Y(_08717_));
 sky130_as_sc_hs__or2_2 _39455_ (.A(_08446_),
    .B(_08717_),
    .Y(_08718_));
 sky130_as_sc_hs__or2_2 _39456_ (.A(_08716_),
    .B(_08718_),
    .Y(_08719_));
 sky130_as_sc_hs__and2_2 _39458_ (.A(_08719_),
    .B(_08720_),
    .Y(_08721_));
 sky130_as_sc_hs__or2_2 _39460_ (.A(_08711_),
    .B(_08721_),
    .Y(_08723_));
 sky130_as_sc_hs__and2_2 _39461_ (.A(_08722_),
    .B(_08723_),
    .Y(_08724_));
 sky130_as_sc_hs__or2_2 _39463_ (.A(_08704_),
    .B(_08724_),
    .Y(_08726_));
 sky130_as_sc_hs__and2_2 _39464_ (.A(_08725_),
    .B(_08726_),
    .Y(_08727_));
 sky130_as_sc_hs__or2_2 _39466_ (.A(_08703_),
    .B(_08727_),
    .Y(_08729_));
 sky130_as_sc_hs__and2_2 _39467_ (.A(_08728_),
    .B(_08729_),
    .Y(_08730_));
 sky130_as_sc_hs__and2_2 _39470_ (.A(net481),
    .B(net440),
    .Y(_08733_));
 sky130_as_sc_hs__and2_2 _39471_ (.A(net476),
    .B(net436),
    .Y(_08734_));
 sky130_as_sc_hs__and2_2 _39472_ (.A(_08733_),
    .B(_08734_),
    .Y(_08735_));
 sky130_as_sc_hs__or2_2 _39473_ (.A(_08733_),
    .B(_08734_),
    .Y(_08736_));
 sky130_as_sc_hs__nor2b_2 _39474_ (.A(_08735_),
    .Y(_08737_),
    .B(_08736_));
 sky130_as_sc_hs__and2_2 _39477_ (.A(net442),
    .B(net434),
    .Y(_08740_));
 sky130_as_sc_hs__and2_2 _39478_ (.A(net444),
    .B(net420),
    .Y(_08741_));
 sky130_as_sc_hs__or2_2 _39480_ (.A(_08740_),
    .B(_08741_),
    .Y(_08743_));
 sky130_as_sc_hs__and2_2 _39481_ (.A(_08742_),
    .B(_08743_),
    .Y(_08744_));
 sky130_as_sc_hs__or2_2 _39483_ (.A(_08739_),
    .B(_08744_),
    .Y(_08746_));
 sky130_as_sc_hs__and2_2 _39484_ (.A(_08745_),
    .B(_08746_),
    .Y(_08747_));
 sky130_as_sc_hs__or2_2 _39486_ (.A(_08738_),
    .B(_08747_),
    .Y(_08749_));
 sky130_as_sc_hs__and2_2 _39487_ (.A(_08748_),
    .B(_08749_),
    .Y(_08750_));
 sky130_as_sc_hs__or2_2 _39490_ (.A(_08750_),
    .B(_08751_),
    .Y(_08753_));
 sky130_as_sc_hs__and2_2 _39491_ (.A(_08752_),
    .B(_08753_),
    .Y(_08754_));
 sky130_as_sc_hs__or2_2 _39493_ (.A(_08737_),
    .B(_08754_),
    .Y(_08756_));
 sky130_as_sc_hs__and2_2 _39494_ (.A(_08755_),
    .B(_08756_),
    .Y(_08757_));
 sky130_as_sc_hs__or2_2 _39496_ (.A(_08732_),
    .B(_08757_),
    .Y(_08759_));
 sky130_as_sc_hs__and2_2 _39497_ (.A(_08758_),
    .B(_08759_),
    .Y(_08760_));
 sky130_as_sc_hs__or2_2 _39499_ (.A(_08731_),
    .B(_08760_),
    .Y(_08762_));
 sky130_as_sc_hs__and2_2 _39500_ (.A(_08761_),
    .B(_08762_),
    .Y(_08763_));
 sky130_as_sc_hs__or2_2 _39506_ (.A(_08766_),
    .B(_08767_),
    .Y(_08769_));
 sky130_as_sc_hs__and2_2 _39507_ (.A(_08768_),
    .B(_08769_),
    .Y(_08770_));
 sky130_as_sc_hs__and2_2 _39508_ (.A(net451),
    .B(net424),
    .Y(_08771_));
 sky130_as_sc_hs__or2_2 _39510_ (.A(_08770_),
    .B(_08771_),
    .Y(_08773_));
 sky130_as_sc_hs__and2_2 _39511_ (.A(_08772_),
    .B(_08773_),
    .Y(_08774_));
 sky130_as_sc_hs__and2_2 _39512_ (.A(_24527_),
    .B(net429),
    .Y(_08775_));
 sky130_as_sc_hs__and2_2 _39513_ (.A(net89),
    .B(net427),
    .Y(_08776_));
 sky130_as_sc_hs__or2_2 _39514_ (.A(_08775_),
    .B(_08776_),
    .Y(_08777_));
 sky130_as_sc_hs__and2_2 _39516_ (.A(_08777_),
    .B(_08778_),
    .Y(_08779_));
 sky130_as_sc_hs__and2_2 _39517_ (.A(net120),
    .B(net88),
    .Y(_08780_));
 sky130_as_sc_hs__or2_2 _39519_ (.A(_08779_),
    .B(_08780_),
    .Y(_08782_));
 sky130_as_sc_hs__and2_2 _39520_ (.A(_08781_),
    .B(_08782_),
    .Y(_08783_));
 sky130_as_sc_hs__or2_2 _39523_ (.A(_08783_),
    .B(_08784_),
    .Y(_08786_));
 sky130_as_sc_hs__and2_2 _39524_ (.A(_08785_),
    .B(_08786_),
    .Y(_08787_));
 sky130_as_sc_hs__or2_2 _39526_ (.A(_08774_),
    .B(_08787_),
    .Y(_08789_));
 sky130_as_sc_hs__and2_2 _39527_ (.A(_08788_),
    .B(_08789_),
    .Y(_08790_));
 sky130_as_sc_hs__or2_2 _39529_ (.A(_08765_),
    .B(_08790_),
    .Y(_08792_));
 sky130_as_sc_hs__and2_2 _39530_ (.A(_08791_),
    .B(_08792_),
    .Y(_08793_));
 sky130_as_sc_hs__or2_2 _39532_ (.A(_08764_),
    .B(_08793_),
    .Y(_08795_));
 sky130_as_sc_hs__and2_2 _39533_ (.A(_08794_),
    .B(_08795_),
    .Y(_08796_));
 sky130_as_sc_hs__and2_2 _39536_ (.A(net474),
    .B(net465),
    .Y(_08799_));
 sky130_as_sc_hs__and2_2 _39537_ (.A(net463),
    .B(net83),
    .Y(_08800_));
 sky130_as_sc_hs__or2_2 _39538_ (.A(_08799_),
    .B(_08800_),
    .Y(_08801_));
 sky130_as_sc_hs__and2_2 _39540_ (.A(_08801_),
    .B(_08802_),
    .Y(_08803_));
 sky130_as_sc_hs__and2_2 _39541_ (.A(net460),
    .B(net431),
    .Y(_08804_));
 sky130_as_sc_hs__or2_2 _39543_ (.A(_08803_),
    .B(_08804_),
    .Y(_08806_));
 sky130_as_sc_hs__and2_2 _39544_ (.A(_08805_),
    .B(_08806_),
    .Y(_08807_));
 sky130_as_sc_hs__or2_2 _39546_ (.A(_08798_),
    .B(_08807_),
    .Y(_08809_));
 sky130_as_sc_hs__and2_2 _39547_ (.A(_08808_),
    .B(_08809_),
    .Y(_08810_));
 sky130_as_sc_hs__or2_2 _39549_ (.A(_08797_),
    .B(_08810_),
    .Y(_08812_));
 sky130_as_sc_hs__and2_2 _39550_ (.A(_08811_),
    .B(_08812_),
    .Y(_08813_));
 sky130_as_sc_hs__and2_2 _39551_ (.A(net466),
    .B(net438),
    .Y(_08814_));
 sky130_as_sc_hs__and2_2 _39552_ (.A(net472),
    .B(net468),
    .Y(_08815_));
 sky130_as_sc_hs__or2_2 _39553_ (.A(_08814_),
    .B(_08815_),
    .Y(_08816_));
 sky130_as_sc_hs__and2_2 _39555_ (.A(_08816_),
    .B(_08817_),
    .Y(_08818_));
 sky130_as_sc_hs__and2_2 _39556_ (.A(net478),
    .B(net471),
    .Y(_08819_));
 sky130_as_sc_hs__or2_2 _39558_ (.A(_08818_),
    .B(_08819_),
    .Y(_08821_));
 sky130_as_sc_hs__and2_2 _39559_ (.A(_08820_),
    .B(_08821_),
    .Y(_08822_));
 sky130_as_sc_hs__and2_2 _39560_ (.A(net454),
    .B(net418),
    .Y(_08823_));
 sky130_as_sc_hs__and2_2 _39561_ (.A(net78),
    .B(_25035_),
    .Y(_08824_));
 sky130_as_sc_hs__or2_2 _39562_ (.A(_08823_),
    .B(_08824_),
    .Y(_08825_));
 sky130_as_sc_hs__and2_2 _39564_ (.A(_08825_),
    .B(_08826_),
    .Y(_08827_));
 sky130_as_sc_hs__and2_2 _39565_ (.A(_23674_),
    .B(net456),
    .Y(_08828_));
 sky130_as_sc_hs__or2_2 _39567_ (.A(_08827_),
    .B(_08828_),
    .Y(_08830_));
 sky130_as_sc_hs__and2_2 _39568_ (.A(_08829_),
    .B(_08830_),
    .Y(_08831_));
 sky130_as_sc_hs__or2_2 _39571_ (.A(_08831_),
    .B(_08832_),
    .Y(_08834_));
 sky130_as_sc_hs__and2_2 _39572_ (.A(_08833_),
    .B(_08834_),
    .Y(_08835_));
 sky130_as_sc_hs__or2_2 _39574_ (.A(_08822_),
    .B(_08835_),
    .Y(_08837_));
 sky130_as_sc_hs__and2_2 _39575_ (.A(_08836_),
    .B(_08837_),
    .Y(_08838_));
 sky130_as_sc_hs__or2_2 _39578_ (.A(_08838_),
    .B(_08839_),
    .Y(_08841_));
 sky130_as_sc_hs__and2_2 _39579_ (.A(_08840_),
    .B(_08841_),
    .Y(_08842_));
 sky130_as_sc_hs__or2_2 _39581_ (.A(_08813_),
    .B(_08842_),
    .Y(_08844_));
 sky130_as_sc_hs__and2_2 _39582_ (.A(_08843_),
    .B(_08844_),
    .Y(_08845_));
 sky130_as_sc_hs__or2_2 _39585_ (.A(_08845_),
    .B(_08846_),
    .Y(_08848_));
 sky130_as_sc_hs__and2_2 _39586_ (.A(_08847_),
    .B(_08848_),
    .Y(_08849_));
 sky130_as_sc_hs__or2_2 _39588_ (.A(_08796_),
    .B(_08849_),
    .Y(_08851_));
 sky130_as_sc_hs__and2_2 _39589_ (.A(_08850_),
    .B(_08851_),
    .Y(_08852_));
 sky130_as_sc_hs__or2_2 _39592_ (.A(_08852_),
    .B(_08853_),
    .Y(_08855_));
 sky130_as_sc_hs__and2_2 _39593_ (.A(_08854_),
    .B(_08855_),
    .Y(_08856_));
 sky130_as_sc_hs__or2_2 _39595_ (.A(_08763_),
    .B(_08856_),
    .Y(_08858_));
 sky130_as_sc_hs__and2_2 _39596_ (.A(_08857_),
    .B(_08858_),
    .Y(_08859_));
 sky130_as_sc_hs__or2_2 _39599_ (.A(_08859_),
    .B(_08860_),
    .Y(_08862_));
 sky130_as_sc_hs__and2_2 _39600_ (.A(_08861_),
    .B(_08862_),
    .Y(_08863_));
 sky130_as_sc_hs__or2_2 _39602_ (.A(_08730_),
    .B(_08863_),
    .Y(_08865_));
 sky130_as_sc_hs__and2_2 _39603_ (.A(_08864_),
    .B(_08865_),
    .Y(_08866_));
 sky130_as_sc_hs__or2_2 _39606_ (.A(_08866_),
    .B(_08867_),
    .Y(_08869_));
 sky130_as_sc_hs__and2_2 _39607_ (.A(_08868_),
    .B(_08869_),
    .Y(_08870_));
 sky130_as_sc_hs__or2_2 _39609_ (.A(_08702_),
    .B(_08870_),
    .Y(_08872_));
 sky130_as_sc_hs__and2_2 _39610_ (.A(_08871_),
    .B(_08872_),
    .Y(_08873_));
 sky130_as_sc_hs__or2_2 _39613_ (.A(_08873_),
    .B(_08874_),
    .Y(_08876_));
 sky130_as_sc_hs__and2_2 _39614_ (.A(_08875_),
    .B(_08876_),
    .Y(_08877_));
 sky130_as_sc_hs__and2_2 _39615_ (.A(_08448_),
    .B(_08449_),
    .Y(_08878_));
 sky130_as_sc_hs__or2_2 _39617_ (.A(_08877_),
    .B(_08878_),
    .Y(_08880_));
 sky130_as_sc_hs__and2_2 _39618_ (.A(_08879_),
    .B(_08880_),
    .Y(_08881_));
 sky130_as_sc_hs__or2_2 _39621_ (.A(_08881_),
    .B(_08882_),
    .Y(_08884_));
 sky130_as_sc_hs__and2_2 _39622_ (.A(_08883_),
    .B(_08884_),
    .Y(_08885_));
 sky130_as_sc_hs__or2_2 _39624_ (.A(_08885_),
    .B(_08886_),
    .Y(_08887_));
 sky130_as_sc_hs__or2_2 _39627_ (.A(_05505_),
    .B(_08638_),
    .Y(_08890_));
 sky130_as_sc_hs__or2_2 _39628_ (.A(_08889_),
    .B(_08890_),
    .Y(_08891_));
 sky130_as_sc_hs__nand3_2 _39630_ (.A(net142),
    .B(_08891_),
    .C(_08892_),
    .Y(_08893_));
 sky130_as_sc_hs__or2_2 _39631_ (.A(_05409_),
    .B(_05505_),
    .Y(_08894_));
 sky130_as_sc_hs__or2_2 _39633_ (.A(_05390_),
    .B(_08894_),
    .Y(_08896_));
 sky130_as_sc_hs__nand3_2 _39634_ (.A(net139),
    .B(_08895_),
    .C(_08896_),
    .Y(_08897_));
 sky130_as_sc_hs__or2_2 _39638_ (.A(_05737_),
    .B(_08899_),
    .Y(_08901_));
 sky130_as_sc_hs__nand3_2 _39644_ (.A(_06523_),
    .B(_08903_),
    .C(_08906_),
    .Y(_08907_));
 sky130_as_sc_hs__or2_2 _39645_ (.A(_05936_),
    .B(_06474_),
    .Y(_08908_));
 sky130_as_sc_hs__or2_2 _39646_ (.A(_05935_),
    .B(_06517_),
    .Y(_08909_));
 sky130_as_sc_hs__nand3_2 _39647_ (.A(_05929_),
    .B(_08908_),
    .C(_08909_),
    .Y(_08910_));
 sky130_as_sc_hs__or2_2 _39648_ (.A(_05929_),
    .B(_08108_),
    .Y(_08911_));
 sky130_as_sc_hs__and2_2 _39649_ (.A(_08910_),
    .B(_08911_),
    .Y(_08912_));
 sky130_as_sc_hs__and2_2 _39653_ (.A(_05926_),
    .B(_08915_),
    .Y(_08916_));
 sky130_as_sc_hs__or2_2 _39654_ (.A(\tholin_riscv.div_res[8] ),
    .B(_08665_),
    .Y(_08917_));
 sky130_as_sc_hs__and2_2 _39655_ (.A(net415),
    .B(_08917_),
    .Y(_08918_));
 sky130_as_sc_hs__or2_2 _39656_ (.A(\tholin_riscv.div_res[9] ),
    .B(_08918_),
    .Y(_08919_));
 sky130_as_sc_hs__nand3_2 _39658_ (.A(net111),
    .B(_08919_),
    .C(_08920_),
    .Y(_08921_));
 sky130_as_sc_hs__or2_2 _39662_ (.A(\tholin_riscv.div_shifter[40] ),
    .B(_08674_),
    .Y(_08925_));
 sky130_as_sc_hs__and2_2 _39663_ (.A(_21655_),
    .B(_08925_),
    .Y(_08926_));
 sky130_as_sc_hs__or2_2 _39665_ (.A(\tholin_riscv.div_shifter[41] ),
    .B(_08926_),
    .Y(_08928_));
 sky130_as_sc_hs__nand3_2 _39666_ (.A(net108),
    .B(_08927_),
    .C(_08928_),
    .Y(_08929_));
 sky130_as_sc_hs__nor2_2 _39667_ (.A(_05735_),
    .B(_06161_),
    .Y(_08930_));
 sky130_as_sc_hs__and2_2 _39670_ (.A(_08931_),
    .B(_08932_),
    .Y(_08933_));
 sky130_as_sc_hs__nand3_2 _39671_ (.A(net412),
    .B(_08929_),
    .C(_08933_),
    .Y(_08934_));
 sky130_as_sc_hs__nor2_2 _39672_ (.A(_08930_),
    .B(_08934_),
    .Y(_08935_));
 sky130_as_sc_hs__nand3_2 _39673_ (.A(_08921_),
    .B(_08924_),
    .C(_08935_),
    .Y(_08936_));
 sky130_as_sc_hs__nor2_2 _39674_ (.A(_08916_),
    .B(_08936_),
    .Y(_08937_));
 sky130_as_sc_hs__and2_2 _39675_ (.A(_08913_),
    .B(_08937_),
    .Y(_08938_));
 sky130_as_sc_hs__and2_2 _39676_ (.A(_08907_),
    .B(_08938_),
    .Y(_08939_));
 sky130_as_sc_hs__nand3_2 _39677_ (.A(_08893_),
    .B(_08897_),
    .C(_08939_),
    .Y(_08940_));
 sky130_as_sc_hs__and2_2 _39678_ (.A(\tholin_riscv.PC[9] ),
    .B(_08690_),
    .Y(_08941_));
 sky130_as_sc_hs__nor2_2 _39679_ (.A(\tholin_riscv.PC[9] ),
    .B(_08690_),
    .Y(_08942_));
 sky130_as_sc_hs__nor2_2 _39680_ (.A(_08941_),
    .B(_08942_),
    .Y(_08943_));
 sky130_as_sc_hs__nand3_2 _39683_ (.A(_21569_),
    .B(_08944_),
    .C(_08945_),
    .Y(_08946_));
 sky130_as_sc_hs__nand3_2 _39684_ (.A(_21546_),
    .B(_08940_),
    .C(_08946_),
    .Y(_08947_));
 sky130_as_sc_hs__or2_2 _39689_ (.A(_19835_),
    .B(_08428_),
    .Y(_08951_));
 sky130_as_sc_hs__and2_2 _39694_ (.A(_08446_),
    .B(_08716_),
    .Y(_08956_));
 sky130_as_sc_hs__nand3_2 _39695_ (.A(net446),
    .B(_08712_),
    .C(_08713_),
    .Y(_08957_));
 sky130_as_sc_hs__and2_2 _39698_ (.A(_08957_),
    .B(_08959_),
    .Y(_08960_));
 sky130_as_sc_hs__or2_2 _39700_ (.A(_08956_),
    .B(_08960_),
    .Y(_08962_));
 sky130_as_sc_hs__and2_2 _39701_ (.A(_08961_),
    .B(_08962_),
    .Y(_08963_));
 sky130_as_sc_hs__and2_2 _39702_ (.A(net452),
    .B(net129),
    .Y(_08964_));
 sky130_as_sc_hs__or2_2 _39704_ (.A(_08735_),
    .B(_08964_),
    .Y(_08966_));
 sky130_as_sc_hs__or2_2 _39706_ (.A(_08706_),
    .B(_08967_),
    .Y(_08968_));
 sky130_as_sc_hs__and2_2 _39708_ (.A(_08968_),
    .B(_08969_),
    .Y(_08970_));
 sky130_as_sc_hs__or2_2 _39710_ (.A(_08963_),
    .B(_08970_),
    .Y(_08972_));
 sky130_as_sc_hs__and2_2 _39711_ (.A(_08971_),
    .B(_08972_),
    .Y(_08973_));
 sky130_as_sc_hs__or2_2 _39713_ (.A(_08955_),
    .B(_08973_),
    .Y(_08975_));
 sky130_as_sc_hs__and2_2 _39714_ (.A(_08974_),
    .B(_08975_),
    .Y(_08976_));
 sky130_as_sc_hs__or2_2 _39716_ (.A(_08954_),
    .B(_08976_),
    .Y(_08978_));
 sky130_as_sc_hs__and2_2 _39717_ (.A(_08977_),
    .B(_08978_),
    .Y(_08979_));
 sky130_as_sc_hs__and2_2 _39720_ (.A(net476),
    .B(net440),
    .Y(_08982_));
 sky130_as_sc_hs__and2_2 _39721_ (.A(net438),
    .B(net436),
    .Y(_08983_));
 sky130_as_sc_hs__and2_2 _39722_ (.A(_08982_),
    .B(_08983_),
    .Y(_08984_));
 sky130_as_sc_hs__or2_2 _39723_ (.A(_08982_),
    .B(_08983_),
    .Y(_08985_));
 sky130_as_sc_hs__nor2b_2 _39724_ (.A(_08984_),
    .Y(_08986_),
    .B(_08985_));
 sky130_as_sc_hs__and2_2 _39726_ (.A(_23674_),
    .B(net434),
    .Y(_08988_));
 sky130_as_sc_hs__and2_2 _39727_ (.A(net444),
    .B(net74),
    .Y(_08989_));
 sky130_as_sc_hs__or2_2 _39729_ (.A(_08988_),
    .B(_08989_),
    .Y(_08991_));
 sky130_as_sc_hs__and2_2 _39730_ (.A(_08990_),
    .B(_08991_),
    .Y(_08992_));
 sky130_as_sc_hs__or2_2 _39732_ (.A(_08987_),
    .B(_08992_),
    .Y(_08994_));
 sky130_as_sc_hs__or2_2 _39734_ (.A(_08742_),
    .B(_08995_),
    .Y(_08996_));
 sky130_as_sc_hs__and2_2 _39736_ (.A(_08996_),
    .B(_08997_),
    .Y(_08998_));
 sky130_as_sc_hs__or2_2 _39739_ (.A(_08998_),
    .B(_08999_),
    .Y(_09001_));
 sky130_as_sc_hs__and2_2 _39740_ (.A(_09000_),
    .B(_09001_),
    .Y(_09002_));
 sky130_as_sc_hs__or2_2 _39742_ (.A(_08986_),
    .B(_09002_),
    .Y(_09004_));
 sky130_as_sc_hs__and2_2 _39743_ (.A(_09003_),
    .B(_09004_),
    .Y(_09005_));
 sky130_as_sc_hs__or2_2 _39745_ (.A(_08981_),
    .B(_09005_),
    .Y(_09007_));
 sky130_as_sc_hs__and2_2 _39746_ (.A(_09006_),
    .B(_09007_),
    .Y(_09008_));
 sky130_as_sc_hs__or2_2 _39748_ (.A(_08980_),
    .B(_09008_),
    .Y(_09010_));
 sky130_as_sc_hs__and2_2 _39749_ (.A(_09009_),
    .B(_09010_),
    .Y(_09011_));
 sky130_as_sc_hs__and2_2 _39752_ (.A(net449),
    .B(net424),
    .Y(_09014_));
 sky130_as_sc_hs__and2_2 _39753_ (.A(net78),
    .B(net426),
    .Y(_09015_));
 sky130_as_sc_hs__or2_2 _39754_ (.A(_09014_),
    .B(_09015_),
    .Y(_09016_));
 sky130_as_sc_hs__and2_2 _39756_ (.A(_09016_),
    .B(_09017_),
    .Y(_09018_));
 sky130_as_sc_hs__and2_2 _39757_ (.A(net451),
    .B(net420),
    .Y(_09019_));
 sky130_as_sc_hs__or2_2 _39759_ (.A(_09018_),
    .B(_09019_),
    .Y(_09021_));
 sky130_as_sc_hs__and2_2 _39760_ (.A(_09020_),
    .B(_09021_),
    .Y(_09022_));
 sky130_as_sc_hs__or2_2 _39764_ (.A(_09023_),
    .B(_09024_),
    .Y(_09026_));
 sky130_as_sc_hs__and2_2 _39765_ (.A(_09025_),
    .B(_09026_),
    .Y(_09027_));
 sky130_as_sc_hs__and2_2 _39766_ (.A(net123),
    .B(net88),
    .Y(_09028_));
 sky130_as_sc_hs__or2_2 _39768_ (.A(_09027_),
    .B(_09028_),
    .Y(_09030_));
 sky130_as_sc_hs__and2_2 _39769_ (.A(_09029_),
    .B(_09030_),
    .Y(_09031_));
 sky130_as_sc_hs__or2_2 _39772_ (.A(_09031_),
    .B(_09032_),
    .Y(_09034_));
 sky130_as_sc_hs__and2_2 _39773_ (.A(_09033_),
    .B(_09034_),
    .Y(_09035_));
 sky130_as_sc_hs__or2_2 _39775_ (.A(_09022_),
    .B(_09035_),
    .Y(_09037_));
 sky130_as_sc_hs__and2_2 _39776_ (.A(_09036_),
    .B(_09037_),
    .Y(_09038_));
 sky130_as_sc_hs__or2_2 _39778_ (.A(_09013_),
    .B(_09038_),
    .Y(_09040_));
 sky130_as_sc_hs__and2_2 _39779_ (.A(_09039_),
    .B(_09040_),
    .Y(_09041_));
 sky130_as_sc_hs__or2_2 _39781_ (.A(_09012_),
    .B(_09041_),
    .Y(_09043_));
 sky130_as_sc_hs__and2_2 _39782_ (.A(_09042_),
    .B(_09043_),
    .Y(_09044_));
 sky130_as_sc_hs__and2_2 _39785_ (.A(net465),
    .B(net84),
    .Y(_09047_));
 sky130_as_sc_hs__and2_2 _39786_ (.A(net463),
    .B(net432),
    .Y(_09048_));
 sky130_as_sc_hs__or2_2 _39787_ (.A(_09047_),
    .B(_09048_),
    .Y(_09049_));
 sky130_as_sc_hs__and2_2 _39789_ (.A(_09049_),
    .B(_09050_),
    .Y(_09051_));
 sky130_as_sc_hs__and2_2 _39790_ (.A(net460),
    .B(net430),
    .Y(_09052_));
 sky130_as_sc_hs__or2_2 _39792_ (.A(_09051_),
    .B(_09052_),
    .Y(_09054_));
 sky130_as_sc_hs__and2_2 _39793_ (.A(_09053_),
    .B(_09054_),
    .Y(_09055_));
 sky130_as_sc_hs__or2_2 _39795_ (.A(_09046_),
    .B(_09055_),
    .Y(_09057_));
 sky130_as_sc_hs__and2_2 _39796_ (.A(_09056_),
    .B(_09057_),
    .Y(_09058_));
 sky130_as_sc_hs__or2_2 _39798_ (.A(_09045_),
    .B(_09058_),
    .Y(_09060_));
 sky130_as_sc_hs__and2_2 _39799_ (.A(_09059_),
    .B(_09060_),
    .Y(_09061_));
 sky130_as_sc_hs__nand3_2 _39801_ (.A(_24740_),
    .B(_24741_),
    .C(_25035_),
    .Y(_09063_));
 sky130_as_sc_hs__or2_2 _39803_ (.A(_09062_),
    .B(_09063_),
    .Y(_09065_));
 sky130_as_sc_hs__and2_2 _39804_ (.A(_09064_),
    .B(_09065_),
    .Y(_09066_));
 sky130_as_sc_hs__and2_2 _39805_ (.A(net481),
    .B(_24479_),
    .Y(_09067_));
 sky130_as_sc_hs__or2_2 _39807_ (.A(_09066_),
    .B(_09067_),
    .Y(_09069_));
 sky130_as_sc_hs__and2_2 _39808_ (.A(_09068_),
    .B(_09069_),
    .Y(_09070_));
 sky130_as_sc_hs__or2_2 _39811_ (.A(_09070_),
    .B(_09071_),
    .Y(_09073_));
 sky130_as_sc_hs__and2_2 _39812_ (.A(_09072_),
    .B(_09073_),
    .Y(_09074_));
 sky130_as_sc_hs__and2_2 _39813_ (.A(net473),
    .B(net466),
    .Y(_09075_));
 sky130_as_sc_hs__and2_2 _39814_ (.A(net479),
    .B(net468),
    .Y(_09076_));
 sky130_as_sc_hs__or2_2 _39815_ (.A(_09075_),
    .B(_09076_),
    .Y(_09077_));
 sky130_as_sc_hs__and2_2 _39817_ (.A(_09077_),
    .B(_09078_),
    .Y(_09079_));
 sky130_as_sc_hs__and2_2 _39818_ (.A(net475),
    .B(net470),
    .Y(_09080_));
 sky130_as_sc_hs__or2_2 _39820_ (.A(_09079_),
    .B(_09080_),
    .Y(_09082_));
 sky130_as_sc_hs__and2_2 _39821_ (.A(_09081_),
    .B(_09082_),
    .Y(_09083_));
 sky130_as_sc_hs__or2_2 _39823_ (.A(_09074_),
    .B(_09083_),
    .Y(_09085_));
 sky130_as_sc_hs__and2_2 _39824_ (.A(_09084_),
    .B(_09085_),
    .Y(_09086_));
 sky130_as_sc_hs__or2_2 _39827_ (.A(_09086_),
    .B(_09087_),
    .Y(_09089_));
 sky130_as_sc_hs__and2_2 _39828_ (.A(_09088_),
    .B(_09089_),
    .Y(_09090_));
 sky130_as_sc_hs__or2_2 _39830_ (.A(_09061_),
    .B(_09090_),
    .Y(_09092_));
 sky130_as_sc_hs__and2_2 _39831_ (.A(_09091_),
    .B(_09092_),
    .Y(_09093_));
 sky130_as_sc_hs__or2_2 _39834_ (.A(_09093_),
    .B(_09094_),
    .Y(_09096_));
 sky130_as_sc_hs__and2_2 _39835_ (.A(_09095_),
    .B(_09096_),
    .Y(_09097_));
 sky130_as_sc_hs__or2_2 _39837_ (.A(_09044_),
    .B(_09097_),
    .Y(_09099_));
 sky130_as_sc_hs__and2_2 _39838_ (.A(_09098_),
    .B(_09099_),
    .Y(_09100_));
 sky130_as_sc_hs__or2_2 _39841_ (.A(_09100_),
    .B(_09101_),
    .Y(_09103_));
 sky130_as_sc_hs__and2_2 _39842_ (.A(_09102_),
    .B(_09103_),
    .Y(_09104_));
 sky130_as_sc_hs__or2_2 _39844_ (.A(_09011_),
    .B(_09104_),
    .Y(_09106_));
 sky130_as_sc_hs__and2_2 _39845_ (.A(_09105_),
    .B(_09106_),
    .Y(_09107_));
 sky130_as_sc_hs__or2_2 _39848_ (.A(_09107_),
    .B(_09108_),
    .Y(_09110_));
 sky130_as_sc_hs__and2_2 _39849_ (.A(_09109_),
    .B(_09110_),
    .Y(_09111_));
 sky130_as_sc_hs__or2_2 _39851_ (.A(_08979_),
    .B(_09111_),
    .Y(_09113_));
 sky130_as_sc_hs__and2_2 _39852_ (.A(_09112_),
    .B(_09113_),
    .Y(_09114_));
 sky130_as_sc_hs__or2_2 _39855_ (.A(_09114_),
    .B(_09115_),
    .Y(_09117_));
 sky130_as_sc_hs__and2_2 _39856_ (.A(_09116_),
    .B(_09117_),
    .Y(_09118_));
 sky130_as_sc_hs__or2_2 _39858_ (.A(_08953_),
    .B(_09118_),
    .Y(_09120_));
 sky130_as_sc_hs__and2_2 _39859_ (.A(_09119_),
    .B(_09120_),
    .Y(_09121_));
 sky130_as_sc_hs__or2_2 _39862_ (.A(_09121_),
    .B(_09122_),
    .Y(_09124_));
 sky130_as_sc_hs__and2_2 _39863_ (.A(_09123_),
    .B(_09124_),
    .Y(_09125_));
 sky130_as_sc_hs__and2_2 _39864_ (.A(_08716_),
    .B(_08717_),
    .Y(_09126_));
 sky130_as_sc_hs__or2_2 _39866_ (.A(_09125_),
    .B(_09126_),
    .Y(_09128_));
 sky130_as_sc_hs__and2_2 _39867_ (.A(_09127_),
    .B(_09128_),
    .Y(_09129_));
 sky130_as_sc_hs__or2_2 _39870_ (.A(_09129_),
    .B(_09130_),
    .Y(_09132_));
 sky130_as_sc_hs__and2_2 _39871_ (.A(_09131_),
    .B(_09132_),
    .Y(_09133_));
 sky130_as_sc_hs__and2_2 _39874_ (.A(_08620_),
    .B(_08885_),
    .Y(_09136_));
 sky130_as_sc_hs__or2_2 _39878_ (.A(_09133_),
    .B(_09138_),
    .Y(_09140_));
 sky130_as_sc_hs__and2_2 _39882_ (.A(_08637_),
    .B(_09143_),
    .Y(_09144_));
 sky130_as_sc_hs__or2_2 _39884_ (.A(_09141_),
    .B(_09144_),
    .Y(_09146_));
 sky130_as_sc_hs__nand3_2 _39885_ (.A(net142),
    .B(_09145_),
    .C(_09146_),
    .Y(_09147_));
 sky130_as_sc_hs__or2_2 _39886_ (.A(_05410_),
    .B(_05505_),
    .Y(_09148_));
 sky130_as_sc_hs__or2_2 _39887_ (.A(_05388_),
    .B(_09148_),
    .Y(_09149_));
 sky130_as_sc_hs__nand3_2 _39889_ (.A(net139),
    .B(_09149_),
    .C(_09150_),
    .Y(_09151_));
 sky130_as_sc_hs__and2_2 _39891_ (.A(_05735_),
    .B(_09152_),
    .Y(_09153_));
 sky130_as_sc_hs__or2_2 _39892_ (.A(_05726_),
    .B(_09153_),
    .Y(_09154_));
 sky130_as_sc_hs__or2_2 _39896_ (.A(_05726_),
    .B(_05869_),
    .Y(_09158_));
 sky130_as_sc_hs__nand3_2 _39899_ (.A(net119),
    .B(_09157_),
    .C(_09160_),
    .Y(_09161_));
 sky130_as_sc_hs__and2_2 _39902_ (.A(_05926_),
    .B(_09163_),
    .Y(_09164_));
 sky130_as_sc_hs__or2_2 _39903_ (.A(_05935_),
    .B(_06861_),
    .Y(_09165_));
 sky130_as_sc_hs__or2_2 _39904_ (.A(_05936_),
    .B(_06836_),
    .Y(_09166_));
 sky130_as_sc_hs__nand3_2 _39905_ (.A(_05929_),
    .B(_09165_),
    .C(_09166_),
    .Y(_09167_));
 sky130_as_sc_hs__or2_2 _39906_ (.A(_05929_),
    .B(_07818_),
    .Y(_09168_));
 sky130_as_sc_hs__and2_2 _39907_ (.A(_09167_),
    .B(_09168_),
    .Y(_09169_));
 sky130_as_sc_hs__or2_2 _39910_ (.A(_05724_),
    .B(_06161_),
    .Y(_09172_));
 sky130_as_sc_hs__nand3_2 _39911_ (.A(_06158_),
    .B(_09171_),
    .C(_09172_),
    .Y(_09173_));
 sky130_as_sc_hs__and2_2 _39912_ (.A(_05725_),
    .B(_09173_),
    .Y(_09174_));
 sky130_as_sc_hs__or2_2 _39913_ (.A(\tholin_riscv.div_res[9] ),
    .B(_08917_),
    .Y(_09175_));
 sky130_as_sc_hs__and2_2 _39914_ (.A(net415),
    .B(_09175_),
    .Y(_09176_));
 sky130_as_sc_hs__or2_2 _39915_ (.A(\tholin_riscv.div_res[10] ),
    .B(_09176_),
    .Y(_09177_));
 sky130_as_sc_hs__nand3_2 _39917_ (.A(net111),
    .B(_09177_),
    .C(_09178_),
    .Y(_09179_));
 sky130_as_sc_hs__or2_2 _39918_ (.A(\tholin_riscv.div_shifter[41] ),
    .B(_08925_),
    .Y(_09180_));
 sky130_as_sc_hs__and2_2 _39919_ (.A(_21655_),
    .B(_09180_),
    .Y(_09181_));
 sky130_as_sc_hs__or2_2 _39921_ (.A(\tholin_riscv.div_shifter[42] ),
    .B(_09181_),
    .Y(_09183_));
 sky130_as_sc_hs__nand3_2 _39922_ (.A(net108),
    .B(_09182_),
    .C(_09183_),
    .Y(_09184_));
 sky130_as_sc_hs__and2_2 _39925_ (.A(_09185_),
    .B(_09186_),
    .Y(_09187_));
 sky130_as_sc_hs__nand3_2 _39926_ (.A(net412),
    .B(_09184_),
    .C(_09187_),
    .Y(_09188_));
 sky130_as_sc_hs__nor2_2 _39927_ (.A(_09174_),
    .B(_09188_),
    .Y(_09189_));
 sky130_as_sc_hs__nand3_2 _39928_ (.A(_09170_),
    .B(_09179_),
    .C(_09189_),
    .Y(_09190_));
 sky130_as_sc_hs__nor2_2 _39929_ (.A(_09164_),
    .B(_09190_),
    .Y(_09191_));
 sky130_as_sc_hs__and2_2 _39930_ (.A(_09161_),
    .B(_09191_),
    .Y(_09192_));
 sky130_as_sc_hs__nand3_2 _39931_ (.A(_09147_),
    .B(_09151_),
    .C(_09192_),
    .Y(_09193_));
 sky130_as_sc_hs__and2_2 _39932_ (.A(\tholin_riscv.PC[10] ),
    .B(_08941_),
    .Y(_09194_));
 sky130_as_sc_hs__nor2_2 _39933_ (.A(\tholin_riscv.PC[10] ),
    .B(_08941_),
    .Y(_09195_));
 sky130_as_sc_hs__nor2_2 _39934_ (.A(_09194_),
    .B(_09195_),
    .Y(_09196_));
 sky130_as_sc_hs__inv_2 _39935_ (.Y(_09197_),
    .A(_09196_));
 sky130_as_sc_hs__nand3_2 _39938_ (.A(_21569_),
    .B(_09198_),
    .C(_09199_),
    .Y(_09200_));
 sky130_as_sc_hs__nand3_2 _39939_ (.A(_21546_),
    .B(_09193_),
    .C(_09200_),
    .Y(_09201_));
 sky130_as_sc_hs__or2_2 _39944_ (.A(_19843_),
    .B(_08428_),
    .Y(_09205_));
 sky130_as_sc_hs__nor2_2 _39951_ (.A(_08957_),
    .B(_09211_),
    .Y(_09212_));
 sky130_as_sc_hs__and2_2 _39952_ (.A(_08957_),
    .B(_09211_),
    .Y(_09213_));
 sky130_as_sc_hs__nor2_2 _39953_ (.A(_09212_),
    .B(_09213_),
    .Y(_09214_));
 sky130_as_sc_hs__and2_2 _39954_ (.A(net446),
    .B(net128),
    .Y(_09215_));
 sky130_as_sc_hs__or2_2 _39956_ (.A(_08984_),
    .B(_09215_),
    .Y(_09217_));
 sky130_as_sc_hs__or2_2 _39958_ (.A(_08965_),
    .B(_09218_),
    .Y(_09219_));
 sky130_as_sc_hs__and2_2 _39960_ (.A(_09219_),
    .B(_09220_),
    .Y(_09221_));
 sky130_as_sc_hs__or2_2 _39962_ (.A(_09214_),
    .B(_09221_),
    .Y(_09223_));
 sky130_as_sc_hs__and2_2 _39963_ (.A(_09222_),
    .B(_09223_),
    .Y(_09224_));
 sky130_as_sc_hs__or2_2 _39965_ (.A(_09210_),
    .B(_09224_),
    .Y(_09226_));
 sky130_as_sc_hs__and2_2 _39966_ (.A(_09225_),
    .B(_09226_),
    .Y(_09227_));
 sky130_as_sc_hs__or2_2 _39968_ (.A(_09209_),
    .B(_09227_),
    .Y(_09229_));
 sky130_as_sc_hs__and2_2 _39969_ (.A(_09228_),
    .B(_09229_),
    .Y(_09230_));
 sky130_as_sc_hs__and2_2 _39972_ (.A(net440),
    .B(net438),
    .Y(_09233_));
 sky130_as_sc_hs__and2_2 _39973_ (.A(net472),
    .B(net436),
    .Y(_09234_));
 sky130_as_sc_hs__and2_2 _39974_ (.A(_09233_),
    .B(_09234_),
    .Y(_09235_));
 sky130_as_sc_hs__or2_2 _39975_ (.A(_09233_),
    .B(_09234_),
    .Y(_09236_));
 sky130_as_sc_hs__nor2b_2 _39976_ (.A(_09235_),
    .Y(_09237_),
    .B(_09236_));
 sky130_as_sc_hs__and2_2 _39977_ (.A(net480),
    .B(net435),
    .Y(_09238_));
 sky130_as_sc_hs__or2_2 _39980_ (.A(_09238_),
    .B(_09239_),
    .Y(_09241_));
 sky130_as_sc_hs__or2_2 _39982_ (.A(_08990_),
    .B(_09242_),
    .Y(_09243_));
 sky130_as_sc_hs__and2_2 _39984_ (.A(_09243_),
    .B(_09244_),
    .Y(_09245_));
 sky130_as_sc_hs__or2_2 _39987_ (.A(_09245_),
    .B(_09246_),
    .Y(_09248_));
 sky130_as_sc_hs__and2_2 _39988_ (.A(_09247_),
    .B(_09248_),
    .Y(_09249_));
 sky130_as_sc_hs__or2_2 _39990_ (.A(_09237_),
    .B(_09249_),
    .Y(_09251_));
 sky130_as_sc_hs__and2_2 _39991_ (.A(_09250_),
    .B(_09251_),
    .Y(_09252_));
 sky130_as_sc_hs__or2_2 _39993_ (.A(_09232_),
    .B(_09252_),
    .Y(_09254_));
 sky130_as_sc_hs__and2_2 _39994_ (.A(_09253_),
    .B(_09254_),
    .Y(_09255_));
 sky130_as_sc_hs__or2_2 _39996_ (.A(_09231_),
    .B(_09255_),
    .Y(_09257_));
 sky130_as_sc_hs__and2_2 _39997_ (.A(_09256_),
    .B(_09257_),
    .Y(_09258_));
 sky130_as_sc_hs__and2_2 _40000_ (.A(net442),
    .B(net426),
    .Y(_09261_));
 sky130_as_sc_hs__and2_2 _40001_ (.A(net449),
    .B(net420),
    .Y(_09262_));
 sky130_as_sc_hs__or2_2 _40002_ (.A(_09261_),
    .B(_09262_),
    .Y(_09263_));
 sky130_as_sc_hs__and2_2 _40004_ (.A(_09263_),
    .B(_09264_),
    .Y(_09265_));
 sky130_as_sc_hs__and2_2 _40005_ (.A(net451),
    .B(net74),
    .Y(_09266_));
 sky130_as_sc_hs__or2_2 _40007_ (.A(_09265_),
    .B(_09266_),
    .Y(_09268_));
 sky130_as_sc_hs__and2_2 _40008_ (.A(_09267_),
    .B(_09268_),
    .Y(_09269_));
 sky130_as_sc_hs__or2_2 _40012_ (.A(_09270_),
    .B(_09271_),
    .Y(_09273_));
 sky130_as_sc_hs__and2_2 _40013_ (.A(_09272_),
    .B(_09273_),
    .Y(_09274_));
 sky130_as_sc_hs__and2_2 _40014_ (.A(net88),
    .B(net424),
    .Y(_09275_));
 sky130_as_sc_hs__or2_2 _40016_ (.A(_09274_),
    .B(_09275_),
    .Y(_09277_));
 sky130_as_sc_hs__and2_2 _40017_ (.A(_09276_),
    .B(_09277_),
    .Y(_09278_));
 sky130_as_sc_hs__or2_2 _40020_ (.A(_09278_),
    .B(_09279_),
    .Y(_09281_));
 sky130_as_sc_hs__and2_2 _40021_ (.A(_09280_),
    .B(_09281_),
    .Y(_09282_));
 sky130_as_sc_hs__or2_2 _40023_ (.A(_09269_),
    .B(_09282_),
    .Y(_09284_));
 sky130_as_sc_hs__and2_2 _40024_ (.A(_09283_),
    .B(_09284_),
    .Y(_09285_));
 sky130_as_sc_hs__or2_2 _40026_ (.A(_09260_),
    .B(_09285_),
    .Y(_09287_));
 sky130_as_sc_hs__and2_2 _40027_ (.A(_09286_),
    .B(_09287_),
    .Y(_09288_));
 sky130_as_sc_hs__or2_2 _40029_ (.A(_09259_),
    .B(_09288_),
    .Y(_09290_));
 sky130_as_sc_hs__and2_2 _40030_ (.A(_09289_),
    .B(_09290_),
    .Y(_09291_));
 sky130_as_sc_hs__or2_2 _40034_ (.A(_09292_),
    .B(_09293_),
    .Y(_09295_));
 sky130_as_sc_hs__and2_2 _40035_ (.A(_09294_),
    .B(_09295_),
    .Y(_09296_));
 sky130_as_sc_hs__and2_2 _40036_ (.A(net476),
    .B(net457),
    .Y(_09297_));
 sky130_as_sc_hs__or2_2 _40038_ (.A(_09296_),
    .B(_09297_),
    .Y(_09299_));
 sky130_as_sc_hs__and2_2 _40039_ (.A(_09298_),
    .B(_09299_),
    .Y(_09300_));
 sky130_as_sc_hs__or2_2 _40042_ (.A(_09300_),
    .B(_09301_),
    .Y(_09303_));
 sky130_as_sc_hs__and2_2 _40043_ (.A(_09302_),
    .B(_09303_),
    .Y(_09304_));
 sky130_as_sc_hs__and2_2 _40044_ (.A(net478),
    .B(net466),
    .Y(_09305_));
 sky130_as_sc_hs__and2_2 _40045_ (.A(net474),
    .B(net468),
    .Y(_09306_));
 sky130_as_sc_hs__or2_2 _40046_ (.A(_09305_),
    .B(_09306_),
    .Y(_09307_));
 sky130_as_sc_hs__and2_2 _40048_ (.A(_09307_),
    .B(_09308_),
    .Y(_09309_));
 sky130_as_sc_hs__and2_2 _40049_ (.A(net471),
    .B(net83),
    .Y(_09310_));
 sky130_as_sc_hs__or2_2 _40051_ (.A(_09309_),
    .B(_09310_),
    .Y(_09312_));
 sky130_as_sc_hs__and2_2 _40052_ (.A(_09311_),
    .B(_09312_),
    .Y(_09313_));
 sky130_as_sc_hs__or2_2 _40054_ (.A(_09304_),
    .B(_09313_),
    .Y(_09315_));
 sky130_as_sc_hs__and2_2 _40055_ (.A(_09314_),
    .B(_09315_),
    .Y(_09316_));
 sky130_as_sc_hs__or2_2 _40058_ (.A(_09316_),
    .B(_09317_),
    .Y(_09319_));
 sky130_as_sc_hs__and2_2 _40059_ (.A(_09318_),
    .B(_09319_),
    .Y(_09320_));
 sky130_as_sc_hs__and2_2 _40062_ (.A(net465),
    .B(net431),
    .Y(_09323_));
 sky130_as_sc_hs__and2_2 _40063_ (.A(net463),
    .B(net429),
    .Y(_09324_));
 sky130_as_sc_hs__or2_2 _40064_ (.A(_09323_),
    .B(_09324_),
    .Y(_09325_));
 sky130_as_sc_hs__and2_2 _40066_ (.A(_09325_),
    .B(_09326_),
    .Y(_09327_));
 sky130_as_sc_hs__and2_2 _40067_ (.A(net460),
    .B(net427),
    .Y(_09328_));
 sky130_as_sc_hs__or2_2 _40069_ (.A(_09327_),
    .B(_09328_),
    .Y(_09330_));
 sky130_as_sc_hs__and2_2 _40070_ (.A(_09329_),
    .B(_09330_),
    .Y(_09331_));
 sky130_as_sc_hs__or2_2 _40072_ (.A(_09322_),
    .B(_09331_),
    .Y(_09333_));
 sky130_as_sc_hs__and2_2 _40073_ (.A(_09332_),
    .B(_09333_),
    .Y(_09334_));
 sky130_as_sc_hs__or2_2 _40075_ (.A(_09321_),
    .B(_09334_),
    .Y(_09336_));
 sky130_as_sc_hs__and2_2 _40076_ (.A(_09335_),
    .B(_09336_),
    .Y(_09337_));
 sky130_as_sc_hs__or2_2 _40078_ (.A(_09320_),
    .B(_09337_),
    .Y(_09339_));
 sky130_as_sc_hs__and2_2 _40079_ (.A(_09338_),
    .B(_09339_),
    .Y(_09340_));
 sky130_as_sc_hs__or2_2 _40082_ (.A(_09340_),
    .B(_09341_),
    .Y(_09343_));
 sky130_as_sc_hs__and2_2 _40083_ (.A(_09342_),
    .B(_09343_),
    .Y(_09344_));
 sky130_as_sc_hs__or2_2 _40085_ (.A(_09291_),
    .B(_09344_),
    .Y(_09346_));
 sky130_as_sc_hs__and2_2 _40086_ (.A(_09345_),
    .B(_09346_),
    .Y(_09347_));
 sky130_as_sc_hs__or2_2 _40089_ (.A(_09347_),
    .B(_09348_),
    .Y(_09350_));
 sky130_as_sc_hs__and2_2 _40090_ (.A(_09349_),
    .B(_09350_),
    .Y(_09351_));
 sky130_as_sc_hs__or2_2 _40092_ (.A(_09258_),
    .B(_09351_),
    .Y(_09353_));
 sky130_as_sc_hs__and2_2 _40093_ (.A(_09352_),
    .B(_09353_),
    .Y(_09354_));
 sky130_as_sc_hs__or2_2 _40096_ (.A(_09354_),
    .B(_09355_),
    .Y(_09357_));
 sky130_as_sc_hs__and2_2 _40097_ (.A(_09356_),
    .B(_09357_),
    .Y(_09358_));
 sky130_as_sc_hs__or2_2 _40099_ (.A(_09230_),
    .B(_09358_),
    .Y(_09360_));
 sky130_as_sc_hs__and2_2 _40100_ (.A(_09359_),
    .B(_09360_),
    .Y(_09361_));
 sky130_as_sc_hs__or2_2 _40103_ (.A(_09361_),
    .B(_09362_),
    .Y(_09364_));
 sky130_as_sc_hs__and2_2 _40104_ (.A(_09363_),
    .B(_09364_),
    .Y(_09365_));
 sky130_as_sc_hs__or2_2 _40106_ (.A(_09208_),
    .B(_09365_),
    .Y(_09367_));
 sky130_as_sc_hs__and2_2 _40107_ (.A(_09366_),
    .B(_09367_),
    .Y(_09368_));
 sky130_as_sc_hs__or2_2 _40110_ (.A(_09368_),
    .B(_09369_),
    .Y(_09371_));
 sky130_as_sc_hs__or2_2 _40112_ (.A(_08961_),
    .B(_09372_),
    .Y(_09373_));
 sky130_as_sc_hs__and2_2 _40114_ (.A(_09373_),
    .B(_09374_),
    .Y(_09375_));
 sky130_as_sc_hs__or2_2 _40116_ (.A(_09207_),
    .B(_09375_),
    .Y(_09377_));
 sky130_as_sc_hs__and2_2 _40117_ (.A(_09376_),
    .B(_09377_),
    .Y(_09378_));
 sky130_as_sc_hs__and2_2 _40118_ (.A(_09131_),
    .B(_09139_),
    .Y(_09379_));
 sky130_as_sc_hs__or2_2 _40120_ (.A(_09378_),
    .B(_09379_),
    .Y(_09381_));
 sky130_as_sc_hs__and2_2 _40121_ (.A(_09380_),
    .B(_09381_),
    .Y(_09382_));
 sky130_as_sc_hs__nor2b_2 _40122_ (.A(_09142_),
    .Y(_09383_),
    .B(_09141_));
 sky130_as_sc_hs__or2_2 _40123_ (.A(_05505_),
    .B(_09383_),
    .Y(_09384_));
 sky130_as_sc_hs__and2_2 _40124_ (.A(_08637_),
    .B(_09384_),
    .Y(_09385_));
 sky130_as_sc_hs__or2_2 _40126_ (.A(_09382_),
    .B(_09385_),
    .Y(_09387_));
 sky130_as_sc_hs__nand3_2 _40127_ (.A(net142),
    .B(_09386_),
    .C(_09387_),
    .Y(_09388_));
 sky130_as_sc_hs__or2_2 _40130_ (.A(_05416_),
    .B(_09389_),
    .Y(_09391_));
 sky130_as_sc_hs__nand3_2 _40131_ (.A(net138),
    .B(_09390_),
    .C(_09391_),
    .Y(_09392_));
 sky130_as_sc_hs__and2_2 _40132_ (.A(_05724_),
    .B(_09154_),
    .Y(_09393_));
 sky130_as_sc_hs__or2_2 _40133_ (.A(_05715_),
    .B(_09393_),
    .Y(_09394_));
 sky130_as_sc_hs__or2_2 _40137_ (.A(_05715_),
    .B(_05871_),
    .Y(_09398_));
 sky130_as_sc_hs__nand3_2 _40140_ (.A(_06523_),
    .B(_09397_),
    .C(_09400_),
    .Y(_09401_));
 sky130_as_sc_hs__and2_2 _40143_ (.A(_05926_),
    .B(_09403_),
    .Y(_09404_));
 sky130_as_sc_hs__or2_2 _40144_ (.A(_05935_),
    .B(_07227_),
    .Y(_09405_));
 sky130_as_sc_hs__or2_2 _40145_ (.A(_05936_),
    .B(_07202_),
    .Y(_09406_));
 sky130_as_sc_hs__nand3_2 _40146_ (.A(_05929_),
    .B(_09405_),
    .C(_09406_),
    .Y(_09407_));
 sky130_as_sc_hs__or2_2 _40147_ (.A(_05929_),
    .B(_07526_),
    .Y(_09408_));
 sky130_as_sc_hs__and2_2 _40148_ (.A(_09407_),
    .B(_09408_),
    .Y(_09409_));
 sky130_as_sc_hs__or2_2 _40151_ (.A(_05713_),
    .B(_06161_),
    .Y(_09412_));
 sky130_as_sc_hs__nand3_2 _40152_ (.A(_06158_),
    .B(_09411_),
    .C(_09412_),
    .Y(_09413_));
 sky130_as_sc_hs__and2_2 _40153_ (.A(_05714_),
    .B(_09413_),
    .Y(_09414_));
 sky130_as_sc_hs__or2_2 _40154_ (.A(\tholin_riscv.div_res[10] ),
    .B(_09175_),
    .Y(_09415_));
 sky130_as_sc_hs__and2_2 _40155_ (.A(net415),
    .B(_09415_),
    .Y(_09416_));
 sky130_as_sc_hs__or2_2 _40156_ (.A(\tholin_riscv.div_res[11] ),
    .B(_09416_),
    .Y(_09417_));
 sky130_as_sc_hs__nand3_2 _40158_ (.A(net111),
    .B(_09417_),
    .C(_09418_),
    .Y(_09419_));
 sky130_as_sc_hs__or2_2 _40159_ (.A(\tholin_riscv.div_shifter[42] ),
    .B(_09180_),
    .Y(_09420_));
 sky130_as_sc_hs__and2_2 _40160_ (.A(_21655_),
    .B(_09420_),
    .Y(_09421_));
 sky130_as_sc_hs__or2_2 _40162_ (.A(\tholin_riscv.div_shifter[43] ),
    .B(_09421_),
    .Y(_09423_));
 sky130_as_sc_hs__nand3_2 _40163_ (.A(net108),
    .B(_09422_),
    .C(_09423_),
    .Y(_09424_));
 sky130_as_sc_hs__and2_2 _40166_ (.A(_09425_),
    .B(_09426_),
    .Y(_09427_));
 sky130_as_sc_hs__nand3_2 _40167_ (.A(net412),
    .B(_09424_),
    .C(_09427_),
    .Y(_09428_));
 sky130_as_sc_hs__nor2_2 _40168_ (.A(_09414_),
    .B(_09428_),
    .Y(_09429_));
 sky130_as_sc_hs__nand3_2 _40169_ (.A(_09410_),
    .B(_09419_),
    .C(_09429_),
    .Y(_09430_));
 sky130_as_sc_hs__nor2_2 _40170_ (.A(_09404_),
    .B(_09430_),
    .Y(_09431_));
 sky130_as_sc_hs__and2_2 _40171_ (.A(_09401_),
    .B(_09431_),
    .Y(_09432_));
 sky130_as_sc_hs__nand3_2 _40172_ (.A(_09388_),
    .B(_09392_),
    .C(_09432_),
    .Y(_09433_));
 sky130_as_sc_hs__and2_2 _40173_ (.A(\tholin_riscv.PC[11] ),
    .B(_09194_),
    .Y(_09434_));
 sky130_as_sc_hs__nor2_2 _40174_ (.A(\tholin_riscv.PC[11] ),
    .B(_09194_),
    .Y(_09435_));
 sky130_as_sc_hs__nor2_2 _40175_ (.A(_09434_),
    .B(_09435_),
    .Y(_09436_));
 sky130_as_sc_hs__inv_2 _40176_ (.Y(_09437_),
    .A(_09436_));
 sky130_as_sc_hs__nand3_2 _40179_ (.A(_21569_),
    .B(_09438_),
    .C(_09439_),
    .Y(_09440_));
 sky130_as_sc_hs__nand3_2 _40180_ (.A(_21546_),
    .B(_09433_),
    .C(_09440_),
    .Y(_09441_));
 sky130_as_sc_hs__or2_2 _40185_ (.A(_19851_),
    .B(_08428_),
    .Y(_09445_));
 sky130_as_sc_hs__and2_2 _40190_ (.A(net78),
    .B(net128),
    .Y(_09450_));
 sky130_as_sc_hs__or2_2 _40192_ (.A(_09235_),
    .B(_09450_),
    .Y(_09452_));
 sky130_as_sc_hs__or2_2 _40194_ (.A(_09216_),
    .B(_09453_),
    .Y(_09454_));
 sky130_as_sc_hs__and2_2 _40196_ (.A(_09454_),
    .B(_09455_),
    .Y(_09456_));
 sky130_as_sc_hs__and2_2 _40197_ (.A(net442),
    .B(net421),
    .Y(_09457_));
 sky130_as_sc_hs__or2_2 _40199_ (.A(_09456_),
    .B(_09457_),
    .Y(_09459_));
 sky130_as_sc_hs__and2_2 _40200_ (.A(_09458_),
    .B(_09459_),
    .Y(_09460_));
 sky130_as_sc_hs__or2_2 _40202_ (.A(_09449_),
    .B(_09460_),
    .Y(_09462_));
 sky130_as_sc_hs__and2_2 _40203_ (.A(_09461_),
    .B(_09462_),
    .Y(_09463_));
 sky130_as_sc_hs__or2_2 _40205_ (.A(_09448_),
    .B(_09463_),
    .Y(_09465_));
 sky130_as_sc_hs__and2_2 _40206_ (.A(_09464_),
    .B(_09465_),
    .Y(_09466_));
 sky130_as_sc_hs__and2_2 _40209_ (.A(net472),
    .B(net440),
    .Y(_09469_));
 sky130_as_sc_hs__and2_2 _40210_ (.A(net478),
    .B(net436),
    .Y(_09470_));
 sky130_as_sc_hs__or2_2 _40212_ (.A(_09469_),
    .B(_09470_),
    .Y(_09472_));
 sky130_as_sc_hs__and2_2 _40213_ (.A(_09471_),
    .B(_09472_),
    .Y(_09473_));
 sky130_as_sc_hs__and2_2 _40214_ (.A(net476),
    .B(net434),
    .Y(_09474_));
 sky130_as_sc_hs__or2_2 _40217_ (.A(_09474_),
    .B(_09475_),
    .Y(_09477_));
 sky130_as_sc_hs__and2_2 _40218_ (.A(_09476_),
    .B(_09477_),
    .Y(_09478_));
 sky130_as_sc_hs__or2_2 _40221_ (.A(_09478_),
    .B(_09479_),
    .Y(_09481_));
 sky130_as_sc_hs__and2_2 _40222_ (.A(_09480_),
    .B(_09481_),
    .Y(_09482_));
 sky130_as_sc_hs__or2_2 _40224_ (.A(_09473_),
    .B(_09482_),
    .Y(_09484_));
 sky130_as_sc_hs__and2_2 _40225_ (.A(_09483_),
    .B(_09484_),
    .Y(_09485_));
 sky130_as_sc_hs__or2_2 _40227_ (.A(_09468_),
    .B(_09485_),
    .Y(_09487_));
 sky130_as_sc_hs__and2_2 _40228_ (.A(_09486_),
    .B(_09487_),
    .Y(_09488_));
 sky130_as_sc_hs__or2_2 _40230_ (.A(_09467_),
    .B(_09488_),
    .Y(_09490_));
 sky130_as_sc_hs__and2_2 _40231_ (.A(_09489_),
    .B(_09490_),
    .Y(_09491_));
 sky130_as_sc_hs__and2_2 _40232_ (.A(net446),
    .B(net418),
    .Y(_09492_));
 sky130_as_sc_hs__and2_2 _40233_ (.A(net480),
    .B(net433),
    .Y(_09493_));
 sky130_as_sc_hs__or2_2 _40234_ (.A(_09492_),
    .B(_09493_),
    .Y(_09494_));
 sky130_as_sc_hs__and2_2 _40236_ (.A(_09494_),
    .B(_09495_),
    .Y(_09496_));
 sky130_as_sc_hs__and2_2 _40237_ (.A(net457),
    .B(net438),
    .Y(_09497_));
 sky130_as_sc_hs__or2_2 _40239_ (.A(_09496_),
    .B(_09497_),
    .Y(_09499_));
 sky130_as_sc_hs__and2_2 _40240_ (.A(_09498_),
    .B(_09499_),
    .Y(_09500_));
 sky130_as_sc_hs__or2_2 _40243_ (.A(_09500_),
    .B(_09501_),
    .Y(_09503_));
 sky130_as_sc_hs__and2_2 _40244_ (.A(_09502_),
    .B(_09503_),
    .Y(_09504_));
 sky130_as_sc_hs__and2_2 _40245_ (.A(net474),
    .B(net466),
    .Y(_09505_));
 sky130_as_sc_hs__and2_2 _40246_ (.A(net468),
    .B(net83),
    .Y(_09506_));
 sky130_as_sc_hs__or2_2 _40247_ (.A(_09505_),
    .B(_09506_),
    .Y(_09507_));
 sky130_as_sc_hs__and2_2 _40249_ (.A(_09507_),
    .B(_09508_),
    .Y(_09509_));
 sky130_as_sc_hs__and2_2 _40250_ (.A(net471),
    .B(net431),
    .Y(_09510_));
 sky130_as_sc_hs__or2_2 _40252_ (.A(_09509_),
    .B(_09510_),
    .Y(_09512_));
 sky130_as_sc_hs__and2_2 _40253_ (.A(_09511_),
    .B(_09512_),
    .Y(_09513_));
 sky130_as_sc_hs__or2_2 _40255_ (.A(_09504_),
    .B(_09513_),
    .Y(_09515_));
 sky130_as_sc_hs__and2_2 _40256_ (.A(_09514_),
    .B(_09515_),
    .Y(_09516_));
 sky130_as_sc_hs__or2_2 _40259_ (.A(_09516_),
    .B(_09517_),
    .Y(_09519_));
 sky130_as_sc_hs__and2_2 _40260_ (.A(_09518_),
    .B(_09519_),
    .Y(_09520_));
 sky130_as_sc_hs__and2_2 _40263_ (.A(net465),
    .B(net429),
    .Y(_09523_));
 sky130_as_sc_hs__and2_2 _40264_ (.A(net463),
    .B(net427),
    .Y(_09524_));
 sky130_as_sc_hs__or2_2 _40265_ (.A(_09523_),
    .B(_09524_),
    .Y(_09525_));
 sky130_as_sc_hs__and2_2 _40267_ (.A(_09525_),
    .B(_09526_),
    .Y(_09527_));
 sky130_as_sc_hs__and2_2 _40268_ (.A(net120),
    .B(net460),
    .Y(_09528_));
 sky130_as_sc_hs__or2_2 _40270_ (.A(_09527_),
    .B(_09528_),
    .Y(_09530_));
 sky130_as_sc_hs__and2_2 _40271_ (.A(_09529_),
    .B(_09530_),
    .Y(_09531_));
 sky130_as_sc_hs__or2_2 _40273_ (.A(_09522_),
    .B(_09531_),
    .Y(_09533_));
 sky130_as_sc_hs__and2_2 _40274_ (.A(_09532_),
    .B(_09533_),
    .Y(_09534_));
 sky130_as_sc_hs__or2_2 _40276_ (.A(_09521_),
    .B(_09534_),
    .Y(_09536_));
 sky130_as_sc_hs__and2_2 _40277_ (.A(_09535_),
    .B(_09536_),
    .Y(_09537_));
 sky130_as_sc_hs__or2_2 _40279_ (.A(_09520_),
    .B(_09537_),
    .Y(_09539_));
 sky130_as_sc_hs__and2_2 _40280_ (.A(_09538_),
    .B(_09539_),
    .Y(_09540_));
 sky130_as_sc_hs__or2_2 _40283_ (.A(_09540_),
    .B(_09541_),
    .Y(_09543_));
 sky130_as_sc_hs__and2_2 _40284_ (.A(_09542_),
    .B(_09543_),
    .Y(_09544_));
 sky130_as_sc_hs__and2_2 _40287_ (.A(_23674_),
    .B(net426),
    .Y(_09547_));
 sky130_as_sc_hs__and2_2 _40288_ (.A(net449),
    .B(net74),
    .Y(_09548_));
 sky130_as_sc_hs__or2_2 _40290_ (.A(_09547_),
    .B(_09548_),
    .Y(_09550_));
 sky130_as_sc_hs__and2_2 _40291_ (.A(_09549_),
    .B(_09550_),
    .Y(_09551_));
 sky130_as_sc_hs__and2_2 _40292_ (.A(net122),
    .B(_24527_),
    .Y(_09552_));
 sky130_as_sc_hs__and2_2 _40293_ (.A(net89),
    .B(net424),
    .Y(_09553_));
 sky130_as_sc_hs__or2_2 _40294_ (.A(_09552_),
    .B(_09553_),
    .Y(_09554_));
 sky130_as_sc_hs__and2_2 _40296_ (.A(_09554_),
    .B(_09555_),
    .Y(_09556_));
 sky130_as_sc_hs__and2_2 _40297_ (.A(net88),
    .B(net419),
    .Y(_09557_));
 sky130_as_sc_hs__or2_2 _40299_ (.A(_09556_),
    .B(_09557_),
    .Y(_09559_));
 sky130_as_sc_hs__and2_2 _40300_ (.A(_09558_),
    .B(_09559_),
    .Y(_09560_));
 sky130_as_sc_hs__or2_2 _40303_ (.A(_09560_),
    .B(_09561_),
    .Y(_09563_));
 sky130_as_sc_hs__and2_2 _40304_ (.A(_09562_),
    .B(_09563_),
    .Y(_09564_));
 sky130_as_sc_hs__or2_2 _40306_ (.A(_09551_),
    .B(_09564_),
    .Y(_09566_));
 sky130_as_sc_hs__and2_2 _40307_ (.A(_09565_),
    .B(_09566_),
    .Y(_09567_));
 sky130_as_sc_hs__or2_2 _40309_ (.A(_09546_),
    .B(_09567_),
    .Y(_09569_));
 sky130_as_sc_hs__and2_2 _40310_ (.A(_09568_),
    .B(_09569_),
    .Y(_09570_));
 sky130_as_sc_hs__or2_2 _40312_ (.A(_09545_),
    .B(_09570_),
    .Y(_09572_));
 sky130_as_sc_hs__and2_2 _40313_ (.A(_09571_),
    .B(_09572_),
    .Y(_09573_));
 sky130_as_sc_hs__or2_2 _40315_ (.A(_09544_),
    .B(_09573_),
    .Y(_09575_));
 sky130_as_sc_hs__and2_2 _40316_ (.A(_09574_),
    .B(_09575_),
    .Y(_09576_));
 sky130_as_sc_hs__or2_2 _40319_ (.A(_09576_),
    .B(_09577_),
    .Y(_09579_));
 sky130_as_sc_hs__and2_2 _40320_ (.A(_09578_),
    .B(_09579_),
    .Y(_09580_));
 sky130_as_sc_hs__or2_2 _40322_ (.A(_09491_),
    .B(_09580_),
    .Y(_09582_));
 sky130_as_sc_hs__and2_2 _40323_ (.A(_09581_),
    .B(_09582_),
    .Y(_09583_));
 sky130_as_sc_hs__or2_2 _40326_ (.A(_09583_),
    .B(_09584_),
    .Y(_09586_));
 sky130_as_sc_hs__and2_2 _40327_ (.A(_09585_),
    .B(_09586_),
    .Y(_09587_));
 sky130_as_sc_hs__or2_2 _40329_ (.A(_09466_),
    .B(_09587_),
    .Y(_09589_));
 sky130_as_sc_hs__and2_2 _40330_ (.A(_09588_),
    .B(_09589_),
    .Y(_09590_));
 sky130_as_sc_hs__or2_2 _40333_ (.A(_09590_),
    .B(_09591_),
    .Y(_09593_));
 sky130_as_sc_hs__and2_2 _40334_ (.A(_09592_),
    .B(_09593_),
    .Y(_09594_));
 sky130_as_sc_hs__or2_2 _40336_ (.A(_09447_),
    .B(_09594_),
    .Y(_09596_));
 sky130_as_sc_hs__and2_2 _40337_ (.A(_09595_),
    .B(_09596_),
    .Y(_09597_));
 sky130_as_sc_hs__or2_2 _40340_ (.A(_09597_),
    .B(_09598_),
    .Y(_09600_));
 sky130_as_sc_hs__and2_2 _40341_ (.A(_09599_),
    .B(_09600_),
    .Y(_09601_));
 sky130_as_sc_hs__or2_2 _40343_ (.A(_09212_),
    .B(_09601_),
    .Y(_09603_));
 sky130_as_sc_hs__and2_2 _40344_ (.A(_09602_),
    .B(_09603_),
    .Y(_09604_));
 sky130_as_sc_hs__or2_2 _40347_ (.A(_09604_),
    .B(_09605_),
    .Y(_09607_));
 sky130_as_sc_hs__and2_2 _40348_ (.A(_09606_),
    .B(_09607_),
    .Y(_09608_));
 sky130_as_sc_hs__and2_2 _40349_ (.A(_09133_),
    .B(_09378_),
    .Y(_09609_));
 sky130_as_sc_hs__nand2b_2 _40350_ (.B(_09609_),
    .Y(_09610_),
    .A(_09135_));
 sky130_as_sc_hs__nand2b_2 _40351_ (.B(_09377_),
    .Y(_09611_),
    .A(_09131_));
 sky130_as_sc_hs__and2_2 _40352_ (.A(_09376_),
    .B(_09611_),
    .Y(_09612_));
 sky130_as_sc_hs__and2_2 _40353_ (.A(_09610_),
    .B(_09612_),
    .Y(_09613_));
 sky130_as_sc_hs__and2_2 _40354_ (.A(_09136_),
    .B(_09609_),
    .Y(_09614_));
 sky130_as_sc_hs__or2_2 _40358_ (.A(_09608_),
    .B(_09616_),
    .Y(_09618_));
 sky130_as_sc_hs__and2_2 _40360_ (.A(_09382_),
    .B(_09383_),
    .Y(_09620_));
 sky130_as_sc_hs__or2_2 _40361_ (.A(_05505_),
    .B(_09620_),
    .Y(_09621_));
 sky130_as_sc_hs__and2_2 _40362_ (.A(_08637_),
    .B(_09621_),
    .Y(_09622_));
 sky130_as_sc_hs__or2_2 _40363_ (.A(_09619_),
    .B(_09622_),
    .Y(_09623_));
 sky130_as_sc_hs__nand3_2 _40365_ (.A(net142),
    .B(_09623_),
    .C(_09624_),
    .Y(_09625_));
 sky130_as_sc_hs__or2_2 _40366_ (.A(_05417_),
    .B(_05505_),
    .Y(_09626_));
 sky130_as_sc_hs__or2_2 _40367_ (.A(_05386_),
    .B(_09626_),
    .Y(_09627_));
 sky130_as_sc_hs__nand3_2 _40369_ (.A(net139),
    .B(_09627_),
    .C(_09628_),
    .Y(_09629_));
 sky130_as_sc_hs__and2_2 _40370_ (.A(_05713_),
    .B(_09394_),
    .Y(_09630_));
 sky130_as_sc_hs__or2_2 _40371_ (.A(_05706_),
    .B(_09630_),
    .Y(_09631_));
 sky130_as_sc_hs__or2_2 _40375_ (.A(_05706_),
    .B(_05873_),
    .Y(_09635_));
 sky130_as_sc_hs__nand3_2 _40378_ (.A(net119),
    .B(_09634_),
    .C(_09637_),
    .Y(_09638_));
 sky130_as_sc_hs__or2_2 _40379_ (.A(_05935_),
    .B(_07517_),
    .Y(_09639_));
 sky130_as_sc_hs__nand3_2 _40381_ (.A(_05929_),
    .B(_09639_),
    .C(_09640_),
    .Y(_09641_));
 sky130_as_sc_hs__or2_2 _40382_ (.A(_05929_),
    .B(_07237_),
    .Y(_09642_));
 sky130_as_sc_hs__and2_2 _40383_ (.A(_09641_),
    .B(_09642_),
    .Y(_09643_));
 sky130_as_sc_hs__and2_2 _40387_ (.A(net140),
    .B(_09646_),
    .Y(_09647_));
 sky130_as_sc_hs__or2_2 _40388_ (.A(\tholin_riscv.div_res[11] ),
    .B(_09415_),
    .Y(_09648_));
 sky130_as_sc_hs__and2_2 _40389_ (.A(net414),
    .B(_09648_),
    .Y(_09649_));
 sky130_as_sc_hs__or2_2 _40391_ (.A(\tholin_riscv.div_res[12] ),
    .B(_09649_),
    .Y(_09651_));
 sky130_as_sc_hs__nand3_2 _40392_ (.A(net111),
    .B(_09650_),
    .C(_09651_),
    .Y(_09652_));
 sky130_as_sc_hs__or2_2 _40396_ (.A(\tholin_riscv.div_shifter[43] ),
    .B(_09420_),
    .Y(_09656_));
 sky130_as_sc_hs__and2_2 _40397_ (.A(_21655_),
    .B(_09656_),
    .Y(_09657_));
 sky130_as_sc_hs__or2_2 _40399_ (.A(\tholin_riscv.div_shifter[44] ),
    .B(_09657_),
    .Y(_09659_));
 sky130_as_sc_hs__nand3_2 _40400_ (.A(net108),
    .B(_09658_),
    .C(_09659_),
    .Y(_09660_));
 sky130_as_sc_hs__nor2_2 _40401_ (.A(_05704_),
    .B(_06161_),
    .Y(_09661_));
 sky130_as_sc_hs__nand3_2 _40404_ (.A(net413),
    .B(_09662_),
    .C(_09663_),
    .Y(_09664_));
 sky130_as_sc_hs__nor2_2 _40405_ (.A(_09661_),
    .B(_09664_),
    .Y(_09665_));
 sky130_as_sc_hs__and2_2 _40406_ (.A(_09660_),
    .B(_09665_),
    .Y(_09666_));
 sky130_as_sc_hs__nand3_2 _40407_ (.A(_09652_),
    .B(_09655_),
    .C(_09666_),
    .Y(_09667_));
 sky130_as_sc_hs__nor2_2 _40408_ (.A(_09647_),
    .B(_09667_),
    .Y(_09668_));
 sky130_as_sc_hs__and2_2 _40409_ (.A(_09644_),
    .B(_09668_),
    .Y(_09669_));
 sky130_as_sc_hs__and2_2 _40410_ (.A(_09638_),
    .B(_09669_),
    .Y(_09670_));
 sky130_as_sc_hs__nand3_2 _40411_ (.A(_09625_),
    .B(_09629_),
    .C(_09670_),
    .Y(_09671_));
 sky130_as_sc_hs__and2_2 _40412_ (.A(\tholin_riscv.PC[12] ),
    .B(_09434_),
    .Y(_09672_));
 sky130_as_sc_hs__nor2_2 _40413_ (.A(\tholin_riscv.PC[12] ),
    .B(_09434_),
    .Y(_09673_));
 sky130_as_sc_hs__or2_2 _40414_ (.A(_09672_),
    .B(_09673_),
    .Y(_09674_));
 sky130_as_sc_hs__or2_2 _40415_ (.A(_21572_),
    .B(_09674_),
    .Y(_09675_));
 sky130_as_sc_hs__and2_2 _40416_ (.A(\tholin_riscv.PC[12] ),
    .B(_19472_),
    .Y(_09676_));
 sky130_as_sc_hs__or2_2 _40417_ (.A(\tholin_riscv.Jimm[12] ),
    .B(_09676_),
    .Y(_09677_));
 sky130_as_sc_hs__nand3_2 _40419_ (.A(_21572_),
    .B(_09677_),
    .C(_09678_),
    .Y(_09679_));
 sky130_as_sc_hs__nand3_2 _40420_ (.A(_21569_),
    .B(_09675_),
    .C(_09679_),
    .Y(_09680_));
 sky130_as_sc_hs__nand3_2 _40421_ (.A(_21546_),
    .B(_09671_),
    .C(_09680_),
    .Y(_09681_));
 sky130_as_sc_hs__or2_2 _40426_ (.A(_19859_),
    .B(_08428_),
    .Y(_09685_));
 sky130_as_sc_hs__or2_2 _40434_ (.A(_09471_),
    .B(_09692_),
    .Y(_09693_));
 sky130_as_sc_hs__or2_2 _40437_ (.A(_09451_),
    .B(_09695_),
    .Y(_09696_));
 sky130_as_sc_hs__and2_2 _40439_ (.A(_09696_),
    .B(_09697_),
    .Y(_09698_));
 sky130_as_sc_hs__and2_2 _40440_ (.A(_23674_),
    .B(net421),
    .Y(_09699_));
 sky130_as_sc_hs__or2_2 _40442_ (.A(_09698_),
    .B(_09699_),
    .Y(_09701_));
 sky130_as_sc_hs__and2_2 _40443_ (.A(_09700_),
    .B(_09701_),
    .Y(_09702_));
 sky130_as_sc_hs__or2_2 _40445_ (.A(_09691_),
    .B(_09702_),
    .Y(_09704_));
 sky130_as_sc_hs__and2_2 _40446_ (.A(_09703_),
    .B(_09704_),
    .Y(_09705_));
 sky130_as_sc_hs__or2_2 _40448_ (.A(_09690_),
    .B(_09705_),
    .Y(_09707_));
 sky130_as_sc_hs__and2_2 _40449_ (.A(_09706_),
    .B(_09707_),
    .Y(_09708_));
 sky130_as_sc_hs__and2_2 _40450_ (.A(net78),
    .B(_02550_),
    .Y(_09709_));
 sky130_as_sc_hs__and2_2 _40451_ (.A(net476),
    .B(net433),
    .Y(_09710_));
 sky130_as_sc_hs__or2_2 _40452_ (.A(_09709_),
    .B(_09710_),
    .Y(_09711_));
 sky130_as_sc_hs__and2_2 _40454_ (.A(_09711_),
    .B(_09712_),
    .Y(_09713_));
 sky130_as_sc_hs__and2_2 _40455_ (.A(net472),
    .B(net457),
    .Y(_09714_));
 sky130_as_sc_hs__or2_2 _40457_ (.A(_09713_),
    .B(_09714_),
    .Y(_09716_));
 sky130_as_sc_hs__and2_2 _40458_ (.A(_09715_),
    .B(_09716_),
    .Y(_09717_));
 sky130_as_sc_hs__or2_2 _40461_ (.A(_09717_),
    .B(_09718_),
    .Y(_09720_));
 sky130_as_sc_hs__and2_2 _40462_ (.A(_09719_),
    .B(_09720_),
    .Y(_09721_));
 sky130_as_sc_hs__or2_2 _40466_ (.A(_09722_),
    .B(_09723_),
    .Y(_09725_));
 sky130_as_sc_hs__and2_2 _40467_ (.A(_09724_),
    .B(_09725_),
    .Y(_09726_));
 sky130_as_sc_hs__and2_2 _40468_ (.A(net471),
    .B(net429),
    .Y(_09727_));
 sky130_as_sc_hs__or2_2 _40470_ (.A(_09726_),
    .B(_09727_),
    .Y(_09729_));
 sky130_as_sc_hs__and2_2 _40471_ (.A(_09728_),
    .B(_09729_),
    .Y(_09730_));
 sky130_as_sc_hs__or2_2 _40473_ (.A(_09721_),
    .B(_09730_),
    .Y(_09732_));
 sky130_as_sc_hs__and2_2 _40474_ (.A(_09731_),
    .B(_09732_),
    .Y(_09733_));
 sky130_as_sc_hs__or2_2 _40477_ (.A(_09733_),
    .B(_09734_),
    .Y(_09736_));
 sky130_as_sc_hs__and2_2 _40478_ (.A(_09735_),
    .B(_09736_),
    .Y(_09737_));
 sky130_as_sc_hs__and2_2 _40481_ (.A(net465),
    .B(net427),
    .Y(_09740_));
 sky130_as_sc_hs__and2_2 _40482_ (.A(net120),
    .B(net463),
    .Y(_09741_));
 sky130_as_sc_hs__or2_2 _40483_ (.A(_09740_),
    .B(_09741_),
    .Y(_09742_));
 sky130_as_sc_hs__and2_2 _40485_ (.A(_09742_),
    .B(_09743_),
    .Y(_09744_));
 sky130_as_sc_hs__and2_2 _40486_ (.A(net122),
    .B(net460),
    .Y(_09745_));
 sky130_as_sc_hs__or2_2 _40488_ (.A(_09744_),
    .B(_09745_),
    .Y(_09747_));
 sky130_as_sc_hs__and2_2 _40489_ (.A(_09746_),
    .B(_09747_),
    .Y(_09748_));
 sky130_as_sc_hs__or2_2 _40491_ (.A(_09739_),
    .B(_09748_),
    .Y(_09750_));
 sky130_as_sc_hs__and2_2 _40492_ (.A(_09749_),
    .B(_09750_),
    .Y(_09751_));
 sky130_as_sc_hs__or2_2 _40494_ (.A(_09738_),
    .B(_09751_),
    .Y(_09753_));
 sky130_as_sc_hs__and2_2 _40495_ (.A(_09752_),
    .B(_09753_),
    .Y(_09754_));
 sky130_as_sc_hs__or2_2 _40497_ (.A(_09737_),
    .B(_09754_),
    .Y(_09756_));
 sky130_as_sc_hs__and2_2 _40498_ (.A(_09755_),
    .B(_09756_),
    .Y(_09757_));
 sky130_as_sc_hs__or2_2 _40501_ (.A(_09757_),
    .B(_09758_),
    .Y(_09760_));
 sky130_as_sc_hs__and2_2 _40502_ (.A(_09759_),
    .B(_09760_),
    .Y(_09761_));
 sky130_as_sc_hs__and2_2 _40505_ (.A(net481),
    .B(net426),
    .Y(_09764_));
 sky130_as_sc_hs__and2_2 _40506_ (.A(_24527_),
    .B(net424),
    .Y(_09765_));
 sky130_as_sc_hs__and2_2 _40507_ (.A(net89),
    .B(net419),
    .Y(_09766_));
 sky130_as_sc_hs__or2_2 _40508_ (.A(_09765_),
    .B(_09766_),
    .Y(_09767_));
 sky130_as_sc_hs__and2_2 _40510_ (.A(_09767_),
    .B(_09768_),
    .Y(_09769_));
 sky130_as_sc_hs__and2_2 _40511_ (.A(net88),
    .B(net74),
    .Y(_09770_));
 sky130_as_sc_hs__or2_2 _40513_ (.A(_09769_),
    .B(_09770_),
    .Y(_09772_));
 sky130_as_sc_hs__and2_2 _40514_ (.A(_09771_),
    .B(_09772_),
    .Y(_09773_));
 sky130_as_sc_hs__or2_2 _40517_ (.A(_09773_),
    .B(_09774_),
    .Y(_09776_));
 sky130_as_sc_hs__and2_2 _40518_ (.A(_09775_),
    .B(_09776_),
    .Y(_09777_));
 sky130_as_sc_hs__or2_2 _40520_ (.A(_09764_),
    .B(_09777_),
    .Y(_09779_));
 sky130_as_sc_hs__and2_2 _40521_ (.A(_09778_),
    .B(_09779_),
    .Y(_09780_));
 sky130_as_sc_hs__or2_2 _40523_ (.A(_09763_),
    .B(_09780_),
    .Y(_09782_));
 sky130_as_sc_hs__and2_2 _40524_ (.A(_09781_),
    .B(_09782_),
    .Y(_09783_));
 sky130_as_sc_hs__or2_2 _40526_ (.A(_09762_),
    .B(_09783_),
    .Y(_09785_));
 sky130_as_sc_hs__and2_2 _40527_ (.A(_09784_),
    .B(_09785_),
    .Y(_09786_));
 sky130_as_sc_hs__or2_2 _40529_ (.A(_09761_),
    .B(_09786_),
    .Y(_09788_));
 sky130_as_sc_hs__and2_2 _40530_ (.A(_09787_),
    .B(_09788_),
    .Y(_09789_));
 sky130_as_sc_hs__or2_2 _40533_ (.A(_09789_),
    .B(_09790_),
    .Y(_09792_));
 sky130_as_sc_hs__and2_2 _40534_ (.A(_09791_),
    .B(_09792_),
    .Y(_09793_));
 sky130_as_sc_hs__and2_2 _40537_ (.A(net478),
    .B(net440),
    .Y(_09796_));
 sky130_as_sc_hs__and2_2 _40538_ (.A(net474),
    .B(net436),
    .Y(_09797_));
 sky130_as_sc_hs__and2_2 _40539_ (.A(_09796_),
    .B(_09797_),
    .Y(_09798_));
 sky130_as_sc_hs__or2_2 _40540_ (.A(_09796_),
    .B(_09797_),
    .Y(_09799_));
 sky130_as_sc_hs__nor2b_2 _40541_ (.A(_09798_),
    .Y(_09800_),
    .B(_09799_));
 sky130_as_sc_hs__nor2_2 _40543_ (.A(_09549_),
    .B(_09801_),
    .Y(_09802_));
 sky130_as_sc_hs__and2_2 _40544_ (.A(_09549_),
    .B(_09801_),
    .Y(_09803_));
 sky130_as_sc_hs__or2_2 _40545_ (.A(_09802_),
    .B(_09803_),
    .Y(_09804_));
 sky130_as_sc_hs__or2_2 _40546_ (.A(_09476_),
    .B(_09804_),
    .Y(_09805_));
 sky130_as_sc_hs__and2_2 _40548_ (.A(_09805_),
    .B(_09806_),
    .Y(_09807_));
 sky130_as_sc_hs__or2_2 _40550_ (.A(_09800_),
    .B(_09807_),
    .Y(_09809_));
 sky130_as_sc_hs__and2_2 _40551_ (.A(_09808_),
    .B(_09809_),
    .Y(_09810_));
 sky130_as_sc_hs__or2_2 _40553_ (.A(_09795_),
    .B(_09810_),
    .Y(_09812_));
 sky130_as_sc_hs__and2_2 _40554_ (.A(_09811_),
    .B(_09812_),
    .Y(_09813_));
 sky130_as_sc_hs__or2_2 _40556_ (.A(_09794_),
    .B(_09813_),
    .Y(_09815_));
 sky130_as_sc_hs__and2_2 _40557_ (.A(_09814_),
    .B(_09815_),
    .Y(_09816_));
 sky130_as_sc_hs__or2_2 _40559_ (.A(_09793_),
    .B(_09816_),
    .Y(_09818_));
 sky130_as_sc_hs__and2_2 _40560_ (.A(_09817_),
    .B(_09818_),
    .Y(_09819_));
 sky130_as_sc_hs__or2_2 _40563_ (.A(_09819_),
    .B(_09820_),
    .Y(_09822_));
 sky130_as_sc_hs__and2_2 _40564_ (.A(_09821_),
    .B(_09822_),
    .Y(_09823_));
 sky130_as_sc_hs__or2_2 _40566_ (.A(_09708_),
    .B(_09823_),
    .Y(_09825_));
 sky130_as_sc_hs__and2_2 _40567_ (.A(_09824_),
    .B(_09825_),
    .Y(_09826_));
 sky130_as_sc_hs__or2_2 _40570_ (.A(_09826_),
    .B(_09827_),
    .Y(_09829_));
 sky130_as_sc_hs__and2_2 _40571_ (.A(_09828_),
    .B(_09829_),
    .Y(_09830_));
 sky130_as_sc_hs__or2_2 _40573_ (.A(_09689_),
    .B(_09830_),
    .Y(_09832_));
 sky130_as_sc_hs__and2_2 _40574_ (.A(_09831_),
    .B(_09832_),
    .Y(_09833_));
 sky130_as_sc_hs__or2_2 _40576_ (.A(_09688_),
    .B(_09833_),
    .Y(_09835_));
 sky130_as_sc_hs__and2_2 _40577_ (.A(_09834_),
    .B(_09835_),
    .Y(_09836_));
 sky130_as_sc_hs__or2_2 _40579_ (.A(_09687_),
    .B(_09836_),
    .Y(_09838_));
 sky130_as_sc_hs__and2_2 _40580_ (.A(_09837_),
    .B(_09838_),
    .Y(_09839_));
 sky130_as_sc_hs__and2_2 _40581_ (.A(_09606_),
    .B(_09617_),
    .Y(_09840_));
 sky130_as_sc_hs__or2_2 _40583_ (.A(_09839_),
    .B(_09840_),
    .Y(_09842_));
 sky130_as_sc_hs__and2_2 _40584_ (.A(_09841_),
    .B(_09842_),
    .Y(_09843_));
 sky130_as_sc_hs__or2_2 _40587_ (.A(_09843_),
    .B(_09844_),
    .Y(_09846_));
 sky130_as_sc_hs__nand3_2 _40588_ (.A(net141),
    .B(_09845_),
    .C(_09846_),
    .Y(_09847_));
 sky130_as_sc_hs__or2_2 _40591_ (.A(_05423_),
    .B(_09848_),
    .Y(_09850_));
 sky130_as_sc_hs__nand3_2 _40592_ (.A(net138),
    .B(_09849_),
    .C(_09850_),
    .Y(_09851_));
 sky130_as_sc_hs__and2_2 _40593_ (.A(_05704_),
    .B(_09631_),
    .Y(_09852_));
 sky130_as_sc_hs__or2_2 _40594_ (.A(_05696_),
    .B(_09852_),
    .Y(_09853_));
 sky130_as_sc_hs__or2_2 _40598_ (.A(_05696_),
    .B(_05875_),
    .Y(_09857_));
 sky130_as_sc_hs__nand3_2 _40601_ (.A(net119),
    .B(_09856_),
    .C(_09859_),
    .Y(_09860_));
 sky130_as_sc_hs__or2_2 _40602_ (.A(_05935_),
    .B(_07809_),
    .Y(_09861_));
 sky130_as_sc_hs__nand3_2 _40604_ (.A(_05929_),
    .B(_09861_),
    .C(_09862_),
    .Y(_09863_));
 sky130_as_sc_hs__or2_2 _40605_ (.A(_05929_),
    .B(_06908_),
    .Y(_09864_));
 sky130_as_sc_hs__and2_2 _40606_ (.A(_09863_),
    .B(_09864_),
    .Y(_09865_));
 sky130_as_sc_hs__and2_2 _40610_ (.A(net140),
    .B(_09868_),
    .Y(_09869_));
 sky130_as_sc_hs__or2_2 _40611_ (.A(\tholin_riscv.div_res[12] ),
    .B(_09648_),
    .Y(_09870_));
 sky130_as_sc_hs__and2_2 _40612_ (.A(net414),
    .B(_09870_),
    .Y(_09871_));
 sky130_as_sc_hs__or2_2 _40613_ (.A(\tholin_riscv.div_res[13] ),
    .B(_09871_),
    .Y(_09872_));
 sky130_as_sc_hs__nand3_2 _40615_ (.A(net110),
    .B(_09872_),
    .C(_09873_),
    .Y(_09874_));
 sky130_as_sc_hs__or2_2 _40616_ (.A(\tholin_riscv.div_shifter[44] ),
    .B(_09656_),
    .Y(_09875_));
 sky130_as_sc_hs__and2_2 _40617_ (.A(_21655_),
    .B(_09875_),
    .Y(_09876_));
 sky130_as_sc_hs__or2_2 _40619_ (.A(\tholin_riscv.div_shifter[45] ),
    .B(_09876_),
    .Y(_09878_));
 sky130_as_sc_hs__nand3_2 _40620_ (.A(net108),
    .B(_09877_),
    .C(_09878_),
    .Y(_09879_));
 sky130_as_sc_hs__nor2_2 _40624_ (.A(_05694_),
    .B(_06161_),
    .Y(_09883_));
 sky130_as_sc_hs__nand3_2 _40627_ (.A(net413),
    .B(_09884_),
    .C(_09885_),
    .Y(_09886_));
 sky130_as_sc_hs__nor2_2 _40628_ (.A(_09883_),
    .B(_09886_),
    .Y(_09887_));
 sky130_as_sc_hs__and2_2 _40629_ (.A(_09882_),
    .B(_09887_),
    .Y(_09888_));
 sky130_as_sc_hs__nand3_2 _40630_ (.A(_09874_),
    .B(_09879_),
    .C(_09888_),
    .Y(_09889_));
 sky130_as_sc_hs__nor2_2 _40631_ (.A(_09869_),
    .B(_09889_),
    .Y(_09890_));
 sky130_as_sc_hs__and2_2 _40632_ (.A(_09866_),
    .B(_09890_),
    .Y(_09891_));
 sky130_as_sc_hs__and2_2 _40633_ (.A(_09860_),
    .B(_09891_),
    .Y(_09892_));
 sky130_as_sc_hs__nand3_2 _40634_ (.A(_09847_),
    .B(_09851_),
    .C(_09892_),
    .Y(_09893_));
 sky130_as_sc_hs__and2_2 _40635_ (.A(\tholin_riscv.PC[13] ),
    .B(_09672_),
    .Y(_09894_));
 sky130_as_sc_hs__nor2_2 _40636_ (.A(\tholin_riscv.PC[13] ),
    .B(_09672_),
    .Y(_09895_));
 sky130_as_sc_hs__or2_2 _40637_ (.A(_09894_),
    .B(_09895_),
    .Y(_09896_));
 sky130_as_sc_hs__nor2_2 _40638_ (.A(_21572_),
    .B(_09896_),
    .Y(_09897_));
 sky130_as_sc_hs__and2_2 _40640_ (.A(\tholin_riscv.PC[12] ),
    .B(\tholin_riscv.Jimm[12] ),
    .Y(_09899_));
 sky130_as_sc_hs__or2_2 _40642_ (.A(\tholin_riscv.PC[13] ),
    .B(\tholin_riscv.Jimm[13] ),
    .Y(_09901_));
 sky130_as_sc_hs__and2_2 _40643_ (.A(_09900_),
    .B(_09901_),
    .Y(_09902_));
 sky130_as_sc_hs__or2_2 _40645_ (.A(_09899_),
    .B(_09902_),
    .Y(_09904_));
 sky130_as_sc_hs__nand3_2 _40646_ (.A(net117),
    .B(_09903_),
    .C(_09904_),
    .Y(_09905_));
 sky130_as_sc_hs__nand3_2 _40647_ (.A(_21569_),
    .B(_09898_),
    .C(_09905_),
    .Y(_09906_));
 sky130_as_sc_hs__or2_2 _40648_ (.A(_09897_),
    .B(_09906_),
    .Y(_09907_));
 sky130_as_sc_hs__nand3_2 _40649_ (.A(_21546_),
    .B(_09893_),
    .C(_09907_),
    .Y(_09908_));
 sky130_as_sc_hs__or2_2 _40654_ (.A(_19867_),
    .B(_08428_),
    .Y(_09912_));
 sky130_as_sc_hs__and2_2 _40657_ (.A(net442),
    .B(_02550_),
    .Y(_09915_));
 sky130_as_sc_hs__and2_2 _40658_ (.A(net438),
    .B(net433),
    .Y(_09916_));
 sky130_as_sc_hs__or2_2 _40659_ (.A(_09915_),
    .B(_09916_),
    .Y(_09917_));
 sky130_as_sc_hs__and2_2 _40661_ (.A(_09917_),
    .B(_09918_),
    .Y(_09919_));
 sky130_as_sc_hs__and2_2 _40662_ (.A(net478),
    .B(net456),
    .Y(_09920_));
 sky130_as_sc_hs__or2_2 _40664_ (.A(_09919_),
    .B(_09920_),
    .Y(_09922_));
 sky130_as_sc_hs__and2_2 _40665_ (.A(_09921_),
    .B(_09922_),
    .Y(_09923_));
 sky130_as_sc_hs__or2_2 _40668_ (.A(_09923_),
    .B(_09924_),
    .Y(_09926_));
 sky130_as_sc_hs__and2_2 _40669_ (.A(_09925_),
    .B(_09926_),
    .Y(_09927_));
 sky130_as_sc_hs__and2_2 _40670_ (.A(net466),
    .B(net431),
    .Y(_09928_));
 sky130_as_sc_hs__and2_2 _40671_ (.A(net468),
    .B(net429),
    .Y(_09929_));
 sky130_as_sc_hs__or2_2 _40672_ (.A(_09928_),
    .B(_09929_),
    .Y(_09930_));
 sky130_as_sc_hs__and2_2 _40674_ (.A(_09930_),
    .B(_09931_),
    .Y(_09932_));
 sky130_as_sc_hs__and2_2 _40675_ (.A(net471),
    .B(net427),
    .Y(_09933_));
 sky130_as_sc_hs__or2_2 _40677_ (.A(_09932_),
    .B(_09933_),
    .Y(_09935_));
 sky130_as_sc_hs__and2_2 _40678_ (.A(_09934_),
    .B(_09935_),
    .Y(_09936_));
 sky130_as_sc_hs__or2_2 _40680_ (.A(_09927_),
    .B(_09936_),
    .Y(_09938_));
 sky130_as_sc_hs__and2_2 _40681_ (.A(_09937_),
    .B(_09938_),
    .Y(_09939_));
 sky130_as_sc_hs__or2_2 _40684_ (.A(_09939_),
    .B(_09940_),
    .Y(_09942_));
 sky130_as_sc_hs__and2_2 _40685_ (.A(_09941_),
    .B(_09942_),
    .Y(_09943_));
 sky130_as_sc_hs__and2_2 _40688_ (.A(net120),
    .B(net465),
    .Y(_09946_));
 sky130_as_sc_hs__and2_2 _40689_ (.A(net122),
    .B(net463),
    .Y(_09947_));
 sky130_as_sc_hs__or2_2 _40690_ (.A(_09946_),
    .B(_09947_),
    .Y(_09948_));
 sky130_as_sc_hs__and2_2 _40692_ (.A(_09948_),
    .B(_09949_),
    .Y(_09950_));
 sky130_as_sc_hs__and2_2 _40693_ (.A(net460),
    .B(net424),
    .Y(_09951_));
 sky130_as_sc_hs__or2_2 _40695_ (.A(_09950_),
    .B(_09951_),
    .Y(_09953_));
 sky130_as_sc_hs__and2_2 _40696_ (.A(_09952_),
    .B(_09953_),
    .Y(_09954_));
 sky130_as_sc_hs__or2_2 _40698_ (.A(_09945_),
    .B(_09954_),
    .Y(_09956_));
 sky130_as_sc_hs__and2_2 _40699_ (.A(_09955_),
    .B(_09956_),
    .Y(_09957_));
 sky130_as_sc_hs__or2_2 _40701_ (.A(_09944_),
    .B(_09957_),
    .Y(_09959_));
 sky130_as_sc_hs__and2_2 _40702_ (.A(_09958_),
    .B(_09959_),
    .Y(_09960_));
 sky130_as_sc_hs__or2_2 _40704_ (.A(_09943_),
    .B(_09960_),
    .Y(_09962_));
 sky130_as_sc_hs__and2_2 _40705_ (.A(_09961_),
    .B(_09962_),
    .Y(_09963_));
 sky130_as_sc_hs__or2_2 _40708_ (.A(_09963_),
    .B(_09964_),
    .Y(_09966_));
 sky130_as_sc_hs__and2_2 _40709_ (.A(_09965_),
    .B(_09966_),
    .Y(_09967_));
 sky130_as_sc_hs__and2_2 _40712_ (.A(net476),
    .B(net425),
    .Y(_09970_));
 sky130_as_sc_hs__and2_2 _40713_ (.A(_24527_),
    .B(net419),
    .Y(_09971_));
 sky130_as_sc_hs__and2_2 _40714_ (.A(net89),
    .B(net74),
    .Y(_09972_));
 sky130_as_sc_hs__or2_2 _40715_ (.A(_09971_),
    .B(_09972_),
    .Y(_09973_));
 sky130_as_sc_hs__and2_2 _40717_ (.A(_09973_),
    .B(_09974_),
    .Y(_09975_));
 sky130_as_sc_hs__or2_2 _40720_ (.A(_09975_),
    .B(_09976_),
    .Y(_09978_));
 sky130_as_sc_hs__and2_2 _40721_ (.A(_09977_),
    .B(_09978_),
    .Y(_09979_));
 sky130_as_sc_hs__or2_2 _40723_ (.A(_09970_),
    .B(_09979_),
    .Y(_09981_));
 sky130_as_sc_hs__and2_2 _40724_ (.A(_09980_),
    .B(_09981_),
    .Y(_09982_));
 sky130_as_sc_hs__or2_2 _40726_ (.A(_09969_),
    .B(_09982_),
    .Y(_09984_));
 sky130_as_sc_hs__and2_2 _40727_ (.A(_09983_),
    .B(_09984_),
    .Y(_09985_));
 sky130_as_sc_hs__or2_2 _40729_ (.A(_09968_),
    .B(_09985_),
    .Y(_09987_));
 sky130_as_sc_hs__and2_2 _40730_ (.A(_09986_),
    .B(_09987_),
    .Y(_09988_));
 sky130_as_sc_hs__or2_2 _40732_ (.A(_09967_),
    .B(_09988_),
    .Y(_09990_));
 sky130_as_sc_hs__and2_2 _40733_ (.A(_09989_),
    .B(_09990_),
    .Y(_09991_));
 sky130_as_sc_hs__or2_2 _40736_ (.A(_09991_),
    .B(_09992_),
    .Y(_09994_));
 sky130_as_sc_hs__and2_2 _40737_ (.A(_09993_),
    .B(_09994_),
    .Y(_09995_));
 sky130_as_sc_hs__and2_2 _40740_ (.A(net475),
    .B(net440),
    .Y(_09998_));
 sky130_as_sc_hs__and2_2 _40741_ (.A(net437),
    .B(net83),
    .Y(_09999_));
 sky130_as_sc_hs__and2_2 _40742_ (.A(_09998_),
    .B(_09999_),
    .Y(_10000_));
 sky130_as_sc_hs__or2_2 _40743_ (.A(_09998_),
    .B(_09999_),
    .Y(_10001_));
 sky130_as_sc_hs__nor2b_2 _40744_ (.A(_10000_),
    .Y(_10002_),
    .B(_10001_));
 sky130_as_sc_hs__and2_2 _40745_ (.A(net472),
    .B(net434),
    .Y(_10003_));
 sky130_as_sc_hs__or2_2 _40746_ (.A(_09802_),
    .B(_10003_),
    .Y(_10004_));
 sky130_as_sc_hs__and2_2 _40748_ (.A(_10004_),
    .B(_10005_),
    .Y(_10006_));
 sky130_as_sc_hs__or2_2 _40750_ (.A(_10002_),
    .B(_10006_),
    .Y(_10008_));
 sky130_as_sc_hs__and2_2 _40751_ (.A(_10007_),
    .B(_10008_),
    .Y(_10009_));
 sky130_as_sc_hs__or2_2 _40753_ (.A(_09997_),
    .B(_10009_),
    .Y(_10011_));
 sky130_as_sc_hs__and2_2 _40754_ (.A(_10010_),
    .B(_10011_),
    .Y(_10012_));
 sky130_as_sc_hs__or2_2 _40756_ (.A(_09996_),
    .B(_10012_),
    .Y(_10014_));
 sky130_as_sc_hs__and2_2 _40757_ (.A(_10013_),
    .B(_10014_),
    .Y(_10015_));
 sky130_as_sc_hs__or2_2 _40759_ (.A(_09995_),
    .B(_10015_),
    .Y(_10017_));
 sky130_as_sc_hs__and2_2 _40760_ (.A(_10016_),
    .B(_10017_),
    .Y(_10018_));
 sky130_as_sc_hs__or2_2 _40763_ (.A(_10018_),
    .B(_10019_),
    .Y(_10021_));
 sky130_as_sc_hs__and2_2 _40764_ (.A(_10020_),
    .B(_10021_),
    .Y(_10022_));
 sky130_as_sc_hs__and2_2 _40767_ (.A(_23674_),
    .B(net128),
    .Y(_10025_));
 sky130_as_sc_hs__or2_2 _40769_ (.A(_09798_),
    .B(_10025_),
    .Y(_10027_));
 sky130_as_sc_hs__or2_2 _40771_ (.A(_09693_),
    .B(_10028_),
    .Y(_10029_));
 sky130_as_sc_hs__and2_2 _40773_ (.A(_10029_),
    .B(_10030_),
    .Y(_10031_));
 sky130_as_sc_hs__and2_2 _40774_ (.A(net480),
    .B(net421),
    .Y(_10032_));
 sky130_as_sc_hs__or2_2 _40776_ (.A(_10031_),
    .B(_10032_),
    .Y(_10034_));
 sky130_as_sc_hs__and2_2 _40777_ (.A(_10033_),
    .B(_10034_),
    .Y(_10035_));
 sky130_as_sc_hs__or2_2 _40779_ (.A(_10024_),
    .B(_10035_),
    .Y(_10037_));
 sky130_as_sc_hs__and2_2 _40780_ (.A(_10036_),
    .B(_10037_),
    .Y(_10038_));
 sky130_as_sc_hs__or2_2 _40782_ (.A(_10023_),
    .B(_10038_),
    .Y(_10040_));
 sky130_as_sc_hs__and2_2 _40783_ (.A(_10039_),
    .B(_10040_),
    .Y(_10041_));
 sky130_as_sc_hs__or2_2 _40785_ (.A(_10022_),
    .B(_10041_),
    .Y(_10043_));
 sky130_as_sc_hs__and2_2 _40786_ (.A(_10042_),
    .B(_10043_),
    .Y(_10044_));
 sky130_as_sc_hs__or2_2 _40789_ (.A(_10044_),
    .B(_10045_),
    .Y(_10047_));
 sky130_as_sc_hs__and2_2 _40790_ (.A(_10046_),
    .B(_10047_),
    .Y(_10048_));
 sky130_as_sc_hs__or2_2 _40792_ (.A(_09914_),
    .B(_10048_),
    .Y(_10050_));
 sky130_as_sc_hs__and2_2 _40793_ (.A(_10049_),
    .B(_10050_),
    .Y(_10051_));
 sky130_as_sc_hs__or2_2 _40796_ (.A(_10051_),
    .B(_10052_),
    .Y(_10054_));
 sky130_as_sc_hs__or2_2 _40798_ (.A(_09834_),
    .B(_10055_),
    .Y(_10056_));
 sky130_as_sc_hs__and2_2 _40800_ (.A(_10056_),
    .B(_10057_),
    .Y(_10058_));
 sky130_as_sc_hs__and2_2 _40803_ (.A(_09608_),
    .B(_09839_),
    .Y(_10061_));
 sky130_as_sc_hs__or2_2 _40807_ (.A(_10058_),
    .B(_10063_),
    .Y(_10065_));
 sky130_as_sc_hs__and2_2 _40808_ (.A(_10064_),
    .B(_10065_),
    .Y(_10066_));
 sky130_as_sc_hs__and2_2 _40809_ (.A(_09619_),
    .B(_09843_),
    .Y(_10067_));
 sky130_as_sc_hs__or2_2 _40814_ (.A(_10066_),
    .B(_10070_),
    .Y(_10072_));
 sky130_as_sc_hs__nand3_2 _40815_ (.A(net141),
    .B(_10071_),
    .C(_10072_),
    .Y(_10073_));
 sky130_as_sc_hs__or2_2 _40816_ (.A(_05424_),
    .B(_05505_),
    .Y(_10074_));
 sky130_as_sc_hs__or2_2 _40817_ (.A(_05384_),
    .B(_10074_),
    .Y(_10075_));
 sky130_as_sc_hs__nand3_2 _40819_ (.A(net138),
    .B(_10075_),
    .C(_10076_),
    .Y(_10077_));
 sky130_as_sc_hs__and2_2 _40820_ (.A(_05694_),
    .B(_09853_),
    .Y(_10078_));
 sky130_as_sc_hs__or2_2 _40821_ (.A(_05686_),
    .B(_10078_),
    .Y(_10079_));
 sky130_as_sc_hs__or2_2 _40825_ (.A(_05686_),
    .B(_05877_),
    .Y(_10083_));
 sky130_as_sc_hs__nand3_2 _40828_ (.A(net118),
    .B(_10082_),
    .C(_10085_),
    .Y(_10086_));
 sky130_as_sc_hs__or2_2 _40829_ (.A(_05935_),
    .B(_08099_),
    .Y(_10087_));
 sky130_as_sc_hs__nand3_2 _40831_ (.A(_05929_),
    .B(_10087_),
    .C(_10088_),
    .Y(_10089_));
 sky130_as_sc_hs__or2_2 _40832_ (.A(_05929_),
    .B(_06431_),
    .Y(_10090_));
 sky130_as_sc_hs__and2_2 _40833_ (.A(_10089_),
    .B(_10090_),
    .Y(_10091_));
 sky130_as_sc_hs__and2_2 _40837_ (.A(net140),
    .B(_10094_),
    .Y(_10095_));
 sky130_as_sc_hs__or2_2 _40838_ (.A(\tholin_riscv.div_shifter[45] ),
    .B(_09875_),
    .Y(_10096_));
 sky130_as_sc_hs__and2_2 _40839_ (.A(_21655_),
    .B(_10096_),
    .Y(_10097_));
 sky130_as_sc_hs__or2_2 _40840_ (.A(\tholin_riscv.div_shifter[46] ),
    .B(_10097_),
    .Y(_10098_));
 sky130_as_sc_hs__nand3_2 _40842_ (.A(net107),
    .B(_10098_),
    .C(_10099_),
    .Y(_10100_));
 sky130_as_sc_hs__or2_2 _40843_ (.A(\tholin_riscv.div_res[13] ),
    .B(_09870_),
    .Y(_10101_));
 sky130_as_sc_hs__and2_2 _40844_ (.A(net414),
    .B(_10101_),
    .Y(_10102_));
 sky130_as_sc_hs__or2_2 _40845_ (.A(\tholin_riscv.div_res[14] ),
    .B(_10102_),
    .Y(_10103_));
 sky130_as_sc_hs__nand3_2 _40847_ (.A(net110),
    .B(_10103_),
    .C(_10104_),
    .Y(_10105_));
 sky130_as_sc_hs__nor2_2 _40851_ (.A(_05684_),
    .B(_06161_),
    .Y(_10109_));
 sky130_as_sc_hs__nand3_2 _40854_ (.A(net412),
    .B(_10110_),
    .C(_10111_),
    .Y(_10112_));
 sky130_as_sc_hs__nor2_2 _40855_ (.A(_10109_),
    .B(_10112_),
    .Y(_10113_));
 sky130_as_sc_hs__and2_2 _40856_ (.A(_10108_),
    .B(_10113_),
    .Y(_10114_));
 sky130_as_sc_hs__nand3_2 _40857_ (.A(_10100_),
    .B(_10105_),
    .C(_10114_),
    .Y(_10115_));
 sky130_as_sc_hs__nor2_2 _40858_ (.A(_10095_),
    .B(_10115_),
    .Y(_10116_));
 sky130_as_sc_hs__and2_2 _40859_ (.A(_10092_),
    .B(_10116_),
    .Y(_10117_));
 sky130_as_sc_hs__and2_2 _40860_ (.A(_10086_),
    .B(_10117_),
    .Y(_10118_));
 sky130_as_sc_hs__nand3_2 _40861_ (.A(_10073_),
    .B(_10077_),
    .C(_10118_),
    .Y(_10119_));
 sky130_as_sc_hs__and2_2 _40862_ (.A(\tholin_riscv.PC[14] ),
    .B(_09894_),
    .Y(_10120_));
 sky130_as_sc_hs__nor2_2 _40863_ (.A(\tholin_riscv.PC[14] ),
    .B(_09894_),
    .Y(_10121_));
 sky130_as_sc_hs__or2_2 _40864_ (.A(_10120_),
    .B(_10121_),
    .Y(_10122_));
 sky130_as_sc_hs__or2_2 _40866_ (.A(\tholin_riscv.Jimm[14] ),
    .B(_21590_),
    .Y(_10124_));
 sky130_as_sc_hs__or2_2 _40869_ (.A(\tholin_riscv.PC[14] ),
    .B(net411),
    .Y(_10127_));
 sky130_as_sc_hs__or2_2 _40871_ (.A(_10125_),
    .B(_10128_),
    .Y(_10129_));
 sky130_as_sc_hs__nand3_2 _40873_ (.A(net117),
    .B(_10129_),
    .C(_10130_),
    .Y(_10131_));
 sky130_as_sc_hs__nand3_2 _40874_ (.A(_10123_),
    .B(_10124_),
    .C(_10131_),
    .Y(_10132_));
 sky130_as_sc_hs__nand3_2 _40876_ (.A(_21546_),
    .B(_10119_),
    .C(_10133_),
    .Y(_10134_));
 sky130_as_sc_hs__or2_2 _40881_ (.A(_19875_),
    .B(_08428_),
    .Y(_10138_));
 sky130_as_sc_hs__and2_2 _40883_ (.A(_10056_),
    .B(_10064_),
    .Y(_10140_));
 sky130_as_sc_hs__and2_2 _40884_ (.A(_23674_),
    .B(net418),
    .Y(_10141_));
 sky130_as_sc_hs__and2_2 _40885_ (.A(net472),
    .B(net433),
    .Y(_10142_));
 sky130_as_sc_hs__or2_2 _40886_ (.A(_10141_),
    .B(_10142_),
    .Y(_10143_));
 sky130_as_sc_hs__and2_2 _40888_ (.A(_10143_),
    .B(_10144_),
    .Y(_10145_));
 sky130_as_sc_hs__and2_2 _40889_ (.A(net474),
    .B(net457),
    .Y(_10146_));
 sky130_as_sc_hs__or2_2 _40891_ (.A(_10145_),
    .B(_10146_),
    .Y(_10148_));
 sky130_as_sc_hs__and2_2 _40892_ (.A(_10147_),
    .B(_10148_),
    .Y(_10149_));
 sky130_as_sc_hs__or2_2 _40895_ (.A(_10149_),
    .B(_10150_),
    .Y(_10152_));
 sky130_as_sc_hs__and2_2 _40896_ (.A(_10151_),
    .B(_10152_),
    .Y(_10153_));
 sky130_as_sc_hs__and2_2 _40897_ (.A(net466),
    .B(net429),
    .Y(_10154_));
 sky130_as_sc_hs__and2_2 _40898_ (.A(net468),
    .B(net427),
    .Y(_10155_));
 sky130_as_sc_hs__or2_2 _40899_ (.A(_10154_),
    .B(_10155_),
    .Y(_10156_));
 sky130_as_sc_hs__and2_2 _40901_ (.A(_10156_),
    .B(_10157_),
    .Y(_10158_));
 sky130_as_sc_hs__and2_2 _40902_ (.A(net120),
    .B(net471),
    .Y(_10159_));
 sky130_as_sc_hs__or2_2 _40904_ (.A(_10158_),
    .B(_10159_),
    .Y(_10161_));
 sky130_as_sc_hs__and2_2 _40905_ (.A(_10160_),
    .B(_10161_),
    .Y(_10162_));
 sky130_as_sc_hs__or2_2 _40907_ (.A(_10153_),
    .B(_10162_),
    .Y(_10164_));
 sky130_as_sc_hs__and2_2 _40908_ (.A(_10163_),
    .B(_10164_),
    .Y(_10165_));
 sky130_as_sc_hs__or2_2 _40911_ (.A(_10165_),
    .B(_10166_),
    .Y(_10168_));
 sky130_as_sc_hs__and2_2 _40912_ (.A(_10167_),
    .B(_10168_),
    .Y(_10169_));
 sky130_as_sc_hs__and2_2 _40915_ (.A(net122),
    .B(net465),
    .Y(_10172_));
 sky130_as_sc_hs__and2_2 _40916_ (.A(net463),
    .B(net423),
    .Y(_10173_));
 sky130_as_sc_hs__or2_2 _40917_ (.A(_10172_),
    .B(_10173_),
    .Y(_10174_));
 sky130_as_sc_hs__and2_2 _40919_ (.A(_10174_),
    .B(_10175_),
    .Y(_10176_));
 sky130_as_sc_hs__and2_2 _40920_ (.A(net460),
    .B(net419),
    .Y(_10177_));
 sky130_as_sc_hs__or2_2 _40922_ (.A(_10176_),
    .B(_10177_),
    .Y(_10179_));
 sky130_as_sc_hs__and2_2 _40923_ (.A(_10178_),
    .B(_10179_),
    .Y(_10180_));
 sky130_as_sc_hs__or2_2 _40925_ (.A(_10171_),
    .B(_10180_),
    .Y(_10182_));
 sky130_as_sc_hs__and2_2 _40926_ (.A(_10181_),
    .B(_10182_),
    .Y(_10183_));
 sky130_as_sc_hs__or2_2 _40928_ (.A(_10170_),
    .B(_10183_),
    .Y(_10185_));
 sky130_as_sc_hs__and2_2 _40929_ (.A(_10184_),
    .B(_10185_),
    .Y(_10186_));
 sky130_as_sc_hs__or2_2 _40931_ (.A(_10169_),
    .B(_10186_),
    .Y(_10188_));
 sky130_as_sc_hs__and2_2 _40932_ (.A(_10187_),
    .B(_10188_),
    .Y(_10189_));
 sky130_as_sc_hs__or2_2 _40935_ (.A(_10189_),
    .B(_10190_),
    .Y(_10192_));
 sky130_as_sc_hs__and2_2 _40936_ (.A(_10191_),
    .B(_10192_),
    .Y(_10193_));
 sky130_as_sc_hs__and2_2 _40939_ (.A(net438),
    .B(net425),
    .Y(_10196_));
 sky130_as_sc_hs__nor2_2 _40941_ (.A(_09766_),
    .B(_10197_),
    .Y(_10198_));
 sky130_as_sc_hs__or2_2 _40943_ (.A(_10196_),
    .B(_10198_),
    .Y(_10200_));
 sky130_as_sc_hs__and2_2 _40944_ (.A(_10199_),
    .B(_10200_),
    .Y(_10201_));
 sky130_as_sc_hs__or2_2 _40946_ (.A(_10195_),
    .B(_10201_),
    .Y(_10203_));
 sky130_as_sc_hs__and2_2 _40947_ (.A(_10202_),
    .B(_10203_),
    .Y(_10204_));
 sky130_as_sc_hs__or2_2 _40949_ (.A(_10194_),
    .B(_10204_),
    .Y(_10206_));
 sky130_as_sc_hs__and2_2 _40950_ (.A(_10205_),
    .B(_10206_),
    .Y(_10207_));
 sky130_as_sc_hs__or2_2 _40952_ (.A(_10193_),
    .B(_10207_),
    .Y(_10209_));
 sky130_as_sc_hs__and2_2 _40953_ (.A(_10208_),
    .B(_10209_),
    .Y(_10210_));
 sky130_as_sc_hs__or2_2 _40956_ (.A(_10210_),
    .B(_10211_),
    .Y(_10213_));
 sky130_as_sc_hs__and2_2 _40957_ (.A(_10212_),
    .B(_10213_),
    .Y(_10214_));
 sky130_as_sc_hs__and2_2 _40960_ (.A(net478),
    .B(net434),
    .Y(_10217_));
 sky130_as_sc_hs__and2_2 _40961_ (.A(net440),
    .B(net83),
    .Y(_10218_));
 sky130_as_sc_hs__and2_2 _40962_ (.A(net436),
    .B(net432),
    .Y(_10219_));
 sky130_as_sc_hs__and2_2 _40963_ (.A(_10218_),
    .B(_10219_),
    .Y(_10220_));
 sky130_as_sc_hs__or2_2 _40964_ (.A(_10218_),
    .B(_10219_),
    .Y(_10221_));
 sky130_as_sc_hs__nor2b_2 _40965_ (.A(_10220_),
    .Y(_10222_),
    .B(_10221_));
 sky130_as_sc_hs__or2_2 _40967_ (.A(_10217_),
    .B(_10222_),
    .Y(_10224_));
 sky130_as_sc_hs__and2_2 _40968_ (.A(_10223_),
    .B(_10224_),
    .Y(_10225_));
 sky130_as_sc_hs__or2_2 _40970_ (.A(_10216_),
    .B(_10225_),
    .Y(_10227_));
 sky130_as_sc_hs__and2_2 _40971_ (.A(_10226_),
    .B(_10227_),
    .Y(_10228_));
 sky130_as_sc_hs__or2_2 _40973_ (.A(_10215_),
    .B(_10228_),
    .Y(_10230_));
 sky130_as_sc_hs__and2_2 _40974_ (.A(_10229_),
    .B(_10230_),
    .Y(_10231_));
 sky130_as_sc_hs__or2_2 _40976_ (.A(_10214_),
    .B(_10231_),
    .Y(_10233_));
 sky130_as_sc_hs__and2_2 _40977_ (.A(_10232_),
    .B(_10233_),
    .Y(_10234_));
 sky130_as_sc_hs__or2_2 _40980_ (.A(_10234_),
    .B(_10235_),
    .Y(_10237_));
 sky130_as_sc_hs__and2_2 _40981_ (.A(_10236_),
    .B(_10237_),
    .Y(_10238_));
 sky130_as_sc_hs__and2_2 _40984_ (.A(net480),
    .B(net128),
    .Y(_10241_));
 sky130_as_sc_hs__or2_2 _40986_ (.A(_10000_),
    .B(_10241_),
    .Y(_10243_));
 sky130_as_sc_hs__or2_2 _40988_ (.A(_10026_),
    .B(_10244_),
    .Y(_10245_));
 sky130_as_sc_hs__and2_2 _40990_ (.A(_10245_),
    .B(_10246_),
    .Y(_10247_));
 sky130_as_sc_hs__and2_2 _40991_ (.A(net476),
    .B(net421),
    .Y(_10248_));
 sky130_as_sc_hs__or2_2 _40993_ (.A(_10247_),
    .B(_10248_),
    .Y(_10250_));
 sky130_as_sc_hs__and2_2 _40994_ (.A(_10249_),
    .B(_10250_),
    .Y(_10251_));
 sky130_as_sc_hs__or2_2 _40996_ (.A(_10240_),
    .B(_10251_),
    .Y(_10253_));
 sky130_as_sc_hs__and2_2 _40997_ (.A(_10252_),
    .B(_10253_),
    .Y(_10254_));
 sky130_as_sc_hs__or2_2 _40999_ (.A(_10239_),
    .B(_10254_),
    .Y(_10256_));
 sky130_as_sc_hs__and2_2 _41000_ (.A(_10255_),
    .B(_10256_),
    .Y(_10257_));
 sky130_as_sc_hs__or2_2 _41002_ (.A(_10238_),
    .B(_10257_),
    .Y(_10259_));
 sky130_as_sc_hs__and2_2 _41003_ (.A(_10258_),
    .B(_10259_),
    .Y(_10260_));
 sky130_as_sc_hs__or2_2 _41006_ (.A(_10260_),
    .B(_10261_),
    .Y(_10263_));
 sky130_as_sc_hs__and2_2 _41007_ (.A(_10262_),
    .B(_10263_),
    .Y(_10264_));
 sky130_as_sc_hs__or2_2 _41010_ (.A(_10264_),
    .B(_10265_),
    .Y(_10267_));
 sky130_as_sc_hs__and2_2 _41011_ (.A(_10266_),
    .B(_10267_),
    .Y(_10268_));
 sky130_as_sc_hs__or2_2 _41014_ (.A(_10268_),
    .B(_10269_),
    .Y(_10271_));
 sky130_as_sc_hs__and2_2 _41015_ (.A(_10270_),
    .B(_10271_),
    .Y(_10272_));
 sky130_as_sc_hs__or2_2 _41016_ (.A(_10053_),
    .B(_10272_),
    .Y(_10273_));
 sky130_as_sc_hs__or2_2 _41020_ (.A(_10140_),
    .B(_10275_),
    .Y(_10277_));
 sky130_as_sc_hs__and2_2 _41021_ (.A(_10276_),
    .B(_10277_),
    .Y(_10278_));
 sky130_as_sc_hs__nor2_2 _41022_ (.A(_05500_),
    .B(_10066_),
    .Y(_10279_));
 sky130_as_sc_hs__nand3_2 _41023_ (.A(_09620_),
    .B(_10067_),
    .C(_10279_),
    .Y(_10280_));
 sky130_as_sc_hs__and2_2 _41025_ (.A(_08636_),
    .B(_10281_),
    .Y(_10282_));
 sky130_as_sc_hs__or2_2 _41027_ (.A(_10278_),
    .B(_10282_),
    .Y(_10284_));
 sky130_as_sc_hs__nand3_2 _41028_ (.A(net141),
    .B(_10283_),
    .C(_10284_),
    .Y(_10285_));
 sky130_as_sc_hs__or2_2 _41029_ (.A(_05425_),
    .B(_05505_),
    .Y(_10286_));
 sky130_as_sc_hs__or2_2 _41031_ (.A(_05429_),
    .B(_10286_),
    .Y(_10288_));
 sky130_as_sc_hs__nand3_2 _41032_ (.A(net139),
    .B(_10287_),
    .C(_10288_),
    .Y(_10289_));
 sky130_as_sc_hs__and2_2 _41033_ (.A(_05684_),
    .B(_10079_),
    .Y(_10290_));
 sky130_as_sc_hs__or2_2 _41034_ (.A(_05676_),
    .B(_10290_),
    .Y(_10291_));
 sky130_as_sc_hs__or2_2 _41038_ (.A(_05676_),
    .B(_05879_),
    .Y(_10295_));
 sky130_as_sc_hs__nand3_2 _41041_ (.A(net118),
    .B(_10294_),
    .C(_10297_),
    .Y(_10298_));
 sky130_as_sc_hs__or2_2 _41042_ (.A(_05935_),
    .B(_08382_),
    .Y(_10299_));
 sky130_as_sc_hs__nand3_2 _41044_ (.A(_05929_),
    .B(_10299_),
    .C(_10300_),
    .Y(_10301_));
 sky130_as_sc_hs__or2_2 _41045_ (.A(_05929_),
    .B(_05963_),
    .Y(_10302_));
 sky130_as_sc_hs__and2_2 _41046_ (.A(_10301_),
    .B(_10302_),
    .Y(_10303_));
 sky130_as_sc_hs__and2_2 _41050_ (.A(net140),
    .B(_10306_),
    .Y(_10307_));
 sky130_as_sc_hs__or2_2 _41051_ (.A(\tholin_riscv.div_res[14] ),
    .B(_10101_),
    .Y(_10308_));
 sky130_as_sc_hs__and2_2 _41052_ (.A(net414),
    .B(_10308_),
    .Y(_10309_));
 sky130_as_sc_hs__or2_2 _41053_ (.A(\tholin_riscv.div_res[15] ),
    .B(_10309_),
    .Y(_10310_));
 sky130_as_sc_hs__nand3_2 _41055_ (.A(net110),
    .B(_10310_),
    .C(_10311_),
    .Y(_10312_));
 sky130_as_sc_hs__or2_2 _41056_ (.A(\tholin_riscv.div_shifter[46] ),
    .B(_10096_),
    .Y(_10313_));
 sky130_as_sc_hs__and2_2 _41057_ (.A(_21655_),
    .B(_10313_),
    .Y(_10314_));
 sky130_as_sc_hs__or2_2 _41058_ (.A(\tholin_riscv.div_shifter[47] ),
    .B(_10314_),
    .Y(_10315_));
 sky130_as_sc_hs__nand3_2 _41060_ (.A(net107),
    .B(_10315_),
    .C(_10316_),
    .Y(_10317_));
 sky130_as_sc_hs__nor2_2 _41064_ (.A(_05674_),
    .B(_06161_),
    .Y(_10321_));
 sky130_as_sc_hs__nand3_2 _41067_ (.A(net412),
    .B(_10322_),
    .C(_10323_),
    .Y(_10324_));
 sky130_as_sc_hs__nor2_2 _41068_ (.A(_10321_),
    .B(_10324_),
    .Y(_10325_));
 sky130_as_sc_hs__and2_2 _41069_ (.A(_10320_),
    .B(_10325_),
    .Y(_10326_));
 sky130_as_sc_hs__nand3_2 _41070_ (.A(_10312_),
    .B(_10317_),
    .C(_10326_),
    .Y(_10327_));
 sky130_as_sc_hs__nor2_2 _41071_ (.A(_10307_),
    .B(_10327_),
    .Y(_10328_));
 sky130_as_sc_hs__and2_2 _41072_ (.A(_10304_),
    .B(_10328_),
    .Y(_10329_));
 sky130_as_sc_hs__and2_2 _41073_ (.A(_10298_),
    .B(_10329_),
    .Y(_10330_));
 sky130_as_sc_hs__nand3_2 _41074_ (.A(_10285_),
    .B(_10289_),
    .C(_10330_),
    .Y(_10331_));
 sky130_as_sc_hs__and2_2 _41075_ (.A(\tholin_riscv.PC[15] ),
    .B(_10120_),
    .Y(_10332_));
 sky130_as_sc_hs__nor2_2 _41076_ (.A(\tholin_riscv.PC[15] ),
    .B(_10120_),
    .Y(_10333_));
 sky130_as_sc_hs__or2_2 _41077_ (.A(_10332_),
    .B(_10333_),
    .Y(_10334_));
 sky130_as_sc_hs__or2_2 _41083_ (.A(\tholin_riscv.PC[15] ),
    .B(net373),
    .Y(_10340_));
 sky130_as_sc_hs__or2_2 _41086_ (.A(_10338_),
    .B(_10341_),
    .Y(_10343_));
 sky130_as_sc_hs__nand3_2 _41087_ (.A(net117),
    .B(_10342_),
    .C(_10343_),
    .Y(_10344_));
 sky130_as_sc_hs__nand3_2 _41088_ (.A(_10335_),
    .B(_10336_),
    .C(_10344_),
    .Y(_10345_));
 sky130_as_sc_hs__nand3_2 _41090_ (.A(_21546_),
    .B(_10331_),
    .C(_10346_),
    .Y(_10347_));
 sky130_as_sc_hs__and2_2 _41096_ (.A(_08426_),
    .B(_10351_),
    .Y(_10352_));
 sky130_as_sc_hs__and2_2 _41097_ (.A(net360),
    .B(net371),
    .Y(_10353_));
 sky130_as_sc_hs__or2_2 _41098_ (.A(_10352_),
    .B(_10353_),
    .Y(_10354_));
 sky130_as_sc_hs__and2_2 _41100_ (.A(_10058_),
    .B(_10275_),
    .Y(_10356_));
 sky130_as_sc_hs__and2_2 _41101_ (.A(_10061_),
    .B(_10356_),
    .Y(_10357_));
 sky130_as_sc_hs__inv_2 _41102_ (.Y(_10358_),
    .A(_10357_));
 sky130_as_sc_hs__and2_2 _41103_ (.A(_09614_),
    .B(_10357_),
    .Y(_10359_));
 sky130_as_sc_hs__inv_2 _41104_ (.Y(_10360_),
    .A(_10359_));
 sky130_as_sc_hs__nand3_2 _41105_ (.A(_05123_),
    .B(_08623_),
    .C(_10359_),
    .Y(_10361_));
 sky130_as_sc_hs__or2_2 _41106_ (.A(_08629_),
    .B(_10360_),
    .Y(_10362_));
 sky130_as_sc_hs__or2_2 _41107_ (.A(_09613_),
    .B(_10358_),
    .Y(_10363_));
 sky130_as_sc_hs__nand3_2 _41108_ (.A(_09838_),
    .B(_10059_),
    .C(_10356_),
    .Y(_10364_));
 sky130_as_sc_hs__and2_2 _41111_ (.A(_10364_),
    .B(_10366_),
    .Y(_10367_));
 sky130_as_sc_hs__and2_2 _41112_ (.A(_10363_),
    .B(_10367_),
    .Y(_10368_));
 sky130_as_sc_hs__nand3_2 _41113_ (.A(_10361_),
    .B(_10362_),
    .C(_10368_),
    .Y(_10369_));
 sky130_as_sc_hs__and2_2 _41114_ (.A(net480),
    .B(_02550_),
    .Y(_10370_));
 sky130_as_sc_hs__and2_2 _41115_ (.A(net478),
    .B(net433),
    .Y(_10371_));
 sky130_as_sc_hs__or2_2 _41116_ (.A(_10370_),
    .B(_10371_),
    .Y(_10372_));
 sky130_as_sc_hs__and2_2 _41118_ (.A(_10372_),
    .B(_10373_),
    .Y(_10374_));
 sky130_as_sc_hs__and2_2 _41119_ (.A(net457),
    .B(net83),
    .Y(_10375_));
 sky130_as_sc_hs__or2_2 _41121_ (.A(_10374_),
    .B(_10375_),
    .Y(_10377_));
 sky130_as_sc_hs__and2_2 _41122_ (.A(_10376_),
    .B(_10377_),
    .Y(_10378_));
 sky130_as_sc_hs__or2_2 _41125_ (.A(_10378_),
    .B(_10379_),
    .Y(_10381_));
 sky130_as_sc_hs__and2_2 _41126_ (.A(_10380_),
    .B(_10381_),
    .Y(_10382_));
 sky130_as_sc_hs__and2_2 _41127_ (.A(net466),
    .B(net427),
    .Y(_10383_));
 sky130_as_sc_hs__and2_2 _41128_ (.A(net120),
    .B(net468),
    .Y(_10384_));
 sky130_as_sc_hs__or2_2 _41129_ (.A(_10383_),
    .B(_10384_),
    .Y(_10385_));
 sky130_as_sc_hs__and2_2 _41131_ (.A(_10385_),
    .B(_10386_),
    .Y(_10387_));
 sky130_as_sc_hs__and2_2 _41132_ (.A(net122),
    .B(net471),
    .Y(_10388_));
 sky130_as_sc_hs__or2_2 _41134_ (.A(_10387_),
    .B(_10388_),
    .Y(_10390_));
 sky130_as_sc_hs__and2_2 _41135_ (.A(_10389_),
    .B(_10390_),
    .Y(_10391_));
 sky130_as_sc_hs__or2_2 _41137_ (.A(_10382_),
    .B(_10391_),
    .Y(_10393_));
 sky130_as_sc_hs__and2_2 _41138_ (.A(_10392_),
    .B(_10393_),
    .Y(_10394_));
 sky130_as_sc_hs__or2_2 _41141_ (.A(_10394_),
    .B(_10395_),
    .Y(_10397_));
 sky130_as_sc_hs__and2_2 _41142_ (.A(_10396_),
    .B(_10397_),
    .Y(_10398_));
 sky130_as_sc_hs__and2_2 _41145_ (.A(net465),
    .B(net423),
    .Y(_10401_));
 sky130_as_sc_hs__and2_2 _41146_ (.A(net463),
    .B(net419),
    .Y(_10402_));
 sky130_as_sc_hs__or2_2 _41147_ (.A(_10401_),
    .B(_10402_),
    .Y(_10403_));
 sky130_as_sc_hs__and2_2 _41149_ (.A(_10403_),
    .B(_10404_),
    .Y(_10405_));
 sky130_as_sc_hs__and2_2 _41150_ (.A(net460),
    .B(net74),
    .Y(_10406_));
 sky130_as_sc_hs__or2_2 _41152_ (.A(_10405_),
    .B(_10406_),
    .Y(_10408_));
 sky130_as_sc_hs__and2_2 _41153_ (.A(_10407_),
    .B(_10408_),
    .Y(_10409_));
 sky130_as_sc_hs__or2_2 _41155_ (.A(_10400_),
    .B(_10409_),
    .Y(_10411_));
 sky130_as_sc_hs__and2_2 _41156_ (.A(_10410_),
    .B(_10411_),
    .Y(_10412_));
 sky130_as_sc_hs__or2_2 _41158_ (.A(_10399_),
    .B(_10412_),
    .Y(_10414_));
 sky130_as_sc_hs__and2_2 _41159_ (.A(_10413_),
    .B(_10414_),
    .Y(_10415_));
 sky130_as_sc_hs__or2_2 _41161_ (.A(_10398_),
    .B(_10415_),
    .Y(_10417_));
 sky130_as_sc_hs__and2_2 _41162_ (.A(_10416_),
    .B(_10417_),
    .Y(_10418_));
 sky130_as_sc_hs__or2_2 _41165_ (.A(_10418_),
    .B(_10419_),
    .Y(_10421_));
 sky130_as_sc_hs__and2_2 _41166_ (.A(_10420_),
    .B(_10421_),
    .Y(_10422_));
 sky130_as_sc_hs__and2_2 _41168_ (.A(net472),
    .B(net425),
    .Y(_10424_));
 sky130_as_sc_hs__or2_2 _41171_ (.A(_10424_),
    .B(_10425_),
    .Y(_10427_));
 sky130_as_sc_hs__and2_2 _41172_ (.A(_10426_),
    .B(_10427_),
    .Y(_10428_));
 sky130_as_sc_hs__or2_2 _41174_ (.A(_10423_),
    .B(_10428_),
    .Y(_10430_));
 sky130_as_sc_hs__and2_2 _41175_ (.A(_10429_),
    .B(_10430_),
    .Y(_10431_));
 sky130_as_sc_hs__or2_2 _41177_ (.A(_10422_),
    .B(_10431_),
    .Y(_10433_));
 sky130_as_sc_hs__and2_2 _41178_ (.A(_10432_),
    .B(_10433_),
    .Y(_10434_));
 sky130_as_sc_hs__or2_2 _41181_ (.A(_10434_),
    .B(_10435_),
    .Y(_10437_));
 sky130_as_sc_hs__and2_2 _41182_ (.A(_10436_),
    .B(_10437_),
    .Y(_10438_));
 sky130_as_sc_hs__and2_2 _41184_ (.A(net474),
    .B(net434),
    .Y(_10440_));
 sky130_as_sc_hs__and2_2 _41185_ (.A(net436),
    .B(net429),
    .Y(_10441_));
 sky130_as_sc_hs__and2_2 _41186_ (.A(net440),
    .B(net431),
    .Y(_10442_));
 sky130_as_sc_hs__and2_2 _41187_ (.A(_10441_),
    .B(_10442_),
    .Y(_10443_));
 sky130_as_sc_hs__or2_2 _41188_ (.A(_10441_),
    .B(_10442_),
    .Y(_10444_));
 sky130_as_sc_hs__nor2b_2 _41189_ (.A(_10443_),
    .Y(_10445_),
    .B(_10444_));
 sky130_as_sc_hs__or2_2 _41191_ (.A(_10440_),
    .B(_10445_),
    .Y(_10447_));
 sky130_as_sc_hs__and2_2 _41192_ (.A(_10446_),
    .B(_10447_),
    .Y(_10448_));
 sky130_as_sc_hs__or2_2 _41194_ (.A(_10439_),
    .B(_10448_),
    .Y(_10450_));
 sky130_as_sc_hs__or2_2 _41196_ (.A(_10223_),
    .B(_10451_),
    .Y(_10452_));
 sky130_as_sc_hs__and2_2 _41198_ (.A(_10452_),
    .B(_10453_),
    .Y(_10454_));
 sky130_as_sc_hs__or2_2 _41200_ (.A(_10438_),
    .B(_10454_),
    .Y(_10456_));
 sky130_as_sc_hs__and2_2 _41201_ (.A(_10455_),
    .B(_10456_),
    .Y(_10457_));
 sky130_as_sc_hs__or2_2 _41204_ (.A(_10457_),
    .B(_10458_),
    .Y(_10460_));
 sky130_as_sc_hs__and2_2 _41205_ (.A(_10459_),
    .B(_10460_),
    .Y(_10461_));
 sky130_as_sc_hs__and2_2 _41208_ (.A(net476),
    .B(net128),
    .Y(_10464_));
 sky130_as_sc_hs__or2_2 _41210_ (.A(_10220_),
    .B(_10464_),
    .Y(_10466_));
 sky130_as_sc_hs__or2_2 _41212_ (.A(_10242_),
    .B(_10467_),
    .Y(_10468_));
 sky130_as_sc_hs__and2_2 _41214_ (.A(_10468_),
    .B(_10469_),
    .Y(_10470_));
 sky130_as_sc_hs__and2_2 _41215_ (.A(net438),
    .B(net421),
    .Y(_10471_));
 sky130_as_sc_hs__or2_2 _41217_ (.A(_10470_),
    .B(_10471_),
    .Y(_10473_));
 sky130_as_sc_hs__and2_2 _41218_ (.A(_10472_),
    .B(_10473_),
    .Y(_10474_));
 sky130_as_sc_hs__or2_2 _41220_ (.A(_10463_),
    .B(_10474_),
    .Y(_10476_));
 sky130_as_sc_hs__and2_2 _41221_ (.A(_10475_),
    .B(_10476_),
    .Y(_10477_));
 sky130_as_sc_hs__or2_2 _41223_ (.A(_10462_),
    .B(_10477_),
    .Y(_10479_));
 sky130_as_sc_hs__and2_2 _41224_ (.A(_10478_),
    .B(_10479_),
    .Y(_10480_));
 sky130_as_sc_hs__or2_2 _41226_ (.A(_10461_),
    .B(_10480_),
    .Y(_10482_));
 sky130_as_sc_hs__and2_2 _41227_ (.A(_10481_),
    .B(_10482_),
    .Y(_10483_));
 sky130_as_sc_hs__or2_2 _41230_ (.A(_10483_),
    .B(_10484_),
    .Y(_10486_));
 sky130_as_sc_hs__and2_2 _41231_ (.A(_10485_),
    .B(_10486_),
    .Y(_10487_));
 sky130_as_sc_hs__or2_2 _41234_ (.A(_10487_),
    .B(_10488_),
    .Y(_10490_));
 sky130_as_sc_hs__and2_2 _41235_ (.A(_10489_),
    .B(_10490_),
    .Y(_10491_));
 sky130_as_sc_hs__or2_2 _41238_ (.A(_10491_),
    .B(_10492_),
    .Y(_10494_));
 sky130_as_sc_hs__or2_2 _41240_ (.A(_10270_),
    .B(_10495_),
    .Y(_10496_));
 sky130_as_sc_hs__and2_2 _41242_ (.A(_10496_),
    .B(_10497_),
    .Y(_10498_));
 sky130_as_sc_hs__or2_2 _41244_ (.A(_10369_),
    .B(_10498_),
    .Y(_10500_));
 sky130_as_sc_hs__nand3_2 _41246_ (.A(_08635_),
    .B(_10276_),
    .C(_10277_),
    .Y(_10502_));
 sky130_as_sc_hs__nor2_2 _41247_ (.A(_10280_),
    .B(_10502_),
    .Y(_10503_));
 sky130_as_sc_hs__or2_2 _41248_ (.A(_05505_),
    .B(_10503_),
    .Y(_10504_));
 sky130_as_sc_hs__or2_2 _41250_ (.A(_10501_),
    .B(_10504_),
    .Y(_10506_));
 sky130_as_sc_hs__nand3_2 _41251_ (.A(net141),
    .B(_10505_),
    .C(_10506_),
    .Y(_10507_));
 sky130_as_sc_hs__or2_2 _41252_ (.A(_05430_),
    .B(_05505_),
    .Y(_10508_));
 sky130_as_sc_hs__or2_2 _41253_ (.A(_05377_),
    .B(_10508_),
    .Y(_10509_));
 sky130_as_sc_hs__nand3_2 _41255_ (.A(net138),
    .B(_10509_),
    .C(_10510_),
    .Y(_10511_));
 sky130_as_sc_hs__or2_2 _41258_ (.A(_05666_),
    .B(_10512_),
    .Y(_10514_));
 sky130_as_sc_hs__and2_2 _41259_ (.A(_10513_),
    .B(_10514_),
    .Y(_10515_));
 sky130_as_sc_hs__or2_2 _41261_ (.A(_05666_),
    .B(_05881_),
    .Y(_10517_));
 sky130_as_sc_hs__nand3_2 _41264_ (.A(net119),
    .B(_10516_),
    .C(_10519_),
    .Y(_10520_));
 sky130_as_sc_hs__and2_2 _41266_ (.A(net140),
    .B(_10303_),
    .Y(_10522_));
 sky130_as_sc_hs__or2_2 _41267_ (.A(\tholin_riscv.div_shifter[47] ),
    .B(_10313_),
    .Y(_10523_));
 sky130_as_sc_hs__and2_2 _41268_ (.A(_21655_),
    .B(_10523_),
    .Y(_10524_));
 sky130_as_sc_hs__or2_2 _41269_ (.A(\tholin_riscv.div_shifter[48] ),
    .B(_10524_),
    .Y(_10525_));
 sky130_as_sc_hs__nand3_2 _41271_ (.A(net107),
    .B(_10525_),
    .C(_10526_),
    .Y(_10527_));
 sky130_as_sc_hs__or2_2 _41272_ (.A(\tholin_riscv.div_res[15] ),
    .B(_10308_),
    .Y(_10528_));
 sky130_as_sc_hs__and2_2 _41273_ (.A(net414),
    .B(_10528_),
    .Y(_10529_));
 sky130_as_sc_hs__or2_2 _41274_ (.A(\tholin_riscv.div_res[16] ),
    .B(_10529_),
    .Y(_10530_));
 sky130_as_sc_hs__nand3_2 _41276_ (.A(net110),
    .B(_10530_),
    .C(_10531_),
    .Y(_10532_));
 sky130_as_sc_hs__nor2_2 _41280_ (.A(_05664_),
    .B(_06161_),
    .Y(_10536_));
 sky130_as_sc_hs__nand3_2 _41283_ (.A(net412),
    .B(_10537_),
    .C(_10538_),
    .Y(_10539_));
 sky130_as_sc_hs__nor2_2 _41284_ (.A(_10536_),
    .B(_10539_),
    .Y(_10540_));
 sky130_as_sc_hs__and2_2 _41285_ (.A(_10535_),
    .B(_10540_),
    .Y(_10541_));
 sky130_as_sc_hs__nand3_2 _41286_ (.A(_10527_),
    .B(_10532_),
    .C(_10541_),
    .Y(_10542_));
 sky130_as_sc_hs__nor2_2 _41287_ (.A(_10522_),
    .B(_10542_),
    .Y(_10543_));
 sky130_as_sc_hs__and2_2 _41288_ (.A(_10521_),
    .B(_10543_),
    .Y(_10544_));
 sky130_as_sc_hs__and2_2 _41289_ (.A(_10520_),
    .B(_10544_),
    .Y(_10545_));
 sky130_as_sc_hs__nand3_2 _41290_ (.A(_10507_),
    .B(_10511_),
    .C(_10545_),
    .Y(_10546_));
 sky130_as_sc_hs__and2_2 _41291_ (.A(\tholin_riscv.PC[16] ),
    .B(_10332_),
    .Y(_10547_));
 sky130_as_sc_hs__nor2_2 _41292_ (.A(\tholin_riscv.PC[16] ),
    .B(_10332_),
    .Y(_10548_));
 sky130_as_sc_hs__or2_2 _41293_ (.A(_10547_),
    .B(_10548_),
    .Y(_10549_));
 sky130_as_sc_hs__or2_2 _41299_ (.A(\tholin_riscv.PC[16] ),
    .B(net353),
    .Y(_10555_));
 sky130_as_sc_hs__or2_2 _41301_ (.A(_10553_),
    .B(_10556_),
    .Y(_10557_));
 sky130_as_sc_hs__nand3_2 _41303_ (.A(net117),
    .B(_10557_),
    .C(_10558_),
    .Y(_10559_));
 sky130_as_sc_hs__nand3_2 _41304_ (.A(_10550_),
    .B(_10551_),
    .C(_10559_),
    .Y(_10560_));
 sky130_as_sc_hs__nand3_2 _41306_ (.A(_21546_),
    .B(_10546_),
    .C(_10561_),
    .Y(_10562_));
 sky130_as_sc_hs__and2_2 _41311_ (.A(net347),
    .B(net371),
    .Y(_10566_));
 sky130_as_sc_hs__or2_2 _41312_ (.A(_10352_),
    .B(_10566_),
    .Y(_10567_));
 sky130_as_sc_hs__and2_2 _41314_ (.A(_10496_),
    .B(_10499_),
    .Y(_10569_));
 sky130_as_sc_hs__and2_2 _41315_ (.A(net476),
    .B(net418),
    .Y(_10570_));
 sky130_as_sc_hs__and2_2 _41316_ (.A(net474),
    .B(net433),
    .Y(_10571_));
 sky130_as_sc_hs__or2_2 _41317_ (.A(_10570_),
    .B(_10571_),
    .Y(_10572_));
 sky130_as_sc_hs__and2_2 _41319_ (.A(_10572_),
    .B(_10573_),
    .Y(_10574_));
 sky130_as_sc_hs__and2_2 _41320_ (.A(net457),
    .B(net431),
    .Y(_10575_));
 sky130_as_sc_hs__or2_2 _41322_ (.A(_10574_),
    .B(_10575_),
    .Y(_10577_));
 sky130_as_sc_hs__and2_2 _41323_ (.A(_10576_),
    .B(_10577_),
    .Y(_10578_));
 sky130_as_sc_hs__or2_2 _41326_ (.A(_10578_),
    .B(_10579_),
    .Y(_10581_));
 sky130_as_sc_hs__and2_2 _41327_ (.A(_10580_),
    .B(_10581_),
    .Y(_10582_));
 sky130_as_sc_hs__and2_2 _41328_ (.A(net120),
    .B(net466),
    .Y(_10583_));
 sky130_as_sc_hs__and2_2 _41329_ (.A(net122),
    .B(net468),
    .Y(_10584_));
 sky130_as_sc_hs__or2_2 _41330_ (.A(_10583_),
    .B(_10584_),
    .Y(_10585_));
 sky130_as_sc_hs__and2_2 _41332_ (.A(_10585_),
    .B(_10586_),
    .Y(_10587_));
 sky130_as_sc_hs__and2_2 _41333_ (.A(net471),
    .B(net423),
    .Y(_10588_));
 sky130_as_sc_hs__or2_2 _41335_ (.A(_10587_),
    .B(_10588_),
    .Y(_10590_));
 sky130_as_sc_hs__and2_2 _41336_ (.A(_10589_),
    .B(_10590_),
    .Y(_10591_));
 sky130_as_sc_hs__or2_2 _41338_ (.A(_10582_),
    .B(_10591_),
    .Y(_10593_));
 sky130_as_sc_hs__and2_2 _41339_ (.A(_10592_),
    .B(_10593_),
    .Y(_10594_));
 sky130_as_sc_hs__or2_2 _41342_ (.A(_10594_),
    .B(_10595_),
    .Y(_10597_));
 sky130_as_sc_hs__and2_2 _41343_ (.A(_10596_),
    .B(_10597_),
    .Y(_10598_));
 sky130_as_sc_hs__and2_2 _41346_ (.A(net464),
    .B(net420),
    .Y(_10601_));
 sky130_as_sc_hs__or2_2 _41348_ (.A(_10601_),
    .B(_10602_),
    .Y(_10603_));
 sky130_as_sc_hs__or2_2 _41352_ (.A(_10600_),
    .B(_10605_),
    .Y(_10607_));
 sky130_as_sc_hs__and2_2 _41353_ (.A(_10606_),
    .B(_10607_),
    .Y(_10608_));
 sky130_as_sc_hs__or2_2 _41355_ (.A(_10599_),
    .B(_10608_),
    .Y(_10610_));
 sky130_as_sc_hs__and2_2 _41356_ (.A(_10609_),
    .B(_10610_),
    .Y(_10611_));
 sky130_as_sc_hs__or2_2 _41358_ (.A(_10598_),
    .B(_10611_),
    .Y(_10613_));
 sky130_as_sc_hs__and2_2 _41359_ (.A(_10612_),
    .B(_10613_),
    .Y(_10614_));
 sky130_as_sc_hs__or2_2 _41362_ (.A(_10614_),
    .B(_10615_),
    .Y(_10617_));
 sky130_as_sc_hs__and2_2 _41363_ (.A(_10616_),
    .B(_10617_),
    .Y(_10618_));
 sky130_as_sc_hs__and2_2 _41364_ (.A(net478),
    .B(net425),
    .Y(_10619_));
 sky130_as_sc_hs__or2_2 _41367_ (.A(_10619_),
    .B(_10620_),
    .Y(_10622_));
 sky130_as_sc_hs__and2_2 _41368_ (.A(_10621_),
    .B(_10622_),
    .Y(_10623_));
 sky130_as_sc_hs__or2_2 _41370_ (.A(_10618_),
    .B(_10623_),
    .Y(_10625_));
 sky130_as_sc_hs__and2_2 _41371_ (.A(_10624_),
    .B(_10625_),
    .Y(_10626_));
 sky130_as_sc_hs__or2_2 _41374_ (.A(_10626_),
    .B(_10627_),
    .Y(_10629_));
 sky130_as_sc_hs__and2_2 _41375_ (.A(_10628_),
    .B(_10629_),
    .Y(_10630_));
 sky130_as_sc_hs__and2_2 _41377_ (.A(net434),
    .B(net83),
    .Y(_10632_));
 sky130_as_sc_hs__and2_2 _41378_ (.A(net436),
    .B(net428),
    .Y(_10633_));
 sky130_as_sc_hs__and2_2 _41379_ (.A(net440),
    .B(net430),
    .Y(_10634_));
 sky130_as_sc_hs__and2_2 _41380_ (.A(_10633_),
    .B(_10634_),
    .Y(_10635_));
 sky130_as_sc_hs__or2_2 _41381_ (.A(_10633_),
    .B(_10634_),
    .Y(_10636_));
 sky130_as_sc_hs__nor2b_2 _41382_ (.A(_10635_),
    .Y(_10637_),
    .B(_10636_));
 sky130_as_sc_hs__or2_2 _41384_ (.A(_10632_),
    .B(_10637_),
    .Y(_10639_));
 sky130_as_sc_hs__and2_2 _41385_ (.A(_10638_),
    .B(_10639_),
    .Y(_10640_));
 sky130_as_sc_hs__or2_2 _41387_ (.A(_10631_),
    .B(_10640_),
    .Y(_10642_));
 sky130_as_sc_hs__or2_2 _41389_ (.A(_10446_),
    .B(_10643_),
    .Y(_10644_));
 sky130_as_sc_hs__and2_2 _41391_ (.A(_10644_),
    .B(_10645_),
    .Y(_10646_));
 sky130_as_sc_hs__or2_2 _41393_ (.A(_10630_),
    .B(_10646_),
    .Y(_10648_));
 sky130_as_sc_hs__and2_2 _41394_ (.A(_10647_),
    .B(_10648_),
    .Y(_10649_));
 sky130_as_sc_hs__or2_2 _41397_ (.A(_10649_),
    .B(_10650_),
    .Y(_10652_));
 sky130_as_sc_hs__and2_2 _41398_ (.A(_10651_),
    .B(_10652_),
    .Y(_10653_));
 sky130_as_sc_hs__and2_2 _41401_ (.A(net439),
    .B(net128),
    .Y(_10656_));
 sky130_as_sc_hs__or2_2 _41403_ (.A(_10443_),
    .B(_10656_),
    .Y(_10658_));
 sky130_as_sc_hs__or2_2 _41405_ (.A(_10465_),
    .B(_10659_),
    .Y(_10660_));
 sky130_as_sc_hs__and2_2 _41407_ (.A(_10660_),
    .B(_10661_),
    .Y(_10662_));
 sky130_as_sc_hs__and2_2 _41408_ (.A(net472),
    .B(net421),
    .Y(_10663_));
 sky130_as_sc_hs__or2_2 _41410_ (.A(_10662_),
    .B(_10663_),
    .Y(_10665_));
 sky130_as_sc_hs__and2_2 _41411_ (.A(_10664_),
    .B(_10665_),
    .Y(_10666_));
 sky130_as_sc_hs__or2_2 _41413_ (.A(_10655_),
    .B(_10666_),
    .Y(_10668_));
 sky130_as_sc_hs__and2_2 _41414_ (.A(_10667_),
    .B(_10668_),
    .Y(_10669_));
 sky130_as_sc_hs__or2_2 _41416_ (.A(_10654_),
    .B(_10669_),
    .Y(_10671_));
 sky130_as_sc_hs__and2_2 _41417_ (.A(_10670_),
    .B(_10671_),
    .Y(_10672_));
 sky130_as_sc_hs__or2_2 _41419_ (.A(_10653_),
    .B(_10672_),
    .Y(_10674_));
 sky130_as_sc_hs__and2_2 _41420_ (.A(_10673_),
    .B(_10674_),
    .Y(_10675_));
 sky130_as_sc_hs__or2_2 _41423_ (.A(_10675_),
    .B(_10676_),
    .Y(_10678_));
 sky130_as_sc_hs__and2_2 _41424_ (.A(_10677_),
    .B(_10678_),
    .Y(_10679_));
 sky130_as_sc_hs__or2_2 _41427_ (.A(_10679_),
    .B(_10680_),
    .Y(_10682_));
 sky130_as_sc_hs__and2_2 _41428_ (.A(_10681_),
    .B(_10682_),
    .Y(_10683_));
 sky130_as_sc_hs__or2_2 _41431_ (.A(_10683_),
    .B(_10684_),
    .Y(_10686_));
 sky130_as_sc_hs__and2_2 _41432_ (.A(_10685_),
    .B(_10686_),
    .Y(_10687_));
 sky130_as_sc_hs__nor2_2 _41433_ (.A(_10493_),
    .B(_10687_),
    .Y(_10688_));
 sky130_as_sc_hs__and2_2 _41434_ (.A(_10493_),
    .B(_10687_),
    .Y(_10689_));
 sky130_as_sc_hs__or2_2 _41435_ (.A(_10688_),
    .B(_10689_),
    .Y(_10690_));
 sky130_as_sc_hs__or2_2 _41437_ (.A(_10569_),
    .B(_10690_),
    .Y(_10692_));
 sky130_as_sc_hs__and2_2 _41438_ (.A(_10691_),
    .B(_10692_),
    .Y(_10693_));
 sky130_as_sc_hs__or2_2 _41441_ (.A(_10693_),
    .B(_10694_),
    .Y(_10696_));
 sky130_as_sc_hs__nand3_2 _41442_ (.A(net141),
    .B(_10695_),
    .C(_10696_),
    .Y(_10697_));
 sky130_as_sc_hs__or2_2 _41444_ (.A(_05381_),
    .B(_10698_),
    .Y(_10699_));
 sky130_as_sc_hs__nand3_2 _41446_ (.A(net139),
    .B(_10699_),
    .C(_10700_),
    .Y(_10701_));
 sky130_as_sc_hs__or2_2 _41449_ (.A(_05658_),
    .B(_10703_),
    .Y(_10704_));
 sky130_as_sc_hs__and2_2 _41451_ (.A(_10704_),
    .B(_10705_),
    .Y(_10706_));
 sky130_as_sc_hs__or2_2 _41453_ (.A(_05658_),
    .B(_05884_),
    .Y(_10708_));
 sky130_as_sc_hs__nand3_2 _41456_ (.A(net119),
    .B(_10707_),
    .C(_10710_),
    .Y(_10711_));
 sky130_as_sc_hs__and2_2 _41458_ (.A(net140),
    .B(_10091_),
    .Y(_10713_));
 sky130_as_sc_hs__or2_2 _41459_ (.A(\tholin_riscv.div_res[16] ),
    .B(_10528_),
    .Y(_10714_));
 sky130_as_sc_hs__and2_2 _41460_ (.A(net414),
    .B(_10714_),
    .Y(_10715_));
 sky130_as_sc_hs__or2_2 _41461_ (.A(\tholin_riscv.div_res[17] ),
    .B(_10715_),
    .Y(_10716_));
 sky130_as_sc_hs__nand3_2 _41463_ (.A(net110),
    .B(_10716_),
    .C(_10717_),
    .Y(_10718_));
 sky130_as_sc_hs__or2_2 _41464_ (.A(\tholin_riscv.div_shifter[48] ),
    .B(_10523_),
    .Y(_10719_));
 sky130_as_sc_hs__and2_2 _41465_ (.A(_21655_),
    .B(_10719_),
    .Y(_10720_));
 sky130_as_sc_hs__or2_2 _41466_ (.A(\tholin_riscv.div_shifter[49] ),
    .B(_10720_),
    .Y(_10721_));
 sky130_as_sc_hs__nand3_2 _41468_ (.A(net108),
    .B(_10721_),
    .C(_10722_),
    .Y(_10723_));
 sky130_as_sc_hs__nor2_2 _41472_ (.A(_05656_),
    .B(_06161_),
    .Y(_10727_));
 sky130_as_sc_hs__nand3_2 _41475_ (.A(net412),
    .B(_10728_),
    .C(_10729_),
    .Y(_10730_));
 sky130_as_sc_hs__nor2_2 _41476_ (.A(_10727_),
    .B(_10730_),
    .Y(_10731_));
 sky130_as_sc_hs__and2_2 _41477_ (.A(_10726_),
    .B(_10731_),
    .Y(_10732_));
 sky130_as_sc_hs__nand3_2 _41478_ (.A(_10718_),
    .B(_10723_),
    .C(_10732_),
    .Y(_10733_));
 sky130_as_sc_hs__nor2_2 _41479_ (.A(_10713_),
    .B(_10733_),
    .Y(_10734_));
 sky130_as_sc_hs__and2_2 _41480_ (.A(_10712_),
    .B(_10734_),
    .Y(_10735_));
 sky130_as_sc_hs__and2_2 _41481_ (.A(_10711_),
    .B(_10735_),
    .Y(_10736_));
 sky130_as_sc_hs__nand3_2 _41482_ (.A(_10697_),
    .B(_10701_),
    .C(_10736_),
    .Y(_10737_));
 sky130_as_sc_hs__and2_2 _41483_ (.A(\tholin_riscv.PC[17] ),
    .B(_10547_),
    .Y(_10738_));
 sky130_as_sc_hs__nor2_2 _41484_ (.A(\tholin_riscv.PC[17] ),
    .B(_10547_),
    .Y(_10739_));
 sky130_as_sc_hs__or2_2 _41485_ (.A(_10738_),
    .B(_10739_),
    .Y(_10740_));
 sky130_as_sc_hs__or2_2 _41491_ (.A(\tholin_riscv.PC[17] ),
    .B(net342),
    .Y(_10746_));
 sky130_as_sc_hs__or2_2 _41494_ (.A(_10744_),
    .B(_10747_),
    .Y(_10749_));
 sky130_as_sc_hs__nand3_2 _41495_ (.A(net117),
    .B(_10748_),
    .C(_10749_),
    .Y(_10750_));
 sky130_as_sc_hs__nand3_2 _41496_ (.A(_10741_),
    .B(_10742_),
    .C(_10750_),
    .Y(_10751_));
 sky130_as_sc_hs__nand3_2 _41498_ (.A(_21546_),
    .B(_10737_),
    .C(_10752_),
    .Y(_10753_));
 sky130_as_sc_hs__and2_2 _41503_ (.A(net340),
    .B(net371),
    .Y(_10757_));
 sky130_as_sc_hs__or2_2 _41504_ (.A(_10352_),
    .B(_10757_),
    .Y(_10758_));
 sky130_as_sc_hs__and2_2 _41506_ (.A(net438),
    .B(net418),
    .Y(_10760_));
 sky130_as_sc_hs__and2_2 _41507_ (.A(net83),
    .B(net433),
    .Y(_10761_));
 sky130_as_sc_hs__or2_2 _41508_ (.A(_10760_),
    .B(_10761_),
    .Y(_10762_));
 sky130_as_sc_hs__and2_2 _41510_ (.A(_10762_),
    .B(_10763_),
    .Y(_10764_));
 sky130_as_sc_hs__and2_2 _41511_ (.A(net457),
    .B(net429),
    .Y(_10765_));
 sky130_as_sc_hs__or2_2 _41513_ (.A(_10764_),
    .B(_10765_),
    .Y(_10767_));
 sky130_as_sc_hs__and2_2 _41514_ (.A(_10766_),
    .B(_10767_),
    .Y(_10768_));
 sky130_as_sc_hs__or2_2 _41517_ (.A(_10768_),
    .B(_10769_),
    .Y(_10771_));
 sky130_as_sc_hs__and2_2 _41518_ (.A(_10770_),
    .B(_10771_),
    .Y(_10772_));
 sky130_as_sc_hs__and2_2 _41519_ (.A(net122),
    .B(net466),
    .Y(_10773_));
 sky130_as_sc_hs__and2_2 _41520_ (.A(net468),
    .B(net423),
    .Y(_10774_));
 sky130_as_sc_hs__or2_2 _41521_ (.A(_10773_),
    .B(_10774_),
    .Y(_10775_));
 sky130_as_sc_hs__and2_2 _41523_ (.A(_10775_),
    .B(_10776_),
    .Y(_10777_));
 sky130_as_sc_hs__and2_2 _41524_ (.A(net471),
    .B(net419),
    .Y(_10778_));
 sky130_as_sc_hs__or2_2 _41526_ (.A(_10777_),
    .B(_10778_),
    .Y(_10780_));
 sky130_as_sc_hs__and2_2 _41527_ (.A(_10779_),
    .B(_10780_),
    .Y(_10781_));
 sky130_as_sc_hs__or2_2 _41529_ (.A(_10772_),
    .B(_10781_),
    .Y(_10783_));
 sky130_as_sc_hs__and2_2 _41530_ (.A(_10782_),
    .B(_10783_),
    .Y(_10784_));
 sky130_as_sc_hs__or2_2 _41533_ (.A(_10784_),
    .B(_10785_),
    .Y(_10787_));
 sky130_as_sc_hs__and2_2 _41534_ (.A(_10786_),
    .B(_10787_),
    .Y(_10788_));
 sky130_as_sc_hs__and2_2 _41536_ (.A(net465),
    .B(net74),
    .Y(_10790_));
 sky130_as_sc_hs__nor2b_2 _41537_ (.A(_10402_),
    .Y(_10791_),
    .B(_10790_));
 sky130_as_sc_hs__nor2_2 _41538_ (.A(_10789_),
    .B(_10791_),
    .Y(_10792_));
 sky130_as_sc_hs__and2_2 _41539_ (.A(_10789_),
    .B(_10791_),
    .Y(_10793_));
 sky130_as_sc_hs__nor2_2 _41540_ (.A(_10792_),
    .B(_10793_),
    .Y(_10794_));
 sky130_as_sc_hs__or2_2 _41542_ (.A(_10788_),
    .B(_10794_),
    .Y(_10796_));
 sky130_as_sc_hs__and2_2 _41543_ (.A(_10795_),
    .B(_10796_),
    .Y(_10797_));
 sky130_as_sc_hs__or2_2 _41546_ (.A(_10797_),
    .B(_10798_),
    .Y(_10800_));
 sky130_as_sc_hs__and2_2 _41547_ (.A(_10799_),
    .B(_10800_),
    .Y(_10801_));
 sky130_as_sc_hs__and2_2 _41548_ (.A(net474),
    .B(net425),
    .Y(_10802_));
 sky130_as_sc_hs__or2_2 _41551_ (.A(_10802_),
    .B(_10803_),
    .Y(_10805_));
 sky130_as_sc_hs__and2_2 _41552_ (.A(_10804_),
    .B(_10805_),
    .Y(_10806_));
 sky130_as_sc_hs__or2_2 _41554_ (.A(_10801_),
    .B(_10806_),
    .Y(_10808_));
 sky130_as_sc_hs__and2_2 _41555_ (.A(_10807_),
    .B(_10808_),
    .Y(_10809_));
 sky130_as_sc_hs__or2_2 _41558_ (.A(_10809_),
    .B(_10810_),
    .Y(_10812_));
 sky130_as_sc_hs__and2_2 _41559_ (.A(_10811_),
    .B(_10812_),
    .Y(_10813_));
 sky130_as_sc_hs__and2_2 _41560_ (.A(net434),
    .B(net431),
    .Y(_10814_));
 sky130_as_sc_hs__and2_2 _41561_ (.A(net120),
    .B(net436),
    .Y(_10815_));
 sky130_as_sc_hs__and2_2 _41562_ (.A(net440),
    .B(net428),
    .Y(_10816_));
 sky130_as_sc_hs__and2_2 _41563_ (.A(_10815_),
    .B(_10816_),
    .Y(_10817_));
 sky130_as_sc_hs__nor2_2 _41564_ (.A(_10815_),
    .B(_10816_),
    .Y(_10818_));
 sky130_as_sc_hs__nor2_2 _41565_ (.A(_10817_),
    .B(_10818_),
    .Y(_10819_));
 sky130_as_sc_hs__or2_2 _41567_ (.A(_10814_),
    .B(_10819_),
    .Y(_10821_));
 sky130_as_sc_hs__or2_2 _41569_ (.A(_10621_),
    .B(_10822_),
    .Y(_10823_));
 sky130_as_sc_hs__or2_2 _41572_ (.A(_10638_),
    .B(_10825_),
    .Y(_10826_));
 sky130_as_sc_hs__and2_2 _41574_ (.A(_10826_),
    .B(_10827_),
    .Y(_10828_));
 sky130_as_sc_hs__or2_2 _41576_ (.A(_10813_),
    .B(_10828_),
    .Y(_10830_));
 sky130_as_sc_hs__and2_2 _41577_ (.A(_10829_),
    .B(_10830_),
    .Y(_10831_));
 sky130_as_sc_hs__or2_2 _41580_ (.A(_10831_),
    .B(_10832_),
    .Y(_10834_));
 sky130_as_sc_hs__and2_2 _41581_ (.A(_10833_),
    .B(_10834_),
    .Y(_10835_));
 sky130_as_sc_hs__and2_2 _41584_ (.A(net472),
    .B(net128),
    .Y(_10838_));
 sky130_as_sc_hs__or2_2 _41586_ (.A(_10635_),
    .B(_10838_),
    .Y(_10840_));
 sky130_as_sc_hs__or2_2 _41588_ (.A(_10657_),
    .B(_10841_),
    .Y(_10842_));
 sky130_as_sc_hs__and2_2 _41590_ (.A(_10842_),
    .B(_10843_),
    .Y(_10844_));
 sky130_as_sc_hs__and2_2 _41591_ (.A(net478),
    .B(net421),
    .Y(_10845_));
 sky130_as_sc_hs__or2_2 _41593_ (.A(_10844_),
    .B(_10845_),
    .Y(_10847_));
 sky130_as_sc_hs__and2_2 _41594_ (.A(_10846_),
    .B(_10847_),
    .Y(_10848_));
 sky130_as_sc_hs__or2_2 _41596_ (.A(_10837_),
    .B(_10848_),
    .Y(_10850_));
 sky130_as_sc_hs__and2_2 _41597_ (.A(_10849_),
    .B(_10850_),
    .Y(_10851_));
 sky130_as_sc_hs__or2_2 _41599_ (.A(_10836_),
    .B(_10851_),
    .Y(_10853_));
 sky130_as_sc_hs__and2_2 _41600_ (.A(_10852_),
    .B(_10853_),
    .Y(_10854_));
 sky130_as_sc_hs__or2_2 _41602_ (.A(_10835_),
    .B(_10854_),
    .Y(_10856_));
 sky130_as_sc_hs__and2_2 _41603_ (.A(_10855_),
    .B(_10856_),
    .Y(_10857_));
 sky130_as_sc_hs__or2_2 _41606_ (.A(_10857_),
    .B(_10858_),
    .Y(_10860_));
 sky130_as_sc_hs__and2_2 _41607_ (.A(_10859_),
    .B(_10860_),
    .Y(_10861_));
 sky130_as_sc_hs__or2_2 _41610_ (.A(_10861_),
    .B(_10862_),
    .Y(_10864_));
 sky130_as_sc_hs__and2_2 _41611_ (.A(_10863_),
    .B(_10864_),
    .Y(_10865_));
 sky130_as_sc_hs__or2_2 _41614_ (.A(_10865_),
    .B(_10866_),
    .Y(_10868_));
 sky130_as_sc_hs__or2_2 _41616_ (.A(_10685_),
    .B(_10869_),
    .Y(_10870_));
 sky130_as_sc_hs__and2_2 _41618_ (.A(_10870_),
    .B(_10871_),
    .Y(_10872_));
 sky130_as_sc_hs__and2_2 _41621_ (.A(_10498_),
    .B(_10690_),
    .Y(_10875_));
 sky130_as_sc_hs__or2_2 _41625_ (.A(_10872_),
    .B(_10877_),
    .Y(_10879_));
 sky130_as_sc_hs__and2_2 _41627_ (.A(_10501_),
    .B(_10693_),
    .Y(_10881_));
 sky130_as_sc_hs__or2_2 _41628_ (.A(_05505_),
    .B(_10881_),
    .Y(_10882_));
 sky130_as_sc_hs__and2_2 _41629_ (.A(_10504_),
    .B(_10882_),
    .Y(_10883_));
 sky130_as_sc_hs__or2_2 _41630_ (.A(_10880_),
    .B(_10883_),
    .Y(_10884_));
 sky130_as_sc_hs__nand3_2 _41632_ (.A(net141),
    .B(_10884_),
    .C(_10885_),
    .Y(_10886_));
 sky130_as_sc_hs__or2_2 _41633_ (.A(_05382_),
    .B(_05505_),
    .Y(_10887_));
 sky130_as_sc_hs__and2_2 _41634_ (.A(_10508_),
    .B(_10887_),
    .Y(_10888_));
 sky130_as_sc_hs__or2_2 _41635_ (.A(_05435_),
    .B(_10888_),
    .Y(_10889_));
 sky130_as_sc_hs__nand3_2 _41637_ (.A(net138),
    .B(_10889_),
    .C(_10890_),
    .Y(_10891_));
 sky130_as_sc_hs__or2_2 _41641_ (.A(_05648_),
    .B(_10893_),
    .Y(_10895_));
 sky130_as_sc_hs__or2_2 _41644_ (.A(_05649_),
    .B(_05886_),
    .Y(_10898_));
 sky130_as_sc_hs__nand3_2 _41647_ (.A(net118),
    .B(_10897_),
    .C(_10900_),
    .Y(_10901_));
 sky130_as_sc_hs__and2_2 _41649_ (.A(net140),
    .B(_09865_),
    .Y(_10903_));
 sky130_as_sc_hs__or2_2 _41650_ (.A(\tholin_riscv.div_res[17] ),
    .B(_10714_),
    .Y(_10904_));
 sky130_as_sc_hs__and2_2 _41651_ (.A(net415),
    .B(_10904_),
    .Y(_10905_));
 sky130_as_sc_hs__or2_2 _41653_ (.A(\tholin_riscv.div_res[18] ),
    .B(_10905_),
    .Y(_10907_));
 sky130_as_sc_hs__nand3_2 _41654_ (.A(net110),
    .B(_10906_),
    .C(_10907_),
    .Y(_10908_));
 sky130_as_sc_hs__or2_2 _41655_ (.A(\tholin_riscv.div_shifter[49] ),
    .B(_10719_),
    .Y(_10909_));
 sky130_as_sc_hs__and2_2 _41656_ (.A(_21655_),
    .B(_10909_),
    .Y(_10910_));
 sky130_as_sc_hs__or2_2 _41658_ (.A(\tholin_riscv.div_shifter[50] ),
    .B(_10910_),
    .Y(_10912_));
 sky130_as_sc_hs__nand3_2 _41659_ (.A(net107),
    .B(_10911_),
    .C(_10912_),
    .Y(_10913_));
 sky130_as_sc_hs__and2_2 _41660_ (.A(_05648_),
    .B(_06538_),
    .Y(_10914_));
 sky130_as_sc_hs__or2_2 _41662_ (.A(_05646_),
    .B(_06161_),
    .Y(_10916_));
 sky130_as_sc_hs__and2_2 _41665_ (.A(_10917_),
    .B(_10918_),
    .Y(_10919_));
 sky130_as_sc_hs__and2_2 _41666_ (.A(net413),
    .B(_10919_),
    .Y(_10920_));
 sky130_as_sc_hs__nand3_2 _41667_ (.A(_10915_),
    .B(_10916_),
    .C(_10920_),
    .Y(_10921_));
 sky130_as_sc_hs__nor2_2 _41668_ (.A(_10914_),
    .B(_10921_),
    .Y(_10922_));
 sky130_as_sc_hs__nand3_2 _41669_ (.A(_10908_),
    .B(_10913_),
    .C(_10922_),
    .Y(_10923_));
 sky130_as_sc_hs__nor2_2 _41670_ (.A(_10903_),
    .B(_10923_),
    .Y(_10924_));
 sky130_as_sc_hs__and2_2 _41671_ (.A(_10902_),
    .B(_10924_),
    .Y(_10925_));
 sky130_as_sc_hs__and2_2 _41672_ (.A(_10901_),
    .B(_10925_),
    .Y(_10926_));
 sky130_as_sc_hs__nand3_2 _41673_ (.A(_10886_),
    .B(_10891_),
    .C(_10926_),
    .Y(_10927_));
 sky130_as_sc_hs__and2_2 _41674_ (.A(\tholin_riscv.PC[18] ),
    .B(_10738_),
    .Y(_10928_));
 sky130_as_sc_hs__nor2_2 _41675_ (.A(\tholin_riscv.PC[18] ),
    .B(_10738_),
    .Y(_10929_));
 sky130_as_sc_hs__or2_2 _41676_ (.A(_10928_),
    .B(_10929_),
    .Y(_10930_));
 sky130_as_sc_hs__or2_2 _41682_ (.A(\tholin_riscv.PC[18] ),
    .B(net337),
    .Y(_10936_));
 sky130_as_sc_hs__or2_2 _41684_ (.A(_10934_),
    .B(_10937_),
    .Y(_10938_));
 sky130_as_sc_hs__nand3_2 _41686_ (.A(net117),
    .B(_10938_),
    .C(_10939_),
    .Y(_10940_));
 sky130_as_sc_hs__nand3_2 _41687_ (.A(_10931_),
    .B(_10932_),
    .C(_10940_),
    .Y(_10941_));
 sky130_as_sc_hs__nand3_2 _41689_ (.A(_21546_),
    .B(_10927_),
    .C(_10942_),
    .Y(_10943_));
 sky130_as_sc_hs__and2_2 _41694_ (.A(net335),
    .B(net371),
    .Y(_10947_));
 sky130_as_sc_hs__or2_2 _41695_ (.A(_10352_),
    .B(_10947_),
    .Y(_10948_));
 sky130_as_sc_hs__and2_2 _41697_ (.A(_10870_),
    .B(_10878_),
    .Y(_10950_));
 sky130_as_sc_hs__and2_2 _41698_ (.A(net472),
    .B(net418),
    .Y(_10951_));
 sky130_as_sc_hs__and2_2 _41699_ (.A(net433),
    .B(net431),
    .Y(_10952_));
 sky130_as_sc_hs__or2_2 _41700_ (.A(_10951_),
    .B(_10952_),
    .Y(_10953_));
 sky130_as_sc_hs__and2_2 _41702_ (.A(_10953_),
    .B(_10954_),
    .Y(_10955_));
 sky130_as_sc_hs__and2_2 _41703_ (.A(net457),
    .B(net427),
    .Y(_10956_));
 sky130_as_sc_hs__or2_2 _41705_ (.A(_10955_),
    .B(_10956_),
    .Y(_10958_));
 sky130_as_sc_hs__and2_2 _41706_ (.A(_10957_),
    .B(_10958_),
    .Y(_10959_));
 sky130_as_sc_hs__or2_2 _41709_ (.A(_10959_),
    .B(_10960_),
    .Y(_10962_));
 sky130_as_sc_hs__and2_2 _41710_ (.A(_10961_),
    .B(_10962_),
    .Y(_10963_));
 sky130_as_sc_hs__and2_2 _41711_ (.A(net466),
    .B(net423),
    .Y(_10964_));
 sky130_as_sc_hs__and2_2 _41712_ (.A(net468),
    .B(net419),
    .Y(_10965_));
 sky130_as_sc_hs__or2_2 _41713_ (.A(_10964_),
    .B(_10965_),
    .Y(_10966_));
 sky130_as_sc_hs__and2_2 _41715_ (.A(_10966_),
    .B(_10967_),
    .Y(_10968_));
 sky130_as_sc_hs__and2_2 _41716_ (.A(net471),
    .B(net74),
    .Y(_10969_));
 sky130_as_sc_hs__or2_2 _41718_ (.A(_10968_),
    .B(_10969_),
    .Y(_10971_));
 sky130_as_sc_hs__and2_2 _41719_ (.A(_10970_),
    .B(_10971_),
    .Y(_10972_));
 sky130_as_sc_hs__or2_2 _41721_ (.A(_10963_),
    .B(_10972_),
    .Y(_10974_));
 sky130_as_sc_hs__and2_2 _41722_ (.A(_10973_),
    .B(_10974_),
    .Y(_10975_));
 sky130_as_sc_hs__or2_2 _41725_ (.A(_10975_),
    .B(_10976_),
    .Y(_10978_));
 sky130_as_sc_hs__and2_2 _41726_ (.A(_10977_),
    .B(_10978_),
    .Y(_10979_));
 sky130_as_sc_hs__or2_2 _41729_ (.A(_10979_),
    .B(_10980_),
    .Y(_10982_));
 sky130_as_sc_hs__and2_2 _41730_ (.A(_10981_),
    .B(_10982_),
    .Y(_10983_));
 sky130_as_sc_hs__or2_2 _41733_ (.A(_10983_),
    .B(_10984_),
    .Y(_10986_));
 sky130_as_sc_hs__and2_2 _41734_ (.A(_10985_),
    .B(_10986_),
    .Y(_10987_));
 sky130_as_sc_hs__and2_2 _41735_ (.A(net83),
    .B(net425),
    .Y(_10988_));
 sky130_as_sc_hs__or2_2 _41736_ (.A(_10402_),
    .B(_10789_),
    .Y(_10989_));
 sky130_as_sc_hs__and2_2 _41737_ (.A(_10790_),
    .B(_10989_),
    .Y(_10990_));
 sky130_as_sc_hs__or2_2 _41739_ (.A(_10988_),
    .B(_10990_),
    .Y(_10992_));
 sky130_as_sc_hs__and2_2 _41740_ (.A(_10991_),
    .B(_10992_),
    .Y(_10993_));
 sky130_as_sc_hs__or2_2 _41742_ (.A(_10987_),
    .B(_10993_),
    .Y(_10995_));
 sky130_as_sc_hs__and2_2 _41743_ (.A(_10994_),
    .B(_10995_),
    .Y(_10996_));
 sky130_as_sc_hs__or2_2 _41746_ (.A(_10996_),
    .B(_10997_),
    .Y(_10999_));
 sky130_as_sc_hs__and2_2 _41747_ (.A(_10998_),
    .B(_10999_),
    .Y(_11000_));
 sky130_as_sc_hs__and2_2 _41748_ (.A(net434),
    .B(net430),
    .Y(_11001_));
 sky130_as_sc_hs__and2_2 _41749_ (.A(net122),
    .B(net436),
    .Y(_11002_));
 sky130_as_sc_hs__and2_2 _41750_ (.A(net120),
    .B(net440),
    .Y(_11003_));
 sky130_as_sc_hs__and2_2 _41751_ (.A(_11002_),
    .B(_11003_),
    .Y(_11004_));
 sky130_as_sc_hs__or2_2 _41752_ (.A(_11002_),
    .B(_11003_),
    .Y(_11005_));
 sky130_as_sc_hs__nor2b_2 _41753_ (.A(_11004_),
    .Y(_11006_),
    .B(_11005_));
 sky130_as_sc_hs__or2_2 _41755_ (.A(_11001_),
    .B(_11006_),
    .Y(_11008_));
 sky130_as_sc_hs__or2_2 _41757_ (.A(_10804_),
    .B(_11009_),
    .Y(_11010_));
 sky130_as_sc_hs__or2_2 _41760_ (.A(_10820_),
    .B(_11012_),
    .Y(_11013_));
 sky130_as_sc_hs__and2_2 _41762_ (.A(_11013_),
    .B(_11014_),
    .Y(_11015_));
 sky130_as_sc_hs__or2_2 _41764_ (.A(_11000_),
    .B(_11015_),
    .Y(_11017_));
 sky130_as_sc_hs__and2_2 _41765_ (.A(_11016_),
    .B(_11017_),
    .Y(_11018_));
 sky130_as_sc_hs__or2_2 _41768_ (.A(_11018_),
    .B(_11019_),
    .Y(_11021_));
 sky130_as_sc_hs__and2_2 _41769_ (.A(_11020_),
    .B(_11021_),
    .Y(_11022_));
 sky130_as_sc_hs__and2_2 _41772_ (.A(net478),
    .B(net128),
    .Y(_11025_));
 sky130_as_sc_hs__or2_2 _41774_ (.A(_10817_),
    .B(_11025_),
    .Y(_11027_));
 sky130_as_sc_hs__or2_2 _41776_ (.A(_10839_),
    .B(_11028_),
    .Y(_11029_));
 sky130_as_sc_hs__and2_2 _41778_ (.A(_11029_),
    .B(_11030_),
    .Y(_11031_));
 sky130_as_sc_hs__and2_2 _41779_ (.A(net474),
    .B(net421),
    .Y(_11032_));
 sky130_as_sc_hs__or2_2 _41781_ (.A(_11031_),
    .B(_11032_),
    .Y(_11034_));
 sky130_as_sc_hs__and2_2 _41782_ (.A(_11033_),
    .B(_11034_),
    .Y(_11035_));
 sky130_as_sc_hs__or2_2 _41784_ (.A(_11024_),
    .B(_11035_),
    .Y(_11037_));
 sky130_as_sc_hs__and2_2 _41785_ (.A(_11036_),
    .B(_11037_),
    .Y(_11038_));
 sky130_as_sc_hs__or2_2 _41787_ (.A(_11023_),
    .B(_11038_),
    .Y(_11040_));
 sky130_as_sc_hs__and2_2 _41788_ (.A(_11039_),
    .B(_11040_),
    .Y(_11041_));
 sky130_as_sc_hs__or2_2 _41790_ (.A(_11022_),
    .B(_11041_),
    .Y(_11043_));
 sky130_as_sc_hs__and2_2 _41791_ (.A(_11042_),
    .B(_11043_),
    .Y(_11044_));
 sky130_as_sc_hs__or2_2 _41794_ (.A(_11044_),
    .B(_11045_),
    .Y(_11047_));
 sky130_as_sc_hs__and2_2 _41795_ (.A(_11046_),
    .B(_11047_),
    .Y(_11048_));
 sky130_as_sc_hs__or2_2 _41798_ (.A(_11048_),
    .B(_11049_),
    .Y(_11051_));
 sky130_as_sc_hs__and2_2 _41799_ (.A(_11050_),
    .B(_11051_),
    .Y(_11052_));
 sky130_as_sc_hs__or2_2 _41802_ (.A(_11052_),
    .B(_11053_),
    .Y(_11055_));
 sky130_as_sc_hs__and2_2 _41803_ (.A(_11054_),
    .B(_11055_),
    .Y(_11056_));
 sky130_as_sc_hs__nor2_2 _41804_ (.A(_10867_),
    .B(_11056_),
    .Y(_11057_));
 sky130_as_sc_hs__and2_2 _41805_ (.A(_10867_),
    .B(_11056_),
    .Y(_11058_));
 sky130_as_sc_hs__or2_2 _41806_ (.A(_11057_),
    .B(_11058_),
    .Y(_11059_));
 sky130_as_sc_hs__or2_2 _41808_ (.A(_10950_),
    .B(_11059_),
    .Y(_11061_));
 sky130_as_sc_hs__and2_2 _41809_ (.A(_11060_),
    .B(_11061_),
    .Y(_11062_));
 sky130_as_sc_hs__and2_2 _41810_ (.A(_10880_),
    .B(_10881_),
    .Y(_11063_));
 sky130_as_sc_hs__or2_2 _41811_ (.A(_05505_),
    .B(_11063_),
    .Y(_11064_));
 sky130_as_sc_hs__and2_2 _41812_ (.A(_10504_),
    .B(_11064_),
    .Y(_11065_));
 sky130_as_sc_hs__or2_2 _41813_ (.A(_11062_),
    .B(_11065_),
    .Y(_11066_));
 sky130_as_sc_hs__nand3_2 _41815_ (.A(net142),
    .B(_11066_),
    .C(_11067_),
    .Y(_11068_));
 sky130_as_sc_hs__or2_2 _41816_ (.A(_05437_),
    .B(_05505_),
    .Y(_11069_));
 sky130_as_sc_hs__or2_2 _41817_ (.A(_05441_),
    .B(_11069_),
    .Y(_11070_));
 sky130_as_sc_hs__nand3_2 _41819_ (.A(net138),
    .B(_11070_),
    .C(_11071_),
    .Y(_11072_));
 sky130_as_sc_hs__or2_2 _41822_ (.A(_05638_),
    .B(_11073_),
    .Y(_11075_));
 sky130_as_sc_hs__or2_2 _41825_ (.A(_05639_),
    .B(_05888_),
    .Y(_11078_));
 sky130_as_sc_hs__nand3_2 _41828_ (.A(net119),
    .B(_11077_),
    .C(_11080_),
    .Y(_11081_));
 sky130_as_sc_hs__and2_2 _41830_ (.A(net140),
    .B(_09643_),
    .Y(_11083_));
 sky130_as_sc_hs__or2_2 _41831_ (.A(\tholin_riscv.div_shifter[50] ),
    .B(_10909_),
    .Y(_11084_));
 sky130_as_sc_hs__and2_2 _41832_ (.A(_21655_),
    .B(_11084_),
    .Y(_11085_));
 sky130_as_sc_hs__or2_2 _41834_ (.A(\tholin_riscv.div_shifter[51] ),
    .B(_11085_),
    .Y(_11087_));
 sky130_as_sc_hs__nand3_2 _41835_ (.A(net107),
    .B(_11086_),
    .C(_11087_),
    .Y(_11088_));
 sky130_as_sc_hs__or2_2 _41836_ (.A(\tholin_riscv.div_res[18] ),
    .B(_10904_),
    .Y(_11089_));
 sky130_as_sc_hs__and2_2 _41837_ (.A(net415),
    .B(_11089_),
    .Y(_11090_));
 sky130_as_sc_hs__or2_2 _41839_ (.A(\tholin_riscv.div_res[19] ),
    .B(_11090_),
    .Y(_11092_));
 sky130_as_sc_hs__nand3_2 _41840_ (.A(net111),
    .B(_11091_),
    .C(_11092_),
    .Y(_11093_));
 sky130_as_sc_hs__and2_2 _41841_ (.A(_05638_),
    .B(_06538_),
    .Y(_11094_));
 sky130_as_sc_hs__or2_2 _41843_ (.A(_05636_),
    .B(_06161_),
    .Y(_11096_));
 sky130_as_sc_hs__and2_2 _41846_ (.A(_11097_),
    .B(_11098_),
    .Y(_11099_));
 sky130_as_sc_hs__and2_2 _41847_ (.A(net413),
    .B(_11099_),
    .Y(_11100_));
 sky130_as_sc_hs__nand3_2 _41848_ (.A(_11095_),
    .B(_11096_),
    .C(_11100_),
    .Y(_11101_));
 sky130_as_sc_hs__nor2_2 _41849_ (.A(_11094_),
    .B(_11101_),
    .Y(_11102_));
 sky130_as_sc_hs__nand3_2 _41850_ (.A(_11088_),
    .B(_11093_),
    .C(_11102_),
    .Y(_11103_));
 sky130_as_sc_hs__nor2_2 _41851_ (.A(_11083_),
    .B(_11103_),
    .Y(_11104_));
 sky130_as_sc_hs__and2_2 _41852_ (.A(_11082_),
    .B(_11104_),
    .Y(_11105_));
 sky130_as_sc_hs__and2_2 _41853_ (.A(_11081_),
    .B(_11105_),
    .Y(_11106_));
 sky130_as_sc_hs__nand3_2 _41854_ (.A(_11068_),
    .B(_11072_),
    .C(_11106_),
    .Y(_11107_));
 sky130_as_sc_hs__and2_2 _41855_ (.A(\tholin_riscv.PC[19] ),
    .B(_10928_),
    .Y(_11108_));
 sky130_as_sc_hs__nor2_2 _41856_ (.A(\tholin_riscv.PC[19] ),
    .B(_10928_),
    .Y(_11109_));
 sky130_as_sc_hs__nor2_2 _41857_ (.A(_11108_),
    .B(_11109_),
    .Y(_11110_));
 sky130_as_sc_hs__inv_2 _41858_ (.Y(_11111_),
    .A(_11110_));
 sky130_as_sc_hs__and2_2 _41859_ (.A(_21573_),
    .B(_11110_),
    .Y(_11112_));
 sky130_as_sc_hs__or2_2 _41863_ (.A(\tholin_riscv.PC[19] ),
    .B(net336),
    .Y(_11116_));
 sky130_as_sc_hs__and2_2 _41864_ (.A(_11115_),
    .B(_11116_),
    .Y(_11117_));
 sky130_as_sc_hs__or2_2 _41866_ (.A(_11114_),
    .B(_11117_),
    .Y(_11119_));
 sky130_as_sc_hs__nand3_2 _41867_ (.A(net117),
    .B(_11118_),
    .C(_11119_),
    .Y(_11120_));
 sky130_as_sc_hs__nand3_2 _41869_ (.A(_21569_),
    .B(_11120_),
    .C(_11121_),
    .Y(_11122_));
 sky130_as_sc_hs__or2_2 _41870_ (.A(_11112_),
    .B(_11122_),
    .Y(_11123_));
 sky130_as_sc_hs__nand3_2 _41871_ (.A(_21546_),
    .B(_11107_),
    .C(_11123_),
    .Y(_11124_));
 sky130_as_sc_hs__and2_2 _41876_ (.A(\tholin_riscv.Iimm[0] ),
    .B(net371),
    .Y(_11128_));
 sky130_as_sc_hs__or2_2 _41877_ (.A(_10352_),
    .B(_11128_),
    .Y(_11129_));
 sky130_as_sc_hs__and2_2 _41879_ (.A(_10872_),
    .B(_11059_),
    .Y(_11131_));
 sky130_as_sc_hs__nand3_2 _41880_ (.A(_10369_),
    .B(_10875_),
    .C(_11131_),
    .Y(_11132_));
 sky130_as_sc_hs__nand2b_2 _41881_ (.B(_11131_),
    .Y(_11133_),
    .A(_10874_));
 sky130_as_sc_hs__nand3_2 _41884_ (.A(_11132_),
    .B(_11133_),
    .C(_11135_),
    .Y(_11136_));
 sky130_as_sc_hs__and2_2 _41885_ (.A(net431),
    .B(net425),
    .Y(_11137_));
 sky130_as_sc_hs__and2_2 _41886_ (.A(net478),
    .B(net418),
    .Y(_11138_));
 sky130_as_sc_hs__and2_2 _41887_ (.A(net433),
    .B(net429),
    .Y(_11139_));
 sky130_as_sc_hs__or2_2 _41889_ (.A(_11138_),
    .B(_11139_),
    .Y(_11141_));
 sky130_as_sc_hs__and2_2 _41890_ (.A(_11140_),
    .B(_11141_),
    .Y(_11142_));
 sky130_as_sc_hs__and2_2 _41891_ (.A(net120),
    .B(net457),
    .Y(_11143_));
 sky130_as_sc_hs__or2_2 _41893_ (.A(_11142_),
    .B(_11143_),
    .Y(_11145_));
 sky130_as_sc_hs__and2_2 _41894_ (.A(_11144_),
    .B(_11145_),
    .Y(_11146_));
 sky130_as_sc_hs__or2_2 _41897_ (.A(_11146_),
    .B(_11147_),
    .Y(_11149_));
 sky130_as_sc_hs__and2_2 _41898_ (.A(_11148_),
    .B(_11149_),
    .Y(_11150_));
 sky130_as_sc_hs__and2_2 _41899_ (.A(net466),
    .B(net419),
    .Y(_11151_));
 sky130_as_sc_hs__and2_2 _41900_ (.A(net468),
    .B(net74),
    .Y(_11152_));
 sky130_as_sc_hs__or2_2 _41902_ (.A(_11151_),
    .B(_11152_),
    .Y(_11154_));
 sky130_as_sc_hs__and2_2 _41903_ (.A(_11153_),
    .B(_11154_),
    .Y(_11155_));
 sky130_as_sc_hs__or2_2 _41905_ (.A(_11150_),
    .B(_11155_),
    .Y(_11157_));
 sky130_as_sc_hs__and2_2 _41906_ (.A(_11156_),
    .B(_11157_),
    .Y(_11158_));
 sky130_as_sc_hs__or2_2 _41909_ (.A(_11158_),
    .B(_11159_),
    .Y(_11161_));
 sky130_as_sc_hs__and2_2 _41910_ (.A(_11160_),
    .B(_11161_),
    .Y(_11162_));
 sky130_as_sc_hs__or2_2 _41913_ (.A(_11162_),
    .B(_11163_),
    .Y(_11165_));
 sky130_as_sc_hs__and2_2 _41914_ (.A(_11164_),
    .B(_11165_),
    .Y(_11166_));
 sky130_as_sc_hs__or2_2 _41917_ (.A(_11166_),
    .B(_11167_),
    .Y(_11169_));
 sky130_as_sc_hs__and2_2 _41918_ (.A(_11168_),
    .B(_11169_),
    .Y(_11170_));
 sky130_as_sc_hs__or2_2 _41920_ (.A(_11137_),
    .B(_11170_),
    .Y(_11172_));
 sky130_as_sc_hs__and2_2 _41921_ (.A(_11171_),
    .B(_11172_),
    .Y(_11173_));
 sky130_as_sc_hs__or2_2 _41924_ (.A(_11173_),
    .B(_11174_),
    .Y(_11176_));
 sky130_as_sc_hs__and2_2 _41925_ (.A(_11175_),
    .B(_11176_),
    .Y(_11177_));
 sky130_as_sc_hs__and2_2 _41926_ (.A(net434),
    .B(net427),
    .Y(_11178_));
 sky130_as_sc_hs__and2_2 _41927_ (.A(net436),
    .B(net423),
    .Y(_11179_));
 sky130_as_sc_hs__and2_2 _41928_ (.A(net123),
    .B(net440),
    .Y(_11180_));
 sky130_as_sc_hs__and2_2 _41929_ (.A(_11179_),
    .B(_11180_),
    .Y(_11181_));
 sky130_as_sc_hs__or2_2 _41930_ (.A(_11179_),
    .B(_11180_),
    .Y(_11182_));
 sky130_as_sc_hs__nor2b_2 _41931_ (.A(_11181_),
    .Y(_11183_),
    .B(_11182_));
 sky130_as_sc_hs__or2_2 _41933_ (.A(_11178_),
    .B(_11183_),
    .Y(_11185_));
 sky130_as_sc_hs__or2_2 _41935_ (.A(_10991_),
    .B(_11186_),
    .Y(_11187_));
 sky130_as_sc_hs__or2_2 _41938_ (.A(_11007_),
    .B(_11189_),
    .Y(_11190_));
 sky130_as_sc_hs__and2_2 _41940_ (.A(_11190_),
    .B(_11191_),
    .Y(_11192_));
 sky130_as_sc_hs__or2_2 _41942_ (.A(_11177_),
    .B(_11192_),
    .Y(_11194_));
 sky130_as_sc_hs__and2_2 _41943_ (.A(_11193_),
    .B(_11194_),
    .Y(_11195_));
 sky130_as_sc_hs__or2_2 _41946_ (.A(_11195_),
    .B(_11196_),
    .Y(_11198_));
 sky130_as_sc_hs__and2_2 _41947_ (.A(_11197_),
    .B(_11198_),
    .Y(_11199_));
 sky130_as_sc_hs__and2_2 _41950_ (.A(net83),
    .B(net421),
    .Y(_11202_));
 sky130_as_sc_hs__and2_2 _41951_ (.A(net474),
    .B(net128),
    .Y(_11203_));
 sky130_as_sc_hs__or2_2 _41953_ (.A(_11004_),
    .B(_11203_),
    .Y(_11205_));
 sky130_as_sc_hs__or2_2 _41955_ (.A(_11026_),
    .B(_11206_),
    .Y(_11207_));
 sky130_as_sc_hs__and2_2 _41957_ (.A(_11207_),
    .B(_11208_),
    .Y(_11209_));
 sky130_as_sc_hs__or2_2 _41959_ (.A(_11202_),
    .B(_11209_),
    .Y(_11211_));
 sky130_as_sc_hs__and2_2 _41960_ (.A(_11210_),
    .B(_11211_),
    .Y(_11212_));
 sky130_as_sc_hs__or2_2 _41962_ (.A(_11201_),
    .B(_11212_),
    .Y(_11214_));
 sky130_as_sc_hs__and2_2 _41963_ (.A(_11213_),
    .B(_11214_),
    .Y(_11215_));
 sky130_as_sc_hs__or2_2 _41965_ (.A(_11200_),
    .B(_11215_),
    .Y(_11217_));
 sky130_as_sc_hs__and2_2 _41966_ (.A(_11216_),
    .B(_11217_),
    .Y(_11218_));
 sky130_as_sc_hs__or2_2 _41968_ (.A(_11199_),
    .B(_11218_),
    .Y(_11220_));
 sky130_as_sc_hs__and2_2 _41969_ (.A(_11219_),
    .B(_11220_),
    .Y(_11221_));
 sky130_as_sc_hs__or2_2 _41972_ (.A(_11221_),
    .B(_11222_),
    .Y(_11224_));
 sky130_as_sc_hs__and2_2 _41973_ (.A(_11223_),
    .B(_11224_),
    .Y(_11225_));
 sky130_as_sc_hs__or2_2 _41976_ (.A(_11225_),
    .B(_11226_),
    .Y(_11228_));
 sky130_as_sc_hs__and2_2 _41977_ (.A(_11227_),
    .B(_11228_),
    .Y(_11229_));
 sky130_as_sc_hs__or2_2 _41980_ (.A(_11229_),
    .B(_11230_),
    .Y(_11232_));
 sky130_as_sc_hs__or2_2 _41982_ (.A(_11054_),
    .B(_11233_),
    .Y(_11234_));
 sky130_as_sc_hs__and2_2 _41984_ (.A(_11234_),
    .B(_11235_),
    .Y(_11236_));
 sky130_as_sc_hs__inv_2 _41986_ (.Y(_11238_),
    .A(_11237_));
 sky130_as_sc_hs__nor2_2 _41987_ (.A(_11136_),
    .B(_11236_),
    .Y(_11239_));
 sky130_as_sc_hs__or2_2 _41988_ (.A(_11238_),
    .B(_11239_),
    .Y(_11240_));
 sky130_as_sc_hs__and2_2 _41989_ (.A(_11062_),
    .B(_11063_),
    .Y(_11241_));
 sky130_as_sc_hs__or2_2 _41993_ (.A(_11240_),
    .B(_11243_),
    .Y(_11245_));
 sky130_as_sc_hs__nand3_2 _41994_ (.A(net141),
    .B(_11244_),
    .C(_11245_),
    .Y(_11246_));
 sky130_as_sc_hs__or2_2 _41995_ (.A(_05442_),
    .B(_05505_),
    .Y(_11247_));
 sky130_as_sc_hs__or2_2 _41996_ (.A(_05445_),
    .B(_11247_),
    .Y(_11248_));
 sky130_as_sc_hs__nand3_2 _41998_ (.A(net138),
    .B(_11248_),
    .C(_11249_),
    .Y(_11250_));
 sky130_as_sc_hs__or2_2 _42001_ (.A(_05628_),
    .B(_11251_),
    .Y(_11253_));
 sky130_as_sc_hs__or2_2 _42004_ (.A(_05629_),
    .B(_05890_),
    .Y(_11256_));
 sky130_as_sc_hs__nand3_2 _42007_ (.A(net118),
    .B(_11255_),
    .C(_11258_),
    .Y(_11259_));
 sky130_as_sc_hs__and2_2 _42008_ (.A(net140),
    .B(_09409_),
    .Y(_11260_));
 sky130_as_sc_hs__or2_2 _42010_ (.A(\tholin_riscv.div_shifter[51] ),
    .B(_11084_),
    .Y(_11262_));
 sky130_as_sc_hs__and2_2 _42011_ (.A(_21655_),
    .B(_11262_),
    .Y(_11263_));
 sky130_as_sc_hs__or2_2 _42013_ (.A(\tholin_riscv.div_shifter[52] ),
    .B(_11263_),
    .Y(_11265_));
 sky130_as_sc_hs__nand3_2 _42014_ (.A(net107),
    .B(_11264_),
    .C(_11265_),
    .Y(_11266_));
 sky130_as_sc_hs__or2_2 _42015_ (.A(\tholin_riscv.div_res[19] ),
    .B(_11089_),
    .Y(_11267_));
 sky130_as_sc_hs__and2_2 _42016_ (.A(net415),
    .B(_11267_),
    .Y(_11268_));
 sky130_as_sc_hs__or2_2 _42018_ (.A(\tholin_riscv.div_res[20] ),
    .B(_11268_),
    .Y(_11270_));
 sky130_as_sc_hs__nand3_2 _42019_ (.A(net111),
    .B(_11269_),
    .C(_11270_),
    .Y(_11271_));
 sky130_as_sc_hs__and2_2 _42020_ (.A(_05628_),
    .B(_06538_),
    .Y(_11272_));
 sky130_as_sc_hs__or2_2 _42022_ (.A(_05626_),
    .B(_06161_),
    .Y(_11274_));
 sky130_as_sc_hs__and2_2 _42025_ (.A(_11275_),
    .B(_11276_),
    .Y(_11277_));
 sky130_as_sc_hs__and2_2 _42026_ (.A(net413),
    .B(_11277_),
    .Y(_11278_));
 sky130_as_sc_hs__nand3_2 _42027_ (.A(_11273_),
    .B(_11274_),
    .C(_11278_),
    .Y(_11279_));
 sky130_as_sc_hs__nor2_2 _42028_ (.A(_11272_),
    .B(_11279_),
    .Y(_11280_));
 sky130_as_sc_hs__nand3_2 _42029_ (.A(_11266_),
    .B(_11271_),
    .C(_11280_),
    .Y(_11281_));
 sky130_as_sc_hs__nor2_2 _42030_ (.A(_11260_),
    .B(_11281_),
    .Y(_11282_));
 sky130_as_sc_hs__and2_2 _42031_ (.A(_11261_),
    .B(_11282_),
    .Y(_11283_));
 sky130_as_sc_hs__and2_2 _42032_ (.A(_11259_),
    .B(_11283_),
    .Y(_11284_));
 sky130_as_sc_hs__nand3_2 _42033_ (.A(_11246_),
    .B(_11250_),
    .C(_11284_),
    .Y(_11285_));
 sky130_as_sc_hs__and2_2 _42034_ (.A(\tholin_riscv.PC[20] ),
    .B(_11108_),
    .Y(_11286_));
 sky130_as_sc_hs__nor2_2 _42035_ (.A(\tholin_riscv.PC[20] ),
    .B(_11108_),
    .Y(_11287_));
 sky130_as_sc_hs__or2_2 _42036_ (.A(_11286_),
    .B(_11287_),
    .Y(_11288_));
 sky130_as_sc_hs__or2_2 _42038_ (.A(\tholin_riscv.Iimm[0] ),
    .B(_21590_),
    .Y(_11290_));
 sky130_as_sc_hs__or2_2 _42042_ (.A(\tholin_riscv.PC[20] ),
    .B(\tholin_riscv.Iimm[0] ),
    .Y(_11294_));
 sky130_as_sc_hs__or2_2 _42044_ (.A(_11292_),
    .B(_11295_),
    .Y(_11296_));
 sky130_as_sc_hs__nand3_2 _42046_ (.A(net117),
    .B(_11296_),
    .C(_11297_),
    .Y(_11298_));
 sky130_as_sc_hs__nand3_2 _42047_ (.A(_11289_),
    .B(_11290_),
    .C(_11298_),
    .Y(_11299_));
 sky130_as_sc_hs__nand3_2 _42049_ (.A(_21546_),
    .B(_11285_),
    .C(_11300_),
    .Y(_11301_));
 sky130_as_sc_hs__and2_2 _42054_ (.A(\tholin_riscv.Iimm[1] ),
    .B(net371),
    .Y(_11305_));
 sky130_as_sc_hs__or2_2 _42055_ (.A(_10352_),
    .B(_11305_),
    .Y(_11306_));
 sky130_as_sc_hs__and2_2 _42057_ (.A(_11234_),
    .B(_11237_),
    .Y(_11308_));
 sky130_as_sc_hs__and2_2 _42058_ (.A(net430),
    .B(net425),
    .Y(_11309_));
 sky130_as_sc_hs__and2_2 _42059_ (.A(net466),
    .B(net74),
    .Y(_11310_));
 sky130_as_sc_hs__and2_2 _42060_ (.A(net474),
    .B(net418),
    .Y(_11311_));
 sky130_as_sc_hs__and2_2 _42061_ (.A(net433),
    .B(net427),
    .Y(_11312_));
 sky130_as_sc_hs__or2_2 _42063_ (.A(_11311_),
    .B(_11312_),
    .Y(_11314_));
 sky130_as_sc_hs__and2_2 _42064_ (.A(_11313_),
    .B(_11314_),
    .Y(_11315_));
 sky130_as_sc_hs__and2_2 _42065_ (.A(net122),
    .B(net457),
    .Y(_11316_));
 sky130_as_sc_hs__or2_2 _42067_ (.A(_11315_),
    .B(_11316_),
    .Y(_11318_));
 sky130_as_sc_hs__and2_2 _42068_ (.A(_11317_),
    .B(_11318_),
    .Y(_11319_));
 sky130_as_sc_hs__or2_2 _42071_ (.A(_11319_),
    .B(_11320_),
    .Y(_11322_));
 sky130_as_sc_hs__and2_2 _42072_ (.A(_11321_),
    .B(_11322_),
    .Y(_11323_));
 sky130_as_sc_hs__or2_2 _42074_ (.A(_11310_),
    .B(_11323_),
    .Y(_11325_));
 sky130_as_sc_hs__and2_2 _42075_ (.A(_11324_),
    .B(_11325_),
    .Y(_11326_));
 sky130_as_sc_hs__or2_2 _42078_ (.A(_11326_),
    .B(_11327_),
    .Y(_11329_));
 sky130_as_sc_hs__or2_2 _42080_ (.A(_11153_),
    .B(_11330_),
    .Y(_11331_));
 sky130_as_sc_hs__and2_2 _42082_ (.A(_11331_),
    .B(_11332_),
    .Y(_11333_));
 sky130_as_sc_hs__or2_2 _42085_ (.A(_11333_),
    .B(_11334_),
    .Y(_11336_));
 sky130_as_sc_hs__and2_2 _42086_ (.A(_11335_),
    .B(_11336_),
    .Y(_11337_));
 sky130_as_sc_hs__or2_2 _42088_ (.A(_11309_),
    .B(_11337_),
    .Y(_11339_));
 sky130_as_sc_hs__and2_2 _42089_ (.A(_11338_),
    .B(_11339_),
    .Y(_11340_));
 sky130_as_sc_hs__or2_2 _42092_ (.A(_11340_),
    .B(_11341_),
    .Y(_11343_));
 sky130_as_sc_hs__and2_2 _42093_ (.A(_11342_),
    .B(_11343_),
    .Y(_11344_));
 sky130_as_sc_hs__and2_2 _42094_ (.A(net121),
    .B(net434),
    .Y(_11345_));
 sky130_as_sc_hs__and2_2 _42095_ (.A(net436),
    .B(net419),
    .Y(_11346_));
 sky130_as_sc_hs__and2_2 _42096_ (.A(net440),
    .B(net423),
    .Y(_11347_));
 sky130_as_sc_hs__and2_2 _42097_ (.A(_11346_),
    .B(_11347_),
    .Y(_11348_));
 sky130_as_sc_hs__nor2_2 _42098_ (.A(_11346_),
    .B(_11347_),
    .Y(_11349_));
 sky130_as_sc_hs__nor2_2 _42099_ (.A(_11348_),
    .B(_11349_),
    .Y(_11350_));
 sky130_as_sc_hs__or2_2 _42101_ (.A(_11345_),
    .B(_11350_),
    .Y(_11352_));
 sky130_as_sc_hs__or2_2 _42103_ (.A(_11184_),
    .B(_11353_),
    .Y(_11354_));
 sky130_as_sc_hs__and2_2 _42105_ (.A(_11354_),
    .B(_11355_),
    .Y(_11356_));
 sky130_as_sc_hs__or2_2 _42107_ (.A(_11344_),
    .B(_11356_),
    .Y(_11358_));
 sky130_as_sc_hs__and2_2 _42108_ (.A(_11357_),
    .B(_11358_),
    .Y(_11359_));
 sky130_as_sc_hs__or2_2 _42111_ (.A(_11359_),
    .B(_11360_),
    .Y(_11362_));
 sky130_as_sc_hs__and2_2 _42112_ (.A(_11361_),
    .B(_11362_),
    .Y(_11363_));
 sky130_as_sc_hs__and2_2 _42115_ (.A(net432),
    .B(net421),
    .Y(_11366_));
 sky130_as_sc_hs__and2_2 _42116_ (.A(net83),
    .B(net128),
    .Y(_11367_));
 sky130_as_sc_hs__or2_2 _42118_ (.A(_11181_),
    .B(_11367_),
    .Y(_11369_));
 sky130_as_sc_hs__or2_2 _42120_ (.A(_11204_),
    .B(_11370_),
    .Y(_11371_));
 sky130_as_sc_hs__and2_2 _42122_ (.A(_11371_),
    .B(_11372_),
    .Y(_11373_));
 sky130_as_sc_hs__or2_2 _42124_ (.A(_11366_),
    .B(_11373_),
    .Y(_11375_));
 sky130_as_sc_hs__and2_2 _42125_ (.A(_11374_),
    .B(_11375_),
    .Y(_11376_));
 sky130_as_sc_hs__or2_2 _42127_ (.A(_11365_),
    .B(_11376_),
    .Y(_11378_));
 sky130_as_sc_hs__and2_2 _42128_ (.A(_11377_),
    .B(_11378_),
    .Y(_11379_));
 sky130_as_sc_hs__or2_2 _42130_ (.A(_11364_),
    .B(_11379_),
    .Y(_11381_));
 sky130_as_sc_hs__and2_2 _42131_ (.A(_11380_),
    .B(_11381_),
    .Y(_11382_));
 sky130_as_sc_hs__or2_2 _42133_ (.A(_11363_),
    .B(_11382_),
    .Y(_11384_));
 sky130_as_sc_hs__and2_2 _42134_ (.A(_11383_),
    .B(_11384_),
    .Y(_11385_));
 sky130_as_sc_hs__or2_2 _42137_ (.A(_11385_),
    .B(_11386_),
    .Y(_11388_));
 sky130_as_sc_hs__and2_2 _42138_ (.A(_11387_),
    .B(_11388_),
    .Y(_11389_));
 sky130_as_sc_hs__or2_2 _42141_ (.A(_11389_),
    .B(_11390_),
    .Y(_11392_));
 sky130_as_sc_hs__and2_2 _42142_ (.A(_11391_),
    .B(_11392_),
    .Y(_11393_));
 sky130_as_sc_hs__or2_2 _42145_ (.A(_11393_),
    .B(_11394_),
    .Y(_11396_));
 sky130_as_sc_hs__and2_2 _42146_ (.A(_11395_),
    .B(_11396_),
    .Y(_11397_));
 sky130_as_sc_hs__nor2_2 _42147_ (.A(_11231_),
    .B(_11397_),
    .Y(_11398_));
 sky130_as_sc_hs__and2_2 _42148_ (.A(_11231_),
    .B(_11397_),
    .Y(_11399_));
 sky130_as_sc_hs__or2_2 _42149_ (.A(_11398_),
    .B(_11399_),
    .Y(_11400_));
 sky130_as_sc_hs__or2_2 _42151_ (.A(_11308_),
    .B(_11400_),
    .Y(_11402_));
 sky130_as_sc_hs__and2_2 _42152_ (.A(_11401_),
    .B(_11402_),
    .Y(_11403_));
 sky130_as_sc_hs__or2_2 _42155_ (.A(_11403_),
    .B(_11404_),
    .Y(_11406_));
 sky130_as_sc_hs__nand3_2 _42156_ (.A(net141),
    .B(_11405_),
    .C(_11406_),
    .Y(_11407_));
 sky130_as_sc_hs__or2_2 _42158_ (.A(_05449_),
    .B(_11408_),
    .Y(_11409_));
 sky130_as_sc_hs__nand3_2 _42160_ (.A(net138),
    .B(_11409_),
    .C(_11410_),
    .Y(_11411_));
 sky130_as_sc_hs__or2_2 _42163_ (.A(_05618_),
    .B(_11412_),
    .Y(_11414_));
 sky130_as_sc_hs__or2_2 _42166_ (.A(_05619_),
    .B(_05892_),
    .Y(_11417_));
 sky130_as_sc_hs__nand3_2 _42169_ (.A(net118),
    .B(_11416_),
    .C(_11419_),
    .Y(_11420_));
 sky130_as_sc_hs__or2_2 _42170_ (.A(\tholin_riscv.div_res[20] ),
    .B(_11267_),
    .Y(_11421_));
 sky130_as_sc_hs__and2_2 _42171_ (.A(net415),
    .B(_11421_),
    .Y(_11422_));
 sky130_as_sc_hs__or2_2 _42173_ (.A(\tholin_riscv.div_res[21] ),
    .B(_11422_),
    .Y(_11424_));
 sky130_as_sc_hs__nand3_2 _42174_ (.A(net110),
    .B(_11423_),
    .C(_11424_),
    .Y(_11425_));
 sky130_as_sc_hs__or2_2 _42175_ (.A(\tholin_riscv.div_shifter[52] ),
    .B(_11262_),
    .Y(_11426_));
 sky130_as_sc_hs__and2_2 _42176_ (.A(_21655_),
    .B(_11426_),
    .Y(_11427_));
 sky130_as_sc_hs__or2_2 _42178_ (.A(\tholin_riscv.div_shifter[53] ),
    .B(_11427_),
    .Y(_11429_));
 sky130_as_sc_hs__nand3_2 _42179_ (.A(net107),
    .B(_11428_),
    .C(_11429_),
    .Y(_11430_));
 sky130_as_sc_hs__and2_2 _42180_ (.A(_05618_),
    .B(_06538_),
    .Y(_11431_));
 sky130_as_sc_hs__or2_2 _42182_ (.A(_05616_),
    .B(_06161_),
    .Y(_11433_));
 sky130_as_sc_hs__and2_2 _42185_ (.A(_11434_),
    .B(_11435_),
    .Y(_11436_));
 sky130_as_sc_hs__and2_2 _42186_ (.A(net413),
    .B(_11436_),
    .Y(_11437_));
 sky130_as_sc_hs__nand3_2 _42187_ (.A(_11432_),
    .B(_11433_),
    .C(_11437_),
    .Y(_11438_));
 sky130_as_sc_hs__nor2_2 _42188_ (.A(_11431_),
    .B(_11438_),
    .Y(_11439_));
 sky130_as_sc_hs__nand3_2 _42189_ (.A(_11425_),
    .B(_11430_),
    .C(_11439_),
    .Y(_11440_));
 sky130_as_sc_hs__nor2_2 _42193_ (.A(_11440_),
    .B(_11443_),
    .Y(_11444_));
 sky130_as_sc_hs__and2_2 _42194_ (.A(_11420_),
    .B(_11444_),
    .Y(_11445_));
 sky130_as_sc_hs__nand3_2 _42195_ (.A(_11407_),
    .B(_11411_),
    .C(_11445_),
    .Y(_11446_));
 sky130_as_sc_hs__or2_2 _42199_ (.A(\tholin_riscv.PC[21] ),
    .B(\tholin_riscv.Iimm[1] ),
    .Y(_11450_));
 sky130_as_sc_hs__or2_2 _42201_ (.A(_11448_),
    .B(_11451_),
    .Y(_11452_));
 sky130_as_sc_hs__nand3_2 _42203_ (.A(net117),
    .B(_11452_),
    .C(_11453_),
    .Y(_11454_));
 sky130_as_sc_hs__and2_2 _42204_ (.A(\tholin_riscv.PC[21] ),
    .B(_11286_),
    .Y(_11455_));
 sky130_as_sc_hs__nor2_2 _42205_ (.A(\tholin_riscv.PC[21] ),
    .B(_11286_),
    .Y(_11456_));
 sky130_as_sc_hs__or2_2 _42206_ (.A(_11455_),
    .B(_11456_),
    .Y(_11457_));
 sky130_as_sc_hs__nand3_2 _42209_ (.A(_11454_),
    .B(_11458_),
    .C(_11459_),
    .Y(_11460_));
 sky130_as_sc_hs__nand3_2 _42211_ (.A(_21546_),
    .B(_11446_),
    .C(_11461_),
    .Y(_11462_));
 sky130_as_sc_hs__and2_2 _42216_ (.A(\tholin_riscv.Iimm[2] ),
    .B(\tholin_riscv.io_size[1] ),
    .Y(_11466_));
 sky130_as_sc_hs__or2_2 _42217_ (.A(_10352_),
    .B(_11466_),
    .Y(_11467_));
 sky130_as_sc_hs__and2_2 _42219_ (.A(net427),
    .B(net425),
    .Y(_11469_));
 sky130_as_sc_hs__and2_2 _42220_ (.A(net83),
    .B(net418),
    .Y(_11470_));
 sky130_as_sc_hs__and2_2 _42221_ (.A(net120),
    .B(net433),
    .Y(_11471_));
 sky130_as_sc_hs__or2_2 _42223_ (.A(_11470_),
    .B(_11471_),
    .Y(_11473_));
 sky130_as_sc_hs__and2_2 _42224_ (.A(_11472_),
    .B(_11473_),
    .Y(_11474_));
 sky130_as_sc_hs__and2_2 _42225_ (.A(net457),
    .B(net423),
    .Y(_11475_));
 sky130_as_sc_hs__or2_2 _42227_ (.A(_11474_),
    .B(_11475_),
    .Y(_11477_));
 sky130_as_sc_hs__and2_2 _42228_ (.A(_11476_),
    .B(_11477_),
    .Y(_11478_));
 sky130_as_sc_hs__or2_2 _42231_ (.A(_11478_),
    .B(_11479_),
    .Y(_11481_));
 sky130_as_sc_hs__and2_2 _42232_ (.A(_11480_),
    .B(_11481_),
    .Y(_11482_));
 sky130_as_sc_hs__or2_2 _42235_ (.A(_11482_),
    .B(_11483_),
    .Y(_11485_));
 sky130_as_sc_hs__and2_2 _42236_ (.A(_11484_),
    .B(_11485_),
    .Y(_11486_));
 sky130_as_sc_hs__or2_2 _42239_ (.A(_11486_),
    .B(_11487_),
    .Y(_11489_));
 sky130_as_sc_hs__and2_2 _42240_ (.A(_11488_),
    .B(_11489_),
    .Y(_11490_));
 sky130_as_sc_hs__or2_2 _42242_ (.A(_11469_),
    .B(_11490_),
    .Y(_11492_));
 sky130_as_sc_hs__and2_2 _42243_ (.A(_11491_),
    .B(_11492_),
    .Y(_11493_));
 sky130_as_sc_hs__or2_2 _42246_ (.A(_11493_),
    .B(_11494_),
    .Y(_11496_));
 sky130_as_sc_hs__and2_2 _42247_ (.A(_11495_),
    .B(_11496_),
    .Y(_11497_));
 sky130_as_sc_hs__and2_2 _42248_ (.A(net122),
    .B(net434),
    .Y(_11498_));
 sky130_as_sc_hs__and2_2 _42249_ (.A(net436),
    .B(net75),
    .Y(_11499_));
 sky130_as_sc_hs__and2_2 _42250_ (.A(net440),
    .B(net419),
    .Y(_11500_));
 sky130_as_sc_hs__and2_2 _42251_ (.A(_11499_),
    .B(_11500_),
    .Y(_11501_));
 sky130_as_sc_hs__nor2_2 _42252_ (.A(_11499_),
    .B(_11500_),
    .Y(_11502_));
 sky130_as_sc_hs__nor2_2 _42253_ (.A(_11501_),
    .B(_11502_),
    .Y(_11503_));
 sky130_as_sc_hs__or2_2 _42255_ (.A(_11498_),
    .B(_11503_),
    .Y(_11505_));
 sky130_as_sc_hs__or2_2 _42257_ (.A(_11351_),
    .B(_11506_),
    .Y(_11507_));
 sky130_as_sc_hs__and2_2 _42259_ (.A(_11507_),
    .B(_11508_),
    .Y(_11509_));
 sky130_as_sc_hs__or2_2 _42261_ (.A(_11497_),
    .B(_11509_),
    .Y(_11511_));
 sky130_as_sc_hs__and2_2 _42262_ (.A(_11510_),
    .B(_11511_),
    .Y(_11512_));
 sky130_as_sc_hs__or2_2 _42265_ (.A(_11512_),
    .B(_11513_),
    .Y(_11515_));
 sky130_as_sc_hs__and2_2 _42266_ (.A(_11514_),
    .B(_11515_),
    .Y(_11516_));
 sky130_as_sc_hs__and2_2 _42268_ (.A(net430),
    .B(net421),
    .Y(_11518_));
 sky130_as_sc_hs__and2_2 _42269_ (.A(net431),
    .B(net128),
    .Y(_11519_));
 sky130_as_sc_hs__or2_2 _42271_ (.A(_11348_),
    .B(_11519_),
    .Y(_11521_));
 sky130_as_sc_hs__or2_2 _42273_ (.A(_11368_),
    .B(_11522_),
    .Y(_11523_));
 sky130_as_sc_hs__and2_2 _42275_ (.A(_11523_),
    .B(_11524_),
    .Y(_11525_));
 sky130_as_sc_hs__or2_2 _42277_ (.A(_11518_),
    .B(_11525_),
    .Y(_11527_));
 sky130_as_sc_hs__or2_2 _42279_ (.A(_11354_),
    .B(_11528_),
    .Y(_11529_));
 sky130_as_sc_hs__and2_2 _42281_ (.A(_11529_),
    .B(_11530_),
    .Y(_11531_));
 sky130_as_sc_hs__or2_2 _42283_ (.A(_11517_),
    .B(_11531_),
    .Y(_11533_));
 sky130_as_sc_hs__and2_2 _42284_ (.A(_11532_),
    .B(_11533_),
    .Y(_11534_));
 sky130_as_sc_hs__or2_2 _42286_ (.A(_11516_),
    .B(_11534_),
    .Y(_11536_));
 sky130_as_sc_hs__and2_2 _42287_ (.A(_11535_),
    .B(_11536_),
    .Y(_11537_));
 sky130_as_sc_hs__or2_2 _42290_ (.A(_11537_),
    .B(_11538_),
    .Y(_11540_));
 sky130_as_sc_hs__and2_2 _42291_ (.A(_11539_),
    .B(_11540_),
    .Y(_11541_));
 sky130_as_sc_hs__or2_2 _42294_ (.A(_11541_),
    .B(_11542_),
    .Y(_11544_));
 sky130_as_sc_hs__and2_2 _42295_ (.A(_11543_),
    .B(_11544_),
    .Y(_11545_));
 sky130_as_sc_hs__or2_2 _42298_ (.A(_11545_),
    .B(_11546_),
    .Y(_11548_));
 sky130_as_sc_hs__or2_2 _42300_ (.A(_11395_),
    .B(_11549_),
    .Y(_11550_));
 sky130_as_sc_hs__and2_2 _42302_ (.A(_11550_),
    .B(_11551_),
    .Y(_11552_));
 sky130_as_sc_hs__and2_2 _42305_ (.A(_11236_),
    .B(_11400_),
    .Y(_11555_));
 sky130_as_sc_hs__or2_2 _42309_ (.A(_11552_),
    .B(_11557_),
    .Y(_11559_));
 sky130_as_sc_hs__and2_2 _42311_ (.A(_11240_),
    .B(_11403_),
    .Y(_11561_));
 sky130_as_sc_hs__or2_2 _42312_ (.A(_05505_),
    .B(_11561_),
    .Y(_11562_));
 sky130_as_sc_hs__and2_2 _42313_ (.A(_11243_),
    .B(_11562_),
    .Y(_11563_));
 sky130_as_sc_hs__or2_2 _42314_ (.A(_11560_),
    .B(_11563_),
    .Y(_11564_));
 sky130_as_sc_hs__nand3_2 _42316_ (.A(net141),
    .B(_11564_),
    .C(_11565_),
    .Y(_11566_));
 sky130_as_sc_hs__or2_2 _42318_ (.A(_05374_),
    .B(_11567_),
    .Y(_11568_));
 sky130_as_sc_hs__nand3_2 _42320_ (.A(net138),
    .B(_11568_),
    .C(_11569_),
    .Y(_11570_));
 sky130_as_sc_hs__nor2_2 _42322_ (.A(_05606_),
    .B(_06161_),
    .Y(_11572_));
 sky130_as_sc_hs__and2_2 _42324_ (.A(\tholin_riscv.div_res[22] ),
    .B(_06564_),
    .Y(_11574_));
 sky130_as_sc_hs__nor2_2 _42326_ (.A(net118),
    .B(_11574_),
    .Y(_11576_));
 sky130_as_sc_hs__nand3_2 _42327_ (.A(_11573_),
    .B(_11575_),
    .C(_11576_),
    .Y(_11577_));
 sky130_as_sc_hs__nor2_2 _42328_ (.A(_11572_),
    .B(_11577_),
    .Y(_11578_));
 sky130_as_sc_hs__nand3_2 _42330_ (.A(_11571_),
    .B(_11578_),
    .C(_11579_),
    .Y(_11580_));
 sky130_as_sc_hs__or2_2 _42331_ (.A(\tholin_riscv.div_res[21] ),
    .B(_11421_),
    .Y(_11581_));
 sky130_as_sc_hs__and2_2 _42332_ (.A(net414),
    .B(_11581_),
    .Y(_11582_));
 sky130_as_sc_hs__or2_2 _42334_ (.A(\tholin_riscv.div_res[22] ),
    .B(_11582_),
    .Y(_11584_));
 sky130_as_sc_hs__nand3_2 _42335_ (.A(net111),
    .B(_11583_),
    .C(_11584_),
    .Y(_11585_));
 sky130_as_sc_hs__or2_2 _42336_ (.A(\tholin_riscv.div_shifter[53] ),
    .B(_11426_),
    .Y(_11586_));
 sky130_as_sc_hs__and2_2 _42337_ (.A(_21655_),
    .B(_11586_),
    .Y(_11587_));
 sky130_as_sc_hs__or2_2 _42339_ (.A(\tholin_riscv.div_shifter[54] ),
    .B(_11587_),
    .Y(_11589_));
 sky130_as_sc_hs__nand3_2 _42340_ (.A(net107),
    .B(_11588_),
    .C(_11589_),
    .Y(_11590_));
 sky130_as_sc_hs__nand3_2 _42342_ (.A(_11585_),
    .B(_11590_),
    .C(_11591_),
    .Y(_11592_));
 sky130_as_sc_hs__nor2_2 _42343_ (.A(_11580_),
    .B(_11592_),
    .Y(_11593_));
 sky130_as_sc_hs__nand3_2 _42344_ (.A(_11566_),
    .B(_11570_),
    .C(_11593_),
    .Y(_11594_));
 sky130_as_sc_hs__or2_2 _42345_ (.A(_05609_),
    .B(_05894_),
    .Y(_11595_));
 sky130_as_sc_hs__or2_2 _42348_ (.A(_05608_),
    .B(_11596_),
    .Y(_11598_));
 sky130_as_sc_hs__nand3_2 _42350_ (.A(_05895_),
    .B(_06527_),
    .C(_11595_),
    .Y(_11600_));
 sky130_as_sc_hs__or2_2 _42351_ (.A(_06527_),
    .B(_11599_),
    .Y(_11601_));
 sky130_as_sc_hs__nand3_2 _42352_ (.A(net119),
    .B(_11600_),
    .C(_11601_),
    .Y(_11602_));
 sky130_as_sc_hs__or2_2 _42358_ (.A(\tholin_riscv.PC[22] ),
    .B(\tholin_riscv.Iimm[2] ),
    .Y(_11608_));
 sky130_as_sc_hs__or2_2 _42360_ (.A(_11606_),
    .B(_11609_),
    .Y(_11610_));
 sky130_as_sc_hs__nand3_2 _42362_ (.A(net117),
    .B(_11610_),
    .C(_11611_),
    .Y(_11612_));
 sky130_as_sc_hs__or2_2 _42363_ (.A(\tholin_riscv.Iimm[2] ),
    .B(_21590_),
    .Y(_11613_));
 sky130_as_sc_hs__and2_2 _42364_ (.A(\tholin_riscv.PC[22] ),
    .B(_11455_),
    .Y(_11614_));
 sky130_as_sc_hs__nor2_2 _42365_ (.A(\tholin_riscv.PC[22] ),
    .B(_11455_),
    .Y(_11615_));
 sky130_as_sc_hs__or2_2 _42366_ (.A(_11614_),
    .B(_11615_),
    .Y(_11616_));
 sky130_as_sc_hs__nand3_2 _42368_ (.A(_11612_),
    .B(_11613_),
    .C(_11617_),
    .Y(_11618_));
 sky130_as_sc_hs__nand3_2 _42370_ (.A(_21546_),
    .B(_11604_),
    .C(_11619_),
    .Y(_11620_));
 sky130_as_sc_hs__and2_2 _42375_ (.A(\tholin_riscv.Iimm[3] ),
    .B(net371),
    .Y(_11624_));
 sky130_as_sc_hs__or2_2 _42376_ (.A(_10352_),
    .B(_11624_),
    .Y(_11625_));
 sky130_as_sc_hs__and2_2 _42378_ (.A(_11550_),
    .B(_11558_),
    .Y(_11627_));
 sky130_as_sc_hs__and2_2 _42379_ (.A(net121),
    .B(net425),
    .Y(_11628_));
 sky130_as_sc_hs__and2_2 _42380_ (.A(net431),
    .B(net418),
    .Y(_11629_));
 sky130_as_sc_hs__and2_2 _42381_ (.A(net122),
    .B(net433),
    .Y(_11630_));
 sky130_as_sc_hs__or2_2 _42383_ (.A(_11629_),
    .B(_11630_),
    .Y(_11632_));
 sky130_as_sc_hs__and2_2 _42384_ (.A(_11631_),
    .B(_11632_),
    .Y(_11633_));
 sky130_as_sc_hs__and2_2 _42385_ (.A(net457),
    .B(net419),
    .Y(_11634_));
 sky130_as_sc_hs__or2_2 _42387_ (.A(_11633_),
    .B(_11634_),
    .Y(_11636_));
 sky130_as_sc_hs__and2_2 _42388_ (.A(_11635_),
    .B(_11636_),
    .Y(_11637_));
 sky130_as_sc_hs__or2_2 _42391_ (.A(_11637_),
    .B(_11638_),
    .Y(_11640_));
 sky130_as_sc_hs__or2_2 _42394_ (.A(_11641_),
    .B(_11642_),
    .Y(_11643_));
 sky130_as_sc_hs__or2_2 _42398_ (.A(_11628_),
    .B(_11645_),
    .Y(_11647_));
 sky130_as_sc_hs__and2_2 _42399_ (.A(_11646_),
    .B(_11647_),
    .Y(_11648_));
 sky130_as_sc_hs__or2_2 _42402_ (.A(_11648_),
    .B(_11649_),
    .Y(_11651_));
 sky130_as_sc_hs__and2_2 _42403_ (.A(_11650_),
    .B(_11651_),
    .Y(_11652_));
 sky130_as_sc_hs__and2_2 _42404_ (.A(net440),
    .B(net74),
    .Y(_11653_));
 sky130_as_sc_hs__and2_2 _42405_ (.A(net434),
    .B(net423),
    .Y(_11654_));
 sky130_as_sc_hs__or2_2 _42407_ (.A(_11653_),
    .B(_11654_),
    .Y(_11656_));
 sky130_as_sc_hs__or2_2 _42409_ (.A(_11504_),
    .B(_11657_),
    .Y(_11658_));
 sky130_as_sc_hs__and2_2 _42411_ (.A(_11658_),
    .B(_11659_),
    .Y(_11660_));
 sky130_as_sc_hs__or2_2 _42413_ (.A(_11652_),
    .B(_11660_),
    .Y(_11662_));
 sky130_as_sc_hs__and2_2 _42414_ (.A(_11661_),
    .B(_11662_),
    .Y(_11663_));
 sky130_as_sc_hs__or2_2 _42417_ (.A(_11663_),
    .B(_11664_),
    .Y(_11666_));
 sky130_as_sc_hs__and2_2 _42418_ (.A(_11665_),
    .B(_11666_),
    .Y(_11667_));
 sky130_as_sc_hs__and2_2 _42420_ (.A(net428),
    .B(net422),
    .Y(_11669_));
 sky130_as_sc_hs__and2_2 _42421_ (.A(net429),
    .B(net128),
    .Y(_11670_));
 sky130_as_sc_hs__or2_2 _42423_ (.A(_11501_),
    .B(_11670_),
    .Y(_11672_));
 sky130_as_sc_hs__or2_2 _42425_ (.A(_11520_),
    .B(_11673_),
    .Y(_11674_));
 sky130_as_sc_hs__and2_2 _42427_ (.A(_11674_),
    .B(_11675_),
    .Y(_11676_));
 sky130_as_sc_hs__or2_2 _42429_ (.A(_11669_),
    .B(_11676_),
    .Y(_11678_));
 sky130_as_sc_hs__or2_2 _42431_ (.A(_11507_),
    .B(_11679_),
    .Y(_11680_));
 sky130_as_sc_hs__and2_2 _42433_ (.A(_11680_),
    .B(_11681_),
    .Y(_11682_));
 sky130_as_sc_hs__or2_2 _42435_ (.A(_11668_),
    .B(_11682_),
    .Y(_11684_));
 sky130_as_sc_hs__and2_2 _42436_ (.A(_11683_),
    .B(_11684_),
    .Y(_11685_));
 sky130_as_sc_hs__or2_2 _42438_ (.A(_11667_),
    .B(_11685_),
    .Y(_11687_));
 sky130_as_sc_hs__and2_2 _42439_ (.A(_11686_),
    .B(_11687_),
    .Y(_11688_));
 sky130_as_sc_hs__or2_2 _42442_ (.A(_11688_),
    .B(_11689_),
    .Y(_11691_));
 sky130_as_sc_hs__and2_2 _42443_ (.A(_11690_),
    .B(_11691_),
    .Y(_11692_));
 sky130_as_sc_hs__or2_2 _42446_ (.A(_11692_),
    .B(_11693_),
    .Y(_11695_));
 sky130_as_sc_hs__and2_2 _42447_ (.A(_11694_),
    .B(_11695_),
    .Y(_11696_));
 sky130_as_sc_hs__or2_2 _42450_ (.A(_11696_),
    .B(_11697_),
    .Y(_11699_));
 sky130_as_sc_hs__and2_2 _42451_ (.A(_11698_),
    .B(_11699_),
    .Y(_11700_));
 sky130_as_sc_hs__or2_2 _42452_ (.A(_11547_),
    .B(_11700_),
    .Y(_11701_));
 sky130_as_sc_hs__or2_2 _42456_ (.A(_11627_),
    .B(_11703_),
    .Y(_11705_));
 sky130_as_sc_hs__and2_2 _42457_ (.A(_11704_),
    .B(_11705_),
    .Y(_11706_));
 sky130_as_sc_hs__and2_2 _42458_ (.A(_11241_),
    .B(_11560_),
    .Y(_11707_));
 sky130_as_sc_hs__and2_2 _42459_ (.A(_11561_),
    .B(_11707_),
    .Y(_11708_));
 sky130_as_sc_hs__and2_2 _42460_ (.A(_10503_),
    .B(_11708_),
    .Y(_11709_));
 sky130_as_sc_hs__or2_2 _42461_ (.A(_05505_),
    .B(_11709_),
    .Y(_11710_));
 sky130_as_sc_hs__or2_2 _42463_ (.A(_11706_),
    .B(_11710_),
    .Y(_11712_));
 sky130_as_sc_hs__nand3_2 _42464_ (.A(net141),
    .B(_11711_),
    .C(_11712_),
    .Y(_11713_));
 sky130_as_sc_hs__and2_2 _42465_ (.A(_05452_),
    .B(_05504_),
    .Y(_11714_));
 sky130_as_sc_hs__or2_2 _42467_ (.A(_05456_),
    .B(_11714_),
    .Y(_11716_));
 sky130_as_sc_hs__nand3_2 _42468_ (.A(net138),
    .B(_11715_),
    .C(_11716_),
    .Y(_11717_));
 sky130_as_sc_hs__or2_2 _42471_ (.A(_05598_),
    .B(_11718_),
    .Y(_11720_));
 sky130_as_sc_hs__or2_2 _42474_ (.A(_05599_),
    .B(_05896_),
    .Y(_11723_));
 sky130_as_sc_hs__nand3_2 _42477_ (.A(net118),
    .B(_11722_),
    .C(_11725_),
    .Y(_11726_));
 sky130_as_sc_hs__and2_2 _42478_ (.A(net140),
    .B(_08663_),
    .Y(_11727_));
 sky130_as_sc_hs__and2_2 _42481_ (.A(_05597_),
    .B(_06157_),
    .Y(_11730_));
 sky130_as_sc_hs__or2_2 _42482_ (.A(_05596_),
    .B(_06161_),
    .Y(_11731_));
 sky130_as_sc_hs__nand3_2 _42485_ (.A(net413),
    .B(_11732_),
    .C(_11733_),
    .Y(_11734_));
 sky130_as_sc_hs__nor2_2 _42486_ (.A(_11730_),
    .B(_11734_),
    .Y(_11735_));
 sky130_as_sc_hs__nand3_2 _42487_ (.A(_11729_),
    .B(_11731_),
    .C(_11735_),
    .Y(_11736_));
 sky130_as_sc_hs__nor2_2 _42488_ (.A(_11727_),
    .B(_11736_),
    .Y(_11737_));
 sky130_as_sc_hs__and2_2 _42489_ (.A(_11728_),
    .B(_11737_),
    .Y(_11738_));
 sky130_as_sc_hs__or2_2 _42490_ (.A(\tholin_riscv.div_shifter[54] ),
    .B(_11586_),
    .Y(_11739_));
 sky130_as_sc_hs__and2_2 _42491_ (.A(_21655_),
    .B(_11739_),
    .Y(_11740_));
 sky130_as_sc_hs__or2_2 _42493_ (.A(\tholin_riscv.div_shifter[55] ),
    .B(_11740_),
    .Y(_11742_));
 sky130_as_sc_hs__nand3_2 _42494_ (.A(net107),
    .B(_11741_),
    .C(_11742_),
    .Y(_11743_));
 sky130_as_sc_hs__or2_2 _42495_ (.A(\tholin_riscv.div_res[22] ),
    .B(_11581_),
    .Y(_11744_));
 sky130_as_sc_hs__and2_2 _42496_ (.A(net414),
    .B(_11744_),
    .Y(_11745_));
 sky130_as_sc_hs__or2_2 _42498_ (.A(\tholin_riscv.div_res[23] ),
    .B(_11745_),
    .Y(_11747_));
 sky130_as_sc_hs__nand3_2 _42499_ (.A(net110),
    .B(_11746_),
    .C(_11747_),
    .Y(_11748_));
 sky130_as_sc_hs__and2_2 _42500_ (.A(_11743_),
    .B(_11748_),
    .Y(_11749_));
 sky130_as_sc_hs__and2_2 _42501_ (.A(_11738_),
    .B(_11749_),
    .Y(_11750_));
 sky130_as_sc_hs__and2_2 _42502_ (.A(_11726_),
    .B(_11750_),
    .Y(_11751_));
 sky130_as_sc_hs__nand3_2 _42503_ (.A(_11713_),
    .B(_11717_),
    .C(_11751_),
    .Y(_11752_));
 sky130_as_sc_hs__or2_2 _42505_ (.A(\tholin_riscv.PC[23] ),
    .B(\tholin_riscv.Iimm[3] ),
    .Y(_11754_));
 sky130_as_sc_hs__and2_2 _42508_ (.A(_11607_),
    .B(_11756_),
    .Y(_11757_));
 sky130_as_sc_hs__or2_2 _42510_ (.A(_11755_),
    .B(_11757_),
    .Y(_11759_));
 sky130_as_sc_hs__nand3_2 _42511_ (.A(net117),
    .B(_11758_),
    .C(_11759_),
    .Y(_11760_));
 sky130_as_sc_hs__and2_2 _42512_ (.A(\tholin_riscv.PC[23] ),
    .B(_11614_),
    .Y(_11761_));
 sky130_as_sc_hs__nor2_2 _42513_ (.A(\tholin_riscv.PC[23] ),
    .B(_11614_),
    .Y(_11762_));
 sky130_as_sc_hs__nor2_2 _42514_ (.A(_11761_),
    .B(_11762_),
    .Y(_11763_));
 sky130_as_sc_hs__inv_2 _42515_ (.Y(_11764_),
    .A(_11763_));
 sky130_as_sc_hs__and2_2 _42518_ (.A(_21569_),
    .B(_11766_),
    .Y(_11767_));
 sky130_as_sc_hs__nand3_2 _42519_ (.A(_11760_),
    .B(_11765_),
    .C(_11767_),
    .Y(_11768_));
 sky130_as_sc_hs__nand3_2 _42520_ (.A(_21546_),
    .B(_11752_),
    .C(_11768_),
    .Y(_11769_));
 sky130_as_sc_hs__and2_2 _42525_ (.A(\tholin_riscv.Iimm[4] ),
    .B(\tholin_riscv.io_size[1] ),
    .Y(_11773_));
 sky130_as_sc_hs__or2_2 _42526_ (.A(_10352_),
    .B(_11773_),
    .Y(_11774_));
 sky130_as_sc_hs__and2_2 _42528_ (.A(_11552_),
    .B(_11703_),
    .Y(_11776_));
 sky130_as_sc_hs__nand3_2 _42529_ (.A(_11136_),
    .B(_11555_),
    .C(_11776_),
    .Y(_11777_));
 sky130_as_sc_hs__nand2b_2 _42530_ (.B(_11776_),
    .Y(_11778_),
    .A(_11554_));
 sky130_as_sc_hs__nand3_2 _42533_ (.A(_11777_),
    .B(_11778_),
    .C(_11780_),
    .Y(_11781_));
 sky130_as_sc_hs__and2_2 _42534_ (.A(net122),
    .B(net425),
    .Y(_11782_));
 sky130_as_sc_hs__and2_2 _42535_ (.A(net429),
    .B(net418),
    .Y(_11783_));
 sky130_as_sc_hs__and2_2 _42536_ (.A(net433),
    .B(net423),
    .Y(_11784_));
 sky130_as_sc_hs__or2_2 _42538_ (.A(_11783_),
    .B(_11784_),
    .Y(_11786_));
 sky130_as_sc_hs__and2_2 _42539_ (.A(_11785_),
    .B(_11786_),
    .Y(_11787_));
 sky130_as_sc_hs__and2_2 _42540_ (.A(net457),
    .B(net74),
    .Y(_11788_));
 sky130_as_sc_hs__or2_2 _42542_ (.A(_11787_),
    .B(_11788_),
    .Y(_11790_));
 sky130_as_sc_hs__and2_2 _42543_ (.A(_11789_),
    .B(_11790_),
    .Y(_11791_));
 sky130_as_sc_hs__and2_2 _42545_ (.A(_11791_),
    .B(_11792_),
    .Y(_11793_));
 sky130_as_sc_hs__nor2_2 _42546_ (.A(_11791_),
    .B(_11792_),
    .Y(_11794_));
 sky130_as_sc_hs__nor2_2 _42547_ (.A(_11793_),
    .B(_11794_),
    .Y(_11795_));
 sky130_as_sc_hs__or2_2 _42548_ (.A(_11480_),
    .B(_11641_),
    .Y(_11796_));
 sky130_as_sc_hs__inv_2 _42549_ (.Y(_11797_),
    .A(_11796_));
 sky130_as_sc_hs__and2_2 _42550_ (.A(_11639_),
    .B(_11796_),
    .Y(_11798_));
 sky130_as_sc_hs__or2_2 _42552_ (.A(_11795_),
    .B(_11798_),
    .Y(_11800_));
 sky130_as_sc_hs__or2_2 _42555_ (.A(_11782_),
    .B(_11801_),
    .Y(_11803_));
 sky130_as_sc_hs__and2_2 _42556_ (.A(_11802_),
    .B(_11803_),
    .Y(_11804_));
 sky130_as_sc_hs__or2_2 _42557_ (.A(_11484_),
    .B(_11641_),
    .Y(_11805_));
 sky130_as_sc_hs__or2_2 _42560_ (.A(_11804_),
    .B(_11806_),
    .Y(_11808_));
 sky130_as_sc_hs__and2_2 _42561_ (.A(_11807_),
    .B(_11808_),
    .Y(_11809_));
 sky130_as_sc_hs__nand3_2 _42562_ (.A(net419),
    .B(_11653_),
    .C(_11654_),
    .Y(_11810_));
 sky130_as_sc_hs__and2_2 _42565_ (.A(_11810_),
    .B(_11812_),
    .Y(_11813_));
 sky130_as_sc_hs__or2_2 _42567_ (.A(_11809_),
    .B(_11813_),
    .Y(_11815_));
 sky130_as_sc_hs__and2_2 _42568_ (.A(_11814_),
    .B(_11815_),
    .Y(_11816_));
 sky130_as_sc_hs__or2_2 _42571_ (.A(_11816_),
    .B(_11817_),
    .Y(_11819_));
 sky130_as_sc_hs__and2_2 _42572_ (.A(_11818_),
    .B(_11819_),
    .Y(_11820_));
 sky130_as_sc_hs__and2_2 _42574_ (.A(net121),
    .B(net421),
    .Y(_11822_));
 sky130_as_sc_hs__nand3_2 _42575_ (.A(net428),
    .B(_11501_),
    .C(_11670_),
    .Y(_11823_));
 sky130_as_sc_hs__and2_2 _42578_ (.A(_11823_),
    .B(_11825_),
    .Y(_11826_));
 sky130_as_sc_hs__or2_2 _42580_ (.A(_11822_),
    .B(_11826_),
    .Y(_11828_));
 sky130_as_sc_hs__or2_2 _42582_ (.A(_11658_),
    .B(_11829_),
    .Y(_11830_));
 sky130_as_sc_hs__and2_2 _42584_ (.A(_11830_),
    .B(_11831_),
    .Y(_11832_));
 sky130_as_sc_hs__or2_2 _42586_ (.A(_11821_),
    .B(_11832_),
    .Y(_11834_));
 sky130_as_sc_hs__and2_2 _42587_ (.A(_11833_),
    .B(_11834_),
    .Y(_11835_));
 sky130_as_sc_hs__or2_2 _42589_ (.A(_11820_),
    .B(_11835_),
    .Y(_11837_));
 sky130_as_sc_hs__and2_2 _42590_ (.A(_11836_),
    .B(_11837_),
    .Y(_11838_));
 sky130_as_sc_hs__or2_2 _42593_ (.A(_11838_),
    .B(_11839_),
    .Y(_11841_));
 sky130_as_sc_hs__and2_2 _42594_ (.A(_11840_),
    .B(_11841_),
    .Y(_11842_));
 sky130_as_sc_hs__or2_2 _42597_ (.A(_11842_),
    .B(_11843_),
    .Y(_11845_));
 sky130_as_sc_hs__and2_2 _42598_ (.A(_11844_),
    .B(_11845_),
    .Y(_11846_));
 sky130_as_sc_hs__or2_2 _42601_ (.A(_11846_),
    .B(_11847_),
    .Y(_11849_));
 sky130_as_sc_hs__or2_2 _42603_ (.A(_11698_),
    .B(_11850_),
    .Y(_11851_));
 sky130_as_sc_hs__and2_2 _42605_ (.A(_11851_),
    .B(_11852_),
    .Y(_11853_));
 sky130_as_sc_hs__or2_2 _42607_ (.A(_11781_),
    .B(_11853_),
    .Y(_11855_));
 sky130_as_sc_hs__and2_2 _42609_ (.A(_11706_),
    .B(_11709_),
    .Y(_11857_));
 sky130_as_sc_hs__or2_2 _42610_ (.A(_05505_),
    .B(_11857_),
    .Y(_11858_));
 sky130_as_sc_hs__or2_2 _42611_ (.A(_11856_),
    .B(_11858_),
    .Y(_11859_));
 sky130_as_sc_hs__nand3_2 _42613_ (.A(net141),
    .B(_11859_),
    .C(_11860_),
    .Y(_11861_));
 sky130_as_sc_hs__or2_2 _42614_ (.A(_05457_),
    .B(_05505_),
    .Y(_11862_));
 sky130_as_sc_hs__or2_2 _42616_ (.A(_05470_),
    .B(_11862_),
    .Y(_11864_));
 sky130_as_sc_hs__nand3_2 _42617_ (.A(net138),
    .B(_11863_),
    .C(_11864_),
    .Y(_11865_));
 sky130_as_sc_hs__or2_2 _42619_ (.A(_05901_),
    .B(_11866_),
    .Y(_11867_));
 sky130_as_sc_hs__and2_2 _42621_ (.A(_11867_),
    .B(_11868_),
    .Y(_11869_));
 sky130_as_sc_hs__or2_2 _42623_ (.A(_05898_),
    .B(_05901_),
    .Y(_11871_));
 sky130_as_sc_hs__nand3_2 _42626_ (.A(net118),
    .B(_11870_),
    .C(_11873_),
    .Y(_11874_));
 sky130_as_sc_hs__or2_2 _42627_ (.A(\tholin_riscv.div_res[23] ),
    .B(_11744_),
    .Y(_11875_));
 sky130_as_sc_hs__and2_2 _42628_ (.A(net414),
    .B(_11875_),
    .Y(_11876_));
 sky130_as_sc_hs__or2_2 _42629_ (.A(\tholin_riscv.div_res[24] ),
    .B(_11876_),
    .Y(_11877_));
 sky130_as_sc_hs__nand3_2 _42631_ (.A(net110),
    .B(_11877_),
    .C(_11878_),
    .Y(_11879_));
 sky130_as_sc_hs__or2_2 _42632_ (.A(\tholin_riscv.div_shifter[55] ),
    .B(_11739_),
    .Y(_11880_));
 sky130_as_sc_hs__and2_2 _42633_ (.A(_21655_),
    .B(_11880_),
    .Y(_11881_));
 sky130_as_sc_hs__or2_2 _42634_ (.A(\tholin_riscv.div_shifter[56] ),
    .B(_11881_),
    .Y(_11882_));
 sky130_as_sc_hs__nand3_2 _42636_ (.A(net107),
    .B(_11882_),
    .C(_11883_),
    .Y(_11884_));
 sky130_as_sc_hs__and2_2 _42637_ (.A(net140),
    .B(_08388_),
    .Y(_11885_));
 sky130_as_sc_hs__nor2_2 _42642_ (.A(_05899_),
    .B(_06161_),
    .Y(_11890_));
 sky130_as_sc_hs__nand3_2 _42645_ (.A(net412),
    .B(_11891_),
    .C(_11892_),
    .Y(_11893_));
 sky130_as_sc_hs__nor2_2 _42646_ (.A(_11890_),
    .B(_11893_),
    .Y(_11894_));
 sky130_as_sc_hs__nand3_2 _42647_ (.A(_11886_),
    .B(_11889_),
    .C(_11894_),
    .Y(_11895_));
 sky130_as_sc_hs__nor2_2 _42648_ (.A(_11885_),
    .B(_11895_),
    .Y(_11896_));
 sky130_as_sc_hs__and2_2 _42649_ (.A(_11884_),
    .B(_11896_),
    .Y(_11897_));
 sky130_as_sc_hs__and2_2 _42650_ (.A(_11879_),
    .B(_11897_),
    .Y(_11898_));
 sky130_as_sc_hs__and2_2 _42651_ (.A(_11874_),
    .B(_11898_),
    .Y(_11899_));
 sky130_as_sc_hs__nand3_2 _42652_ (.A(_11861_),
    .B(_11865_),
    .C(_11899_),
    .Y(_11900_));
 sky130_as_sc_hs__or2_2 _42655_ (.A(\tholin_riscv.PC[24] ),
    .B(\tholin_riscv.Iimm[4] ),
    .Y(_11903_));
 sky130_as_sc_hs__or2_2 _42657_ (.A(_11901_),
    .B(_11904_),
    .Y(_11905_));
 sky130_as_sc_hs__nand3_2 _42659_ (.A(net117),
    .B(_11905_),
    .C(_11906_),
    .Y(_11907_));
 sky130_as_sc_hs__and2_2 _42661_ (.A(\tholin_riscv.PC[24] ),
    .B(_11761_),
    .Y(_11909_));
 sky130_as_sc_hs__nor2_2 _42662_ (.A(\tholin_riscv.PC[24] ),
    .B(_11761_),
    .Y(_11910_));
 sky130_as_sc_hs__or2_2 _42663_ (.A(_11909_),
    .B(_11910_),
    .Y(_11911_));
 sky130_as_sc_hs__nand3_2 _42665_ (.A(_11907_),
    .B(_11908_),
    .C(_11912_),
    .Y(_11913_));
 sky130_as_sc_hs__nand3_2 _42667_ (.A(_21546_),
    .B(_11900_),
    .C(_11914_),
    .Y(_11915_));
 sky130_as_sc_hs__and2_2 _42672_ (.A(\tholin_riscv.Bimm[5] ),
    .B(net371),
    .Y(_11919_));
 sky130_as_sc_hs__or2_2 _42673_ (.A(_10352_),
    .B(_11919_),
    .Y(_11920_));
 sky130_as_sc_hs__and2_2 _42675_ (.A(_11851_),
    .B(_11854_),
    .Y(_11922_));
 sky130_as_sc_hs__and2_2 _42676_ (.A(net434),
    .B(net74),
    .Y(_11923_));
 sky130_as_sc_hs__and2_2 _42677_ (.A(net425),
    .B(net423),
    .Y(_11924_));
 sky130_as_sc_hs__and2_2 _42678_ (.A(net427),
    .B(net418),
    .Y(_11925_));
 sky130_as_sc_hs__and2_2 _42679_ (.A(net433),
    .B(net419),
    .Y(_11926_));
 sky130_as_sc_hs__or2_2 _42681_ (.A(_11925_),
    .B(_11926_),
    .Y(_11928_));
 sky130_as_sc_hs__and2_2 _42682_ (.A(_11927_),
    .B(_11928_),
    .Y(_11929_));
 sky130_as_sc_hs__or2_2 _42685_ (.A(_11929_),
    .B(_11930_),
    .Y(_11932_));
 sky130_as_sc_hs__and2_2 _42686_ (.A(_11931_),
    .B(_11932_),
    .Y(_11933_));
 sky130_as_sc_hs__nor2b_2 _42687_ (.A(_11639_),
    .Y(_11934_),
    .B(_11795_));
 sky130_as_sc_hs__nor2_2 _42688_ (.A(_11793_),
    .B(_11934_),
    .Y(_11935_));
 sky130_as_sc_hs__or2_2 _42690_ (.A(_11933_),
    .B(_11935_),
    .Y(_11937_));
 sky130_as_sc_hs__or2_2 _42693_ (.A(_11924_),
    .B(_11938_),
    .Y(_11940_));
 sky130_as_sc_hs__and2_2 _42694_ (.A(_11939_),
    .B(_11940_),
    .Y(_11941_));
 sky130_as_sc_hs__or2_2 _42698_ (.A(_11941_),
    .B(_11943_),
    .Y(_11945_));
 sky130_as_sc_hs__and2_2 _42699_ (.A(_11944_),
    .B(_11945_),
    .Y(_11946_));
 sky130_as_sc_hs__or2_2 _42701_ (.A(_11923_),
    .B(_11946_),
    .Y(_11948_));
 sky130_as_sc_hs__and2_2 _42702_ (.A(_11947_),
    .B(_11948_),
    .Y(_11949_));
 sky130_as_sc_hs__or2_2 _42705_ (.A(_11949_),
    .B(_11950_),
    .Y(_11952_));
 sky130_as_sc_hs__and2_2 _42706_ (.A(_11951_),
    .B(_11952_),
    .Y(_11953_));
 sky130_as_sc_hs__and2_2 _42708_ (.A(net123),
    .B(net421),
    .Y(_11955_));
 sky130_as_sc_hs__and2_2 _42709_ (.A(net120),
    .B(net128),
    .Y(_11956_));
 sky130_as_sc_hs__or2_2 _42711_ (.A(_11955_),
    .B(_11956_),
    .Y(_11958_));
 sky130_as_sc_hs__or2_2 _42713_ (.A(_11810_),
    .B(_11959_),
    .Y(_11960_));
 sky130_as_sc_hs__and2_2 _42715_ (.A(_11960_),
    .B(_11961_),
    .Y(_11962_));
 sky130_as_sc_hs__or2_2 _42717_ (.A(_11954_),
    .B(_11962_),
    .Y(_11964_));
 sky130_as_sc_hs__and2_2 _42718_ (.A(_11963_),
    .B(_11964_),
    .Y(_11965_));
 sky130_as_sc_hs__or2_2 _42720_ (.A(_11953_),
    .B(_11965_),
    .Y(_11967_));
 sky130_as_sc_hs__and2_2 _42721_ (.A(_11966_),
    .B(_11967_),
    .Y(_11968_));
 sky130_as_sc_hs__or2_2 _42724_ (.A(_11968_),
    .B(_11969_),
    .Y(_11971_));
 sky130_as_sc_hs__and2_2 _42725_ (.A(_11970_),
    .B(_11971_),
    .Y(_11972_));
 sky130_as_sc_hs__or2_2 _42728_ (.A(_11972_),
    .B(_11973_),
    .Y(_11975_));
 sky130_as_sc_hs__and2_2 _42729_ (.A(_11974_),
    .B(_11975_),
    .Y(_11976_));
 sky130_as_sc_hs__or2_2 _42732_ (.A(_11976_),
    .B(_11977_),
    .Y(_11979_));
 sky130_as_sc_hs__and2_2 _42733_ (.A(_11978_),
    .B(_11979_),
    .Y(_11980_));
 sky130_as_sc_hs__or2_2 _42734_ (.A(_11848_),
    .B(_11980_),
    .Y(_11981_));
 sky130_as_sc_hs__or2_2 _42738_ (.A(_11922_),
    .B(_11983_),
    .Y(_11985_));
 sky130_as_sc_hs__and2_2 _42739_ (.A(_11984_),
    .B(_11985_),
    .Y(_11986_));
 sky130_as_sc_hs__or2_2 _42742_ (.A(_11986_),
    .B(_11987_),
    .Y(_11989_));
 sky130_as_sc_hs__nand3_2 _42743_ (.A(net141),
    .B(_11988_),
    .C(_11989_),
    .Y(_11990_));
 sky130_as_sc_hs__or2_2 _42745_ (.A(_05474_),
    .B(_11991_),
    .Y(_11992_));
 sky130_as_sc_hs__nand3_2 _42747_ (.A(net138),
    .B(_11992_),
    .C(_11993_),
    .Y(_11994_));
 sky130_as_sc_hs__or2_2 _42750_ (.A(_05583_),
    .B(_11996_),
    .Y(_11997_));
 sky130_as_sc_hs__and2_2 _42752_ (.A(_11997_),
    .B(_11998_),
    .Y(_11999_));
 sky130_as_sc_hs__or2_2 _42754_ (.A(_05583_),
    .B(_05903_),
    .Y(_12001_));
 sky130_as_sc_hs__nand3_2 _42757_ (.A(net118),
    .B(_12000_),
    .C(_12003_),
    .Y(_12004_));
 sky130_as_sc_hs__or2_2 _42758_ (.A(\tholin_riscv.div_res[24] ),
    .B(_11875_),
    .Y(_12005_));
 sky130_as_sc_hs__and2_2 _42759_ (.A(net414),
    .B(_12005_),
    .Y(_12006_));
 sky130_as_sc_hs__or2_2 _42761_ (.A(\tholin_riscv.div_res[25] ),
    .B(_12006_),
    .Y(_12008_));
 sky130_as_sc_hs__nand3_2 _42762_ (.A(net110),
    .B(_12007_),
    .C(_12008_),
    .Y(_12009_));
 sky130_as_sc_hs__or2_2 _42763_ (.A(\tholin_riscv.div_shifter[56] ),
    .B(_11880_),
    .Y(_12010_));
 sky130_as_sc_hs__and2_2 _42764_ (.A(_21655_),
    .B(_12010_),
    .Y(_12011_));
 sky130_as_sc_hs__or2_2 _42766_ (.A(\tholin_riscv.div_shifter[57] ),
    .B(_12011_),
    .Y(_12013_));
 sky130_as_sc_hs__nand3_2 _42767_ (.A(net107),
    .B(_12012_),
    .C(_12013_),
    .Y(_12014_));
 sky130_as_sc_hs__and2_2 _42768_ (.A(_05968_),
    .B(_08110_),
    .Y(_12015_));
 sky130_as_sc_hs__nor2_2 _42773_ (.A(_05581_),
    .B(_06161_),
    .Y(_12020_));
 sky130_as_sc_hs__nand3_2 _42776_ (.A(net413),
    .B(_12021_),
    .C(_12022_),
    .Y(_12023_));
 sky130_as_sc_hs__nor2_2 _42777_ (.A(_12020_),
    .B(_12023_),
    .Y(_12024_));
 sky130_as_sc_hs__nand3_2 _42778_ (.A(_12016_),
    .B(_12019_),
    .C(_12024_),
    .Y(_12025_));
 sky130_as_sc_hs__nor2_2 _42779_ (.A(_12015_),
    .B(_12025_),
    .Y(_12026_));
 sky130_as_sc_hs__and2_2 _42780_ (.A(_12014_),
    .B(_12026_),
    .Y(_12027_));
 sky130_as_sc_hs__and2_2 _42781_ (.A(_12009_),
    .B(_12027_),
    .Y(_12028_));
 sky130_as_sc_hs__and2_2 _42782_ (.A(_12004_),
    .B(_12028_),
    .Y(_12029_));
 sky130_as_sc_hs__nand3_2 _42783_ (.A(_11990_),
    .B(_11994_),
    .C(_12029_),
    .Y(_12030_));
 sky130_as_sc_hs__or2_2 _42785_ (.A(\tholin_riscv.PC[25] ),
    .B(\tholin_riscv.Bimm[5] ),
    .Y(_12032_));
 sky130_as_sc_hs__and2_2 _42788_ (.A(_11902_),
    .B(_12034_),
    .Y(_12035_));
 sky130_as_sc_hs__or2_2 _42790_ (.A(_12033_),
    .B(_12035_),
    .Y(_12037_));
 sky130_as_sc_hs__nand3_2 _42791_ (.A(net117),
    .B(_12036_),
    .C(_12037_),
    .Y(_12038_));
 sky130_as_sc_hs__and2_2 _42792_ (.A(\tholin_riscv.PC[25] ),
    .B(_11909_),
    .Y(_12039_));
 sky130_as_sc_hs__nor2_2 _42793_ (.A(\tholin_riscv.PC[25] ),
    .B(_11909_),
    .Y(_12040_));
 sky130_as_sc_hs__nor2_2 _42794_ (.A(_12039_),
    .B(_12040_),
    .Y(_12041_));
 sky130_as_sc_hs__inv_2 _42795_ (.Y(_12042_),
    .A(_12041_));
 sky130_as_sc_hs__and2_2 _42798_ (.A(_21569_),
    .B(_12044_),
    .Y(_12045_));
 sky130_as_sc_hs__nand3_2 _42799_ (.A(_12038_),
    .B(_12043_),
    .C(_12045_),
    .Y(_12046_));
 sky130_as_sc_hs__nand3_2 _42800_ (.A(_21546_),
    .B(_12030_),
    .C(_12046_),
    .Y(_12047_));
 sky130_as_sc_hs__and2_2 _42805_ (.A(\tholin_riscv.Bimm[6] ),
    .B(net371),
    .Y(_12051_));
 sky130_as_sc_hs__or2_2 _42806_ (.A(_10352_),
    .B(_12051_),
    .Y(_12052_));
 sky130_as_sc_hs__and2_2 _42808_ (.A(net425),
    .B(net419),
    .Y(_12054_));
 sky130_as_sc_hs__and2_2 _42809_ (.A(_11793_),
    .B(_11933_),
    .Y(_12055_));
 sky130_as_sc_hs__and2_2 _42810_ (.A(net120),
    .B(net418),
    .Y(_12056_));
 sky130_as_sc_hs__and2_2 _42811_ (.A(net433),
    .B(net74),
    .Y(_12057_));
 sky130_as_sc_hs__or2_2 _42812_ (.A(_12056_),
    .B(_12057_),
    .Y(_12058_));
 sky130_as_sc_hs__and2_2 _42814_ (.A(_12058_),
    .B(_12059_),
    .Y(_12060_));
 sky130_as_sc_hs__or2_2 _42816_ (.A(_12060_),
    .B(_12061_),
    .Y(_12062_));
 sky130_as_sc_hs__and2_2 _42818_ (.A(_12062_),
    .B(_12063_),
    .Y(_12064_));
 sky130_as_sc_hs__or2_2 _42820_ (.A(_12055_),
    .B(_12064_),
    .Y(_12066_));
 sky130_as_sc_hs__and2_2 _42821_ (.A(_12065_),
    .B(_12066_),
    .Y(_12067_));
 sky130_as_sc_hs__or2_2 _42823_ (.A(_12054_),
    .B(_12067_),
    .Y(_12069_));
 sky130_as_sc_hs__and2_2 _42824_ (.A(_12068_),
    .B(_12069_),
    .Y(_12070_));
 sky130_as_sc_hs__or2_2 _42828_ (.A(_12070_),
    .B(_12072_),
    .Y(_12074_));
 sky130_as_sc_hs__and2_2 _42829_ (.A(_12073_),
    .B(_12074_),
    .Y(_12075_));
 sky130_as_sc_hs__or2_2 _42832_ (.A(_12075_),
    .B(_12076_),
    .Y(_12078_));
 sky130_as_sc_hs__and2_2 _42834_ (.A(net123),
    .B(net128),
    .Y(_12080_));
 sky130_as_sc_hs__and2_2 _42835_ (.A(net423),
    .B(net421),
    .Y(_12081_));
 sky130_as_sc_hs__and2_2 _42836_ (.A(_12080_),
    .B(_12081_),
    .Y(_12082_));
 sky130_as_sc_hs__or2_2 _42839_ (.A(_11957_),
    .B(_12082_),
    .Y(_12085_));
 sky130_as_sc_hs__or2_2 _42840_ (.A(_12080_),
    .B(_12081_),
    .Y(_12086_));
 sky130_as_sc_hs__nand3_2 _42841_ (.A(_12084_),
    .B(_12085_),
    .C(_12086_),
    .Y(_12087_));
 sky130_as_sc_hs__or2_2 _42842_ (.A(_12079_),
    .B(_12087_),
    .Y(_12088_));
 sky130_as_sc_hs__and2_2 _42844_ (.A(_12088_),
    .B(_12089_),
    .Y(_12090_));
 sky130_as_sc_hs__or2_2 _42847_ (.A(_12090_),
    .B(_12091_),
    .Y(_12093_));
 sky130_as_sc_hs__and2_2 _42848_ (.A(_12092_),
    .B(_12093_),
    .Y(_12094_));
 sky130_as_sc_hs__or2_2 _42851_ (.A(_12094_),
    .B(_12095_),
    .Y(_12097_));
 sky130_as_sc_hs__and2_2 _42852_ (.A(_12096_),
    .B(_12097_),
    .Y(_12098_));
 sky130_as_sc_hs__or2_2 _42855_ (.A(_12098_),
    .B(_12099_),
    .Y(_12101_));
 sky130_as_sc_hs__or2_2 _42857_ (.A(_11978_),
    .B(_12102_),
    .Y(_12103_));
 sky130_as_sc_hs__and2_2 _42859_ (.A(_12103_),
    .B(_12104_),
    .Y(_12105_));
 sky130_as_sc_hs__nand3_2 _42860_ (.A(_11781_),
    .B(_11853_),
    .C(_11983_),
    .Y(_12106_));
 sky130_as_sc_hs__or2_2 _42865_ (.A(_12105_),
    .B(_12109_),
    .Y(_12111_));
 sky130_as_sc_hs__and2_2 _42867_ (.A(_11856_),
    .B(_11986_),
    .Y(_12113_));
 sky130_as_sc_hs__or2_2 _42868_ (.A(_05505_),
    .B(_12113_),
    .Y(_12114_));
 sky130_as_sc_hs__and2_2 _42869_ (.A(_11858_),
    .B(_12114_),
    .Y(_12115_));
 sky130_as_sc_hs__or2_2 _42870_ (.A(_12112_),
    .B(_12115_),
    .Y(_12116_));
 sky130_as_sc_hs__nand3_2 _42872_ (.A(net141),
    .B(_12116_),
    .C(_12117_),
    .Y(_12118_));
 sky130_as_sc_hs__or2_2 _42873_ (.A(_05475_),
    .B(_05505_),
    .Y(_12119_));
 sky130_as_sc_hs__and2_2 _42874_ (.A(_11862_),
    .B(_12119_),
    .Y(_12120_));
 sky130_as_sc_hs__or2_2 _42875_ (.A(_05467_),
    .B(_12120_),
    .Y(_12121_));
 sky130_as_sc_hs__nand3_2 _42877_ (.A(net138),
    .B(_12121_),
    .C(_12122_),
    .Y(_12123_));
 sky130_as_sc_hs__or2_2 _42880_ (.A(_05574_),
    .B(_12125_),
    .Y(_12126_));
 sky130_as_sc_hs__and2_2 _42882_ (.A(_12126_),
    .B(_12127_),
    .Y(_12128_));
 sky130_as_sc_hs__or2_2 _42884_ (.A(_05574_),
    .B(_05905_),
    .Y(_12130_));
 sky130_as_sc_hs__nand3_2 _42887_ (.A(net118),
    .B(_12129_),
    .C(_12132_),
    .Y(_12133_));
 sky130_as_sc_hs__or2_2 _42888_ (.A(\tholin_riscv.div_res[25] ),
    .B(_12005_),
    .Y(_12134_));
 sky130_as_sc_hs__and2_2 _42889_ (.A(net414),
    .B(_12134_),
    .Y(_12135_));
 sky130_as_sc_hs__or2_2 _42891_ (.A(\tholin_riscv.div_res[26] ),
    .B(_12135_),
    .Y(_12137_));
 sky130_as_sc_hs__nand3_2 _42892_ (.A(net110),
    .B(_12136_),
    .C(_12137_),
    .Y(_12138_));
 sky130_as_sc_hs__or2_2 _42893_ (.A(\tholin_riscv.div_shifter[57] ),
    .B(_12010_),
    .Y(_12139_));
 sky130_as_sc_hs__and2_2 _42894_ (.A(_21655_),
    .B(_12139_),
    .Y(_12140_));
 sky130_as_sc_hs__or2_2 _42896_ (.A(\tholin_riscv.div_shifter[58] ),
    .B(_12140_),
    .Y(_12142_));
 sky130_as_sc_hs__nand3_2 _42897_ (.A(net107),
    .B(_12141_),
    .C(_12142_),
    .Y(_12143_));
 sky130_as_sc_hs__and2_2 _42898_ (.A(net140),
    .B(_07815_),
    .Y(_12144_));
 sky130_as_sc_hs__nor2_2 _42903_ (.A(_05572_),
    .B(_06161_),
    .Y(_12149_));
 sky130_as_sc_hs__nand3_2 _42906_ (.A(net412),
    .B(_12150_),
    .C(_12151_),
    .Y(_12152_));
 sky130_as_sc_hs__nor2_2 _42907_ (.A(_12149_),
    .B(_12152_),
    .Y(_12153_));
 sky130_as_sc_hs__nand3_2 _42908_ (.A(_12145_),
    .B(_12148_),
    .C(_12153_),
    .Y(_12154_));
 sky130_as_sc_hs__nor2_2 _42909_ (.A(_12144_),
    .B(_12154_),
    .Y(_12155_));
 sky130_as_sc_hs__and2_2 _42910_ (.A(_12143_),
    .B(_12155_),
    .Y(_12156_));
 sky130_as_sc_hs__and2_2 _42911_ (.A(_12138_),
    .B(_12156_),
    .Y(_12157_));
 sky130_as_sc_hs__and2_2 _42912_ (.A(_12133_),
    .B(_12157_),
    .Y(_12158_));
 sky130_as_sc_hs__nand3_2 _42913_ (.A(_12118_),
    .B(_12123_),
    .C(_12158_),
    .Y(_12159_));
 sky130_as_sc_hs__or2_2 _42916_ (.A(\tholin_riscv.PC[26] ),
    .B(\tholin_riscv.Bimm[6] ),
    .Y(_12162_));
 sky130_as_sc_hs__or2_2 _42918_ (.A(_12160_),
    .B(_12163_),
    .Y(_12164_));
 sky130_as_sc_hs__nand3_2 _42920_ (.A(net117),
    .B(_12164_),
    .C(_12165_),
    .Y(_12166_));
 sky130_as_sc_hs__or2_2 _42921_ (.A(\tholin_riscv.Bimm[6] ),
    .B(_21590_),
    .Y(_12167_));
 sky130_as_sc_hs__and2_2 _42922_ (.A(\tholin_riscv.PC[26] ),
    .B(_12039_),
    .Y(_12168_));
 sky130_as_sc_hs__nor2_2 _42923_ (.A(\tholin_riscv.PC[26] ),
    .B(_12039_),
    .Y(_12169_));
 sky130_as_sc_hs__or2_2 _42924_ (.A(_12168_),
    .B(_12169_),
    .Y(_12170_));
 sky130_as_sc_hs__nand3_2 _42926_ (.A(_12166_),
    .B(_12167_),
    .C(_12171_),
    .Y(_12172_));
 sky130_as_sc_hs__nand3_2 _42928_ (.A(_21546_),
    .B(_12159_),
    .C(_12173_),
    .Y(_12174_));
 sky130_as_sc_hs__and2_2 _42933_ (.A(\tholin_riscv.Bimm[7] ),
    .B(\tholin_riscv.io_size[1] ),
    .Y(_12178_));
 sky130_as_sc_hs__or2_2 _42934_ (.A(_10352_),
    .B(_12178_),
    .Y(_12179_));
 sky130_as_sc_hs__and2_2 _42936_ (.A(_12103_),
    .B(_12110_),
    .Y(_12181_));
 sky130_as_sc_hs__and2_2 _42937_ (.A(net425),
    .B(net74),
    .Y(_12182_));
 sky130_as_sc_hs__nor2b_2 _42938_ (.A(_11927_),
    .Y(_12183_),
    .B(_12060_));
 sky130_as_sc_hs__nand3_2 _42941_ (.A(net122),
    .B(_12056_),
    .C(_12057_),
    .Y(_12186_));
 sky130_as_sc_hs__inv_2 _42942_ (.Y(_12187_),
    .A(_12186_));
 sky130_as_sc_hs__and2_2 _42943_ (.A(_12185_),
    .B(_12186_),
    .Y(_12188_));
 sky130_as_sc_hs__or2_2 _42945_ (.A(_12183_),
    .B(_12188_),
    .Y(_12190_));
 sky130_as_sc_hs__and2_2 _42946_ (.A(_12189_),
    .B(_12190_),
    .Y(_12191_));
 sky130_as_sc_hs__nor2b_2 _42947_ (.A(_11931_),
    .Y(_12192_),
    .B(_12060_));
 sky130_as_sc_hs__or2_2 _42949_ (.A(_12191_),
    .B(_12192_),
    .Y(_12194_));
 sky130_as_sc_hs__and2_2 _42950_ (.A(_12193_),
    .B(_12194_),
    .Y(_12195_));
 sky130_as_sc_hs__or2_2 _42952_ (.A(_12182_),
    .B(_12195_),
    .Y(_12197_));
 sky130_as_sc_hs__and2_2 _42953_ (.A(_12196_),
    .B(_12197_),
    .Y(_12198_));
 sky130_as_sc_hs__or2_2 _42956_ (.A(_12198_),
    .B(_12199_),
    .Y(_12201_));
 sky130_as_sc_hs__or2_2 _42958_ (.A(_12073_),
    .B(_12202_),
    .Y(_12203_));
 sky130_as_sc_hs__and2_2 _42961_ (.A(net423),
    .B(net128),
    .Y(_12206_));
 sky130_as_sc_hs__and2_2 _42962_ (.A(net421),
    .B(net420),
    .Y(_12207_));
 sky130_as_sc_hs__and2_2 _42963_ (.A(_12206_),
    .B(_12207_),
    .Y(_12208_));
 sky130_as_sc_hs__or2_2 _42965_ (.A(_12083_),
    .B(_12208_),
    .Y(_12210_));
 sky130_as_sc_hs__or2_2 _42966_ (.A(_12206_),
    .B(_12207_),
    .Y(_12211_));
 sky130_as_sc_hs__nand3_2 _42967_ (.A(_12209_),
    .B(_12210_),
    .C(_12211_),
    .Y(_12212_));
 sky130_as_sc_hs__or2_2 _42968_ (.A(_12205_),
    .B(_12212_),
    .Y(_12213_));
 sky130_as_sc_hs__and2_2 _42970_ (.A(_12213_),
    .B(_12214_),
    .Y(_12215_));
 sky130_as_sc_hs__or2_2 _42973_ (.A(_12215_),
    .B(_12216_),
    .Y(_12218_));
 sky130_as_sc_hs__or2_2 _42975_ (.A(_12085_),
    .B(_12219_),
    .Y(_12220_));
 sky130_as_sc_hs__and2_2 _42977_ (.A(_12220_),
    .B(_12221_),
    .Y(_12222_));
 sky130_as_sc_hs__or2_2 _42980_ (.A(_12222_),
    .B(_12223_),
    .Y(_12225_));
 sky130_as_sc_hs__and2_2 _42981_ (.A(_12224_),
    .B(_12225_),
    .Y(_12226_));
 sky130_as_sc_hs__or2_2 _42982_ (.A(_12100_),
    .B(_12226_),
    .Y(_12227_));
 sky130_as_sc_hs__or2_2 _42986_ (.A(_12181_),
    .B(_12229_),
    .Y(_12231_));
 sky130_as_sc_hs__and2_2 _42987_ (.A(_12230_),
    .B(_12231_),
    .Y(_12232_));
 sky130_as_sc_hs__and2_2 _42988_ (.A(_12112_),
    .B(_12113_),
    .Y(_12233_));
 sky130_as_sc_hs__or2_2 _42989_ (.A(_05505_),
    .B(_12233_),
    .Y(_12234_));
 sky130_as_sc_hs__and2_2 _42990_ (.A(_11858_),
    .B(_12234_),
    .Y(_12235_));
 sky130_as_sc_hs__or2_2 _42992_ (.A(_12232_),
    .B(_12235_),
    .Y(_12237_));
 sky130_as_sc_hs__nand3_2 _42993_ (.A(net141),
    .B(_12236_),
    .C(_12237_),
    .Y(_12238_));
 sky130_as_sc_hs__or2_2 _42994_ (.A(_05476_),
    .B(_05505_),
    .Y(_12239_));
 sky130_as_sc_hs__and2_2 _42995_ (.A(_11862_),
    .B(_12239_),
    .Y(_12240_));
 sky130_as_sc_hs__or2_2 _42996_ (.A(_05465_),
    .B(_12240_),
    .Y(_12241_));
 sky130_as_sc_hs__nand3_2 _42998_ (.A(net138),
    .B(_12241_),
    .C(_12242_),
    .Y(_12243_));
 sky130_as_sc_hs__or2_2 _43001_ (.A(_05565_),
    .B(_12245_),
    .Y(_12246_));
 sky130_as_sc_hs__and2_2 _43003_ (.A(_12246_),
    .B(_12247_),
    .Y(_12248_));
 sky130_as_sc_hs__or2_2 _43005_ (.A(_05565_),
    .B(_05907_),
    .Y(_12250_));
 sky130_as_sc_hs__nand3_2 _43008_ (.A(net118),
    .B(_12249_),
    .C(_12252_),
    .Y(_12253_));
 sky130_as_sc_hs__or2_2 _43009_ (.A(\tholin_riscv.div_res[26] ),
    .B(_12134_),
    .Y(_12254_));
 sky130_as_sc_hs__and2_2 _43010_ (.A(net414),
    .B(_12254_),
    .Y(_12255_));
 sky130_as_sc_hs__or2_2 _43012_ (.A(\tholin_riscv.div_res[27] ),
    .B(_12255_),
    .Y(_12257_));
 sky130_as_sc_hs__nand3_2 _43013_ (.A(net110),
    .B(_12256_),
    .C(_12257_),
    .Y(_12258_));
 sky130_as_sc_hs__or2_2 _43014_ (.A(\tholin_riscv.div_shifter[58] ),
    .B(_12139_),
    .Y(_12259_));
 sky130_as_sc_hs__and2_2 _43015_ (.A(_21655_),
    .B(_12259_),
    .Y(_12260_));
 sky130_as_sc_hs__or2_2 _43017_ (.A(\tholin_riscv.div_shifter[59] ),
    .B(_12260_),
    .Y(_12262_));
 sky130_as_sc_hs__nand3_2 _43018_ (.A(net107),
    .B(_12261_),
    .C(_12262_),
    .Y(_12263_));
 sky130_as_sc_hs__and2_2 _43019_ (.A(_05968_),
    .B(_07528_),
    .Y(_12264_));
 sky130_as_sc_hs__nor2_2 _43024_ (.A(_05563_),
    .B(_06161_),
    .Y(_12269_));
 sky130_as_sc_hs__nand3_2 _43027_ (.A(net412),
    .B(_12270_),
    .C(_12271_),
    .Y(_12272_));
 sky130_as_sc_hs__nor2_2 _43028_ (.A(_12269_),
    .B(_12272_),
    .Y(_12273_));
 sky130_as_sc_hs__nand3_2 _43029_ (.A(_12265_),
    .B(_12268_),
    .C(_12273_),
    .Y(_12274_));
 sky130_as_sc_hs__nor2_2 _43030_ (.A(_12264_),
    .B(_12274_),
    .Y(_12275_));
 sky130_as_sc_hs__and2_2 _43031_ (.A(_12263_),
    .B(_12275_),
    .Y(_12276_));
 sky130_as_sc_hs__and2_2 _43032_ (.A(_12258_),
    .B(_12276_),
    .Y(_12277_));
 sky130_as_sc_hs__and2_2 _43033_ (.A(_12253_),
    .B(_12277_),
    .Y(_12278_));
 sky130_as_sc_hs__nand3_2 _43034_ (.A(_12238_),
    .B(_12243_),
    .C(_12278_),
    .Y(_12279_));
 sky130_as_sc_hs__or2_2 _43036_ (.A(\tholin_riscv.PC[27] ),
    .B(\tholin_riscv.Bimm[7] ),
    .Y(_12281_));
 sky130_as_sc_hs__and2_2 _43037_ (.A(_12280_),
    .B(_12281_),
    .Y(_12282_));
 sky130_as_sc_hs__or2_2 _43041_ (.A(_12282_),
    .B(_12284_),
    .Y(_12286_));
 sky130_as_sc_hs__and2_2 _43044_ (.A(\tholin_riscv.PC[27] ),
    .B(_12168_),
    .Y(_12289_));
 sky130_as_sc_hs__nor2_2 _43045_ (.A(\tholin_riscv.PC[27] ),
    .B(_12168_),
    .Y(_12290_));
 sky130_as_sc_hs__or2_2 _43046_ (.A(_12289_),
    .B(_12290_),
    .Y(_12291_));
 sky130_as_sc_hs__nand3_2 _43049_ (.A(_12288_),
    .B(_12292_),
    .C(_12293_),
    .Y(_12294_));
 sky130_as_sc_hs__nand3_2 _43051_ (.A(_21546_),
    .B(_12279_),
    .C(_12295_),
    .Y(_12296_));
 sky130_as_sc_hs__and2_2 _43056_ (.A(\tholin_riscv.Bimm[8] ),
    .B(net371),
    .Y(_12300_));
 sky130_as_sc_hs__or2_2 _43057_ (.A(_10352_),
    .B(_12300_),
    .Y(_12301_));
 sky130_as_sc_hs__and2_2 _43060_ (.A(net423),
    .B(net418),
    .Y(_12304_));
 sky130_as_sc_hs__inv_2 _43063_ (.Y(_12307_),
    .A(_12306_));
 sky130_as_sc_hs__or2_2 _43064_ (.A(_12304_),
    .B(_12305_),
    .Y(_12308_));
 sky130_as_sc_hs__and2_2 _43065_ (.A(_12306_),
    .B(_12308_),
    .Y(_12309_));
 sky130_as_sc_hs__or2_2 _43067_ (.A(_12303_),
    .B(_12309_),
    .Y(_12311_));
 sky130_as_sc_hs__or2_2 _43069_ (.A(_12200_),
    .B(_12312_),
    .Y(_12313_));
 sky130_as_sc_hs__and2_2 _43072_ (.A(net128),
    .B(net420),
    .Y(_12316_));
 sky130_as_sc_hs__and2_2 _43073_ (.A(net421),
    .B(net75),
    .Y(_12317_));
 sky130_as_sc_hs__or2_2 _43075_ (.A(_12208_),
    .B(_12318_),
    .Y(_12319_));
 sky130_as_sc_hs__or2_2 _43077_ (.A(_12316_),
    .B(_12317_),
    .Y(_12321_));
 sky130_as_sc_hs__nand3_2 _43078_ (.A(_12319_),
    .B(_12320_),
    .C(_12321_),
    .Y(_12322_));
 sky130_as_sc_hs__or2_2 _43079_ (.A(_12315_),
    .B(_12322_),
    .Y(_12323_));
 sky130_as_sc_hs__and2_2 _43081_ (.A(_12323_),
    .B(_12324_),
    .Y(_12325_));
 sky130_as_sc_hs__or2_2 _43084_ (.A(_12325_),
    .B(_12326_),
    .Y(_12328_));
 sky130_as_sc_hs__or2_2 _43086_ (.A(_12210_),
    .B(_12329_),
    .Y(_12330_));
 sky130_as_sc_hs__and2_2 _43088_ (.A(_12330_),
    .B(_12331_),
    .Y(_12332_));
 sky130_as_sc_hs__or2_2 _43091_ (.A(_12332_),
    .B(_12333_),
    .Y(_12335_));
 sky130_as_sc_hs__or2_2 _43093_ (.A(_12224_),
    .B(_12336_),
    .Y(_12337_));
 sky130_as_sc_hs__and2_2 _43095_ (.A(_12337_),
    .B(_12338_),
    .Y(_12339_));
 sky130_as_sc_hs__and2_2 _43096_ (.A(_12105_),
    .B(_12229_),
    .Y(_12340_));
 sky130_as_sc_hs__nand2b_2 _43097_ (.B(_12340_),
    .Y(_12341_),
    .A(_12106_));
 sky130_as_sc_hs__nand2b_2 _43098_ (.B(_12340_),
    .Y(_12342_),
    .A(_12108_));
 sky130_as_sc_hs__nand3_2 _43101_ (.A(_12341_),
    .B(_12342_),
    .C(_12344_),
    .Y(_12345_));
 sky130_as_sc_hs__or2_2 _43103_ (.A(_12339_),
    .B(_12345_),
    .Y(_12347_));
 sky130_as_sc_hs__nand3_2 _43105_ (.A(_11857_),
    .B(_12232_),
    .C(_12233_),
    .Y(_12349_));
 sky130_as_sc_hs__or2_2 _43108_ (.A(_12348_),
    .B(_12350_),
    .Y(_12352_));
 sky130_as_sc_hs__nand3_2 _43109_ (.A(net142),
    .B(_12351_),
    .C(_12352_),
    .Y(_12353_));
 sky130_as_sc_hs__or2_2 _43112_ (.A(_05483_),
    .B(_12354_),
    .Y(_12356_));
 sky130_as_sc_hs__nand3_2 _43113_ (.A(net139),
    .B(_12355_),
    .C(_12356_),
    .Y(_12357_));
 sky130_as_sc_hs__or2_2 _43115_ (.A(_05909_),
    .B(_05912_),
    .Y(_12359_));
 sky130_as_sc_hs__nand3_2 _43116_ (.A(_06527_),
    .B(_12358_),
    .C(_12359_),
    .Y(_12360_));
 sky130_as_sc_hs__or2_2 _43119_ (.A(_05912_),
    .B(_12362_),
    .Y(_12363_));
 sky130_as_sc_hs__and2_2 _43121_ (.A(_12363_),
    .B(_12364_),
    .Y(_12365_));
 sky130_as_sc_hs__or2_2 _43122_ (.A(_06527_),
    .B(_12365_),
    .Y(_12366_));
 sky130_as_sc_hs__and2_2 _43124_ (.A(net118),
    .B(_12367_),
    .Y(_12368_));
 sky130_as_sc_hs__or2_2 _43125_ (.A(\tholin_riscv.div_shifter[59] ),
    .B(_12259_),
    .Y(_12369_));
 sky130_as_sc_hs__and2_2 _43126_ (.A(_21655_),
    .B(_12369_),
    .Y(_12370_));
 sky130_as_sc_hs__or2_2 _43128_ (.A(\tholin_riscv.div_shifter[60] ),
    .B(_12370_),
    .Y(_12372_));
 sky130_as_sc_hs__nand3_2 _43129_ (.A(net107),
    .B(_12371_),
    .C(_12372_),
    .Y(_12373_));
 sky130_as_sc_hs__or2_2 _43130_ (.A(\tholin_riscv.div_res[27] ),
    .B(_12254_),
    .Y(_12374_));
 sky130_as_sc_hs__and2_2 _43131_ (.A(net414),
    .B(_12374_),
    .Y(_12375_));
 sky130_as_sc_hs__or2_2 _43133_ (.A(\tholin_riscv.div_res[28] ),
    .B(_12375_),
    .Y(_12377_));
 sky130_as_sc_hs__nand3_2 _43134_ (.A(net110),
    .B(_12376_),
    .C(_12377_),
    .Y(_12378_));
 sky130_as_sc_hs__and2_2 _43135_ (.A(net140),
    .B(_07232_),
    .Y(_12379_));
 sky130_as_sc_hs__nor2_2 _43140_ (.A(_05910_),
    .B(_06161_),
    .Y(_12384_));
 sky130_as_sc_hs__nand3_2 _43143_ (.A(net412),
    .B(_12385_),
    .C(_12386_),
    .Y(_12387_));
 sky130_as_sc_hs__nor2_2 _43144_ (.A(_12384_),
    .B(_12387_),
    .Y(_12388_));
 sky130_as_sc_hs__nand3_2 _43145_ (.A(_12380_),
    .B(_12383_),
    .C(_12388_),
    .Y(_12389_));
 sky130_as_sc_hs__nor2_2 _43146_ (.A(_12379_),
    .B(_12389_),
    .Y(_12390_));
 sky130_as_sc_hs__nand3_2 _43147_ (.A(_12373_),
    .B(_12378_),
    .C(_12390_),
    .Y(_12391_));
 sky130_as_sc_hs__nor2_2 _43148_ (.A(_12368_),
    .B(_12391_),
    .Y(_12392_));
 sky130_as_sc_hs__nand3_2 _43149_ (.A(_12353_),
    .B(_12357_),
    .C(_12392_),
    .Y(_12393_));
 sky130_as_sc_hs__or2_2 _43152_ (.A(\tholin_riscv.PC[28] ),
    .B(\tholin_riscv.Bimm[8] ),
    .Y(_12396_));
 sky130_as_sc_hs__or2_2 _43154_ (.A(_12394_),
    .B(_12397_),
    .Y(_12398_));
 sky130_as_sc_hs__nand3_2 _43156_ (.A(net117),
    .B(_12398_),
    .C(_12399_),
    .Y(_12400_));
 sky130_as_sc_hs__and2_2 _43157_ (.A(\tholin_riscv.PC[28] ),
    .B(_12289_),
    .Y(_12401_));
 sky130_as_sc_hs__nor2_2 _43158_ (.A(\tholin_riscv.PC[28] ),
    .B(_12289_),
    .Y(_12402_));
 sky130_as_sc_hs__or2_2 _43159_ (.A(_12401_),
    .B(_12402_),
    .Y(_12403_));
 sky130_as_sc_hs__nand3_2 _43162_ (.A(_12400_),
    .B(_12404_),
    .C(_12405_),
    .Y(_12406_));
 sky130_as_sc_hs__nand3_2 _43164_ (.A(_21546_),
    .B(_12393_),
    .C(_12407_),
    .Y(_12408_));
 sky130_as_sc_hs__and2_2 _43169_ (.A(net419),
    .B(_12307_),
    .Y(_12412_));
 sky130_as_sc_hs__and2_2 _43170_ (.A(net423),
    .B(_12187_),
    .Y(_12413_));
 sky130_as_sc_hs__or2_2 _43171_ (.A(net419),
    .B(_12413_),
    .Y(_12414_));
 sky130_as_sc_hs__or2_2 _43173_ (.A(_12412_),
    .B(_12415_),
    .Y(_12416_));
 sky130_as_sc_hs__or2_2 _43174_ (.A(_12310_),
    .B(_12416_),
    .Y(_12417_));
 sky130_as_sc_hs__and2_2 _43176_ (.A(_12417_),
    .B(_12418_),
    .Y(_12419_));
 sky130_as_sc_hs__nor2_2 _43178_ (.A(_12207_),
    .B(_12420_),
    .Y(_12421_));
 sky130_as_sc_hs__or2_2 _43180_ (.A(_12419_),
    .B(_12421_),
    .Y(_12423_));
 sky130_as_sc_hs__and2_2 _43181_ (.A(_12422_),
    .B(_12423_),
    .Y(_12424_));
 sky130_as_sc_hs__or2_2 _43184_ (.A(_12424_),
    .B(_12425_),
    .Y(_12427_));
 sky130_as_sc_hs__or2_2 _43186_ (.A(_12320_),
    .B(_12428_),
    .Y(_12429_));
 sky130_as_sc_hs__and2_2 _43188_ (.A(_12429_),
    .B(_12430_),
    .Y(_12431_));
 sky130_as_sc_hs__or2_2 _43191_ (.A(_12431_),
    .B(_12432_),
    .Y(_12434_));
 sky130_as_sc_hs__nor2_2 _43193_ (.A(_12334_),
    .B(_12435_),
    .Y(_12436_));
 sky130_as_sc_hs__and2_2 _43194_ (.A(_12334_),
    .B(_12435_),
    .Y(_12437_));
 sky130_as_sc_hs__nor2_2 _43195_ (.A(_12436_),
    .B(_12437_),
    .Y(_12438_));
 sky130_as_sc_hs__or2_2 _43198_ (.A(_12438_),
    .B(_12439_),
    .Y(_12441_));
 sky130_as_sc_hs__or2_2 _43202_ (.A(_12442_),
    .B(_12443_),
    .Y(_12445_));
 sky130_as_sc_hs__nand3_2 _43203_ (.A(net141),
    .B(_12444_),
    .C(_12445_),
    .Y(_12446_));
 sky130_as_sc_hs__or2_2 _43205_ (.A(_05487_),
    .B(_12447_),
    .Y(_12448_));
 sky130_as_sc_hs__nand3_2 _43207_ (.A(net138),
    .B(_12448_),
    .C(_12449_),
    .Y(_12450_));
 sky130_as_sc_hs__or2_2 _43210_ (.A(_05545_),
    .B(_12452_),
    .Y(_12453_));
 sky130_as_sc_hs__and2_2 _43212_ (.A(_12453_),
    .B(_12454_),
    .Y(_12455_));
 sky130_as_sc_hs__or2_2 _43216_ (.A(_05545_),
    .B(_12457_),
    .Y(_12459_));
 sky130_as_sc_hs__nand3_2 _43219_ (.A(net118),
    .B(_12456_),
    .C(_12461_),
    .Y(_12462_));
 sky130_as_sc_hs__or2_2 _43220_ (.A(\tholin_riscv.div_res[28] ),
    .B(_12374_),
    .Y(_12463_));
 sky130_as_sc_hs__and2_2 _43221_ (.A(net414),
    .B(_12463_),
    .Y(_12464_));
 sky130_as_sc_hs__or2_2 _43223_ (.A(\tholin_riscv.div_res[29] ),
    .B(_12464_),
    .Y(_12466_));
 sky130_as_sc_hs__nand3_2 _43224_ (.A(net110),
    .B(_12465_),
    .C(_12466_),
    .Y(_12467_));
 sky130_as_sc_hs__or2_2 _43225_ (.A(\tholin_riscv.div_shifter[60] ),
    .B(_12369_),
    .Y(_12468_));
 sky130_as_sc_hs__and2_2 _43226_ (.A(_21655_),
    .B(_12468_),
    .Y(_12469_));
 sky130_as_sc_hs__or2_2 _43228_ (.A(\tholin_riscv.div_shifter[61] ),
    .B(_12469_),
    .Y(_12471_));
 sky130_as_sc_hs__nand3_2 _43229_ (.A(net107),
    .B(_12470_),
    .C(_12471_),
    .Y(_12472_));
 sky130_as_sc_hs__and2_2 _43230_ (.A(_05968_),
    .B(_06910_),
    .Y(_12473_));
 sky130_as_sc_hs__nor2_2 _43235_ (.A(_05543_),
    .B(_06161_),
    .Y(_12478_));
 sky130_as_sc_hs__nand3_2 _43238_ (.A(net412),
    .B(_12479_),
    .C(_12480_),
    .Y(_12481_));
 sky130_as_sc_hs__nor2_2 _43239_ (.A(_12478_),
    .B(_12481_),
    .Y(_12482_));
 sky130_as_sc_hs__nand3_2 _43240_ (.A(_12474_),
    .B(_12477_),
    .C(_12482_),
    .Y(_12483_));
 sky130_as_sc_hs__nor2_2 _43241_ (.A(_12473_),
    .B(_12483_),
    .Y(_12484_));
 sky130_as_sc_hs__and2_2 _43242_ (.A(_12472_),
    .B(_12484_),
    .Y(_12485_));
 sky130_as_sc_hs__and2_2 _43243_ (.A(_12467_),
    .B(_12485_),
    .Y(_12486_));
 sky130_as_sc_hs__and2_2 _43244_ (.A(_12462_),
    .B(_12486_),
    .Y(_12487_));
 sky130_as_sc_hs__nand3_2 _43245_ (.A(_12446_),
    .B(_12450_),
    .C(_12487_),
    .Y(_12488_));
 sky130_as_sc_hs__or2_2 _43249_ (.A(\tholin_riscv.PC[29] ),
    .B(\tholin_riscv.Bimm[9] ),
    .Y(_12492_));
 sky130_as_sc_hs__or2_2 _43251_ (.A(_12490_),
    .B(_12493_),
    .Y(_12494_));
 sky130_as_sc_hs__nand3_2 _43253_ (.A(net117),
    .B(_12494_),
    .C(_12495_),
    .Y(_12496_));
 sky130_as_sc_hs__and2_2 _43254_ (.A(\tholin_riscv.PC[29] ),
    .B(_12401_),
    .Y(_12497_));
 sky130_as_sc_hs__nor2_2 _43255_ (.A(\tholin_riscv.PC[29] ),
    .B(_12401_),
    .Y(_12498_));
 sky130_as_sc_hs__or2_2 _43256_ (.A(_12497_),
    .B(_12498_),
    .Y(_12499_));
 sky130_as_sc_hs__or2_2 _43258_ (.A(\tholin_riscv.Bimm[9] ),
    .B(_21590_),
    .Y(_12501_));
 sky130_as_sc_hs__nand3_2 _43259_ (.A(_12496_),
    .B(_12500_),
    .C(_12501_),
    .Y(_12502_));
 sky130_as_sc_hs__nand3_2 _43261_ (.A(_21546_),
    .B(_12488_),
    .C(_12503_),
    .Y(_12504_));
 sky130_as_sc_hs__and2_2 _43262_ (.A(\tholin_riscv.Bimm[9] ),
    .B(net371),
    .Y(_12505_));
 sky130_as_sc_hs__or2_2 _43263_ (.A(_10352_),
    .B(_12505_),
    .Y(_12506_));
 sky130_as_sc_hs__and2_2 _43271_ (.A(net418),
    .B(net74),
    .Y(_12513_));
 sky130_as_sc_hs__or2_2 _43272_ (.A(_12412_),
    .B(_12513_),
    .Y(_12514_));
 sky130_as_sc_hs__and2_2 _43273_ (.A(_12512_),
    .B(_12514_),
    .Y(_12515_));
 sky130_as_sc_hs__or2_2 _43275_ (.A(_12511_),
    .B(_12515_),
    .Y(_12517_));
 sky130_as_sc_hs__or2_2 _43277_ (.A(_12318_),
    .B(_12518_),
    .Y(_12519_));
 sky130_as_sc_hs__and2_2 _43279_ (.A(_12519_),
    .B(_12520_),
    .Y(_12521_));
 sky130_as_sc_hs__or2_2 _43282_ (.A(_12521_),
    .B(_12522_),
    .Y(_12524_));
 sky130_as_sc_hs__or2_2 _43284_ (.A(_12433_),
    .B(_12525_),
    .Y(_12526_));
 sky130_as_sc_hs__and2_2 _43286_ (.A(_12526_),
    .B(_12527_),
    .Y(_12528_));
 sky130_as_sc_hs__nand2b_2 _43287_ (.B(_12440_),
    .Y(_12529_),
    .A(_12436_));
 sky130_as_sc_hs__or2_2 _43289_ (.A(_12528_),
    .B(_12529_),
    .Y(_12531_));
 sky130_as_sc_hs__nor2_2 _43292_ (.A(_12349_),
    .B(_12533_),
    .Y(_12534_));
 sky130_as_sc_hs__or2_2 _43293_ (.A(_05505_),
    .B(_12534_),
    .Y(_12535_));
 sky130_as_sc_hs__or2_2 _43295_ (.A(_12532_),
    .B(_12535_),
    .Y(_12537_));
 sky130_as_sc_hs__nand3_2 _43296_ (.A(net141),
    .B(_12536_),
    .C(_12537_),
    .Y(_12538_));
 sky130_as_sc_hs__nor2_2 _43297_ (.A(_05489_),
    .B(_05505_),
    .Y(_12539_));
 sky130_as_sc_hs__or2_2 _43299_ (.A(_05499_),
    .B(_12539_),
    .Y(_12541_));
 sky130_as_sc_hs__nand3_2 _43300_ (.A(net138),
    .B(_12540_),
    .C(_12541_),
    .Y(_12542_));
 sky130_as_sc_hs__or2_2 _43301_ (.A(\tholin_riscv.div_res[29] ),
    .B(_12463_),
    .Y(_12543_));
 sky130_as_sc_hs__and2_2 _43302_ (.A(net415),
    .B(_12543_),
    .Y(_12544_));
 sky130_as_sc_hs__or2_2 _43304_ (.A(\tholin_riscv.div_res[30] ),
    .B(_12544_),
    .Y(_12546_));
 sky130_as_sc_hs__nand3_2 _43305_ (.A(net111),
    .B(_12545_),
    .C(_12546_),
    .Y(_12547_));
 sky130_as_sc_hs__or2_2 _43306_ (.A(\tholin_riscv.div_shifter[61] ),
    .B(_12468_),
    .Y(_12548_));
 sky130_as_sc_hs__and2_2 _43307_ (.A(_21655_),
    .B(_12548_),
    .Y(_12549_));
 sky130_as_sc_hs__or2_2 _43309_ (.A(\tholin_riscv.div_shifter[62] ),
    .B(_12549_),
    .Y(_12551_));
 sky130_as_sc_hs__nand3_2 _43310_ (.A(net107),
    .B(_12550_),
    .C(_12551_),
    .Y(_12552_));
 sky130_as_sc_hs__and2_2 _43311_ (.A(_05968_),
    .B(_06433_),
    .Y(_12553_));
 sky130_as_sc_hs__or2_2 _43313_ (.A(_05536_),
    .B(_06539_),
    .Y(_12555_));
 sky130_as_sc_hs__and2_2 _43314_ (.A(_05534_),
    .B(_06160_),
    .Y(_12556_));
 sky130_as_sc_hs__or2_2 _43315_ (.A(_05535_),
    .B(_06158_),
    .Y(_12557_));
 sky130_as_sc_hs__and2_2 _43316_ (.A(\tholin_riscv.div_res[30] ),
    .B(_06564_),
    .Y(_12558_));
 sky130_as_sc_hs__nor2_2 _43318_ (.A(net119),
    .B(_12558_),
    .Y(_12560_));
 sky130_as_sc_hs__nand3_2 _43319_ (.A(_12557_),
    .B(_12559_),
    .C(_12560_),
    .Y(_12561_));
 sky130_as_sc_hs__nor2_2 _43320_ (.A(_12556_),
    .B(_12561_),
    .Y(_12562_));
 sky130_as_sc_hs__nand3_2 _43321_ (.A(_12554_),
    .B(_12555_),
    .C(_12562_),
    .Y(_12563_));
 sky130_as_sc_hs__nor2_2 _43322_ (.A(_12553_),
    .B(_12563_),
    .Y(_12564_));
 sky130_as_sc_hs__and2_2 _43323_ (.A(_12552_),
    .B(_12564_),
    .Y(_12565_));
 sky130_as_sc_hs__and2_2 _43324_ (.A(_12547_),
    .B(_12565_),
    .Y(_12566_));
 sky130_as_sc_hs__nand3_2 _43325_ (.A(_12538_),
    .B(_12542_),
    .C(_12566_),
    .Y(_12567_));
 sky130_as_sc_hs__or2_2 _43327_ (.A(_05536_),
    .B(_12568_),
    .Y(_12569_));
 sky130_as_sc_hs__and2_2 _43330_ (.A(_05543_),
    .B(_12571_),
    .Y(_12572_));
 sky130_as_sc_hs__or2_2 _43331_ (.A(_05536_),
    .B(_12572_),
    .Y(_12573_));
 sky130_as_sc_hs__and2_2 _43333_ (.A(_12573_),
    .B(_12574_),
    .Y(_12575_));
 sky130_as_sc_hs__nand3_2 _43334_ (.A(_06527_),
    .B(_12569_),
    .C(_12570_),
    .Y(_12576_));
 sky130_as_sc_hs__nand3_2 _43336_ (.A(net119),
    .B(_12576_),
    .C(_12577_),
    .Y(_12578_));
 sky130_as_sc_hs__or2_2 _43342_ (.A(\tholin_riscv.PC[30] ),
    .B(\tholin_riscv.Bimm[10] ),
    .Y(_12584_));
 sky130_as_sc_hs__or2_2 _43344_ (.A(_12582_),
    .B(_12585_),
    .Y(_12586_));
 sky130_as_sc_hs__nand3_2 _43346_ (.A(_06914_),
    .B(_12586_),
    .C(_12587_),
    .Y(_12588_));
 sky130_as_sc_hs__and2_2 _43347_ (.A(\tholin_riscv.PC[30] ),
    .B(_12497_),
    .Y(_12589_));
 sky130_as_sc_hs__nor2_2 _43348_ (.A(\tholin_riscv.PC[30] ),
    .B(_12497_),
    .Y(_12590_));
 sky130_as_sc_hs__nor2_2 _43349_ (.A(_12589_),
    .B(_12590_),
    .Y(_12591_));
 sky130_as_sc_hs__or2_2 _43350_ (.A(_21572_),
    .B(_12591_),
    .Y(_12592_));
 sky130_as_sc_hs__or2_2 _43351_ (.A(\tholin_riscv.Bimm[10] ),
    .B(_21590_),
    .Y(_12593_));
 sky130_as_sc_hs__nand3_2 _43352_ (.A(_12588_),
    .B(_12592_),
    .C(_12593_),
    .Y(_12594_));
 sky130_as_sc_hs__nand3_2 _43354_ (.A(_21546_),
    .B(_12580_),
    .C(_12595_),
    .Y(_12596_));
 sky130_as_sc_hs__and2_2 _43355_ (.A(\tholin_riscv.Bimm[10] ),
    .B(net371),
    .Y(_12597_));
 sky130_as_sc_hs__or2_2 _43356_ (.A(_10352_),
    .B(_12597_),
    .Y(_12598_));
 sky130_as_sc_hs__and2_2 _43362_ (.A(net334),
    .B(\tholin_riscv.io_size[1] ),
    .Y(_12603_));
 sky130_as_sc_hs__or2_2 _43363_ (.A(_10352_),
    .B(_12603_),
    .Y(_12604_));
 sky130_as_sc_hs__and2_2 _43365_ (.A(_12526_),
    .B(_12530_),
    .Y(_12606_));
 sky130_as_sc_hs__and2_2 _43366_ (.A(_12512_),
    .B(_12516_),
    .Y(_12607_));
 sky130_as_sc_hs__nand3_2 _43367_ (.A(_12519_),
    .B(_12523_),
    .C(_12607_),
    .Y(_12608_));
 sky130_as_sc_hs__or2_2 _43369_ (.A(_12606_),
    .B(_12608_),
    .Y(_12610_));
 sky130_as_sc_hs__and2_2 _43372_ (.A(_05504_),
    .B(_12612_),
    .Y(_12613_));
 sky130_as_sc_hs__or2_2 _43374_ (.A(_12611_),
    .B(_12613_),
    .Y(_12615_));
 sky130_as_sc_hs__nand3_2 _43375_ (.A(net142),
    .B(_12614_),
    .C(_12615_),
    .Y(_12616_));
 sky130_as_sc_hs__nor2b_2 _43376_ (.A(_05534_),
    .Y(_12617_),
    .B(_12573_));
 sky130_as_sc_hs__or2_2 _43377_ (.A(_05526_),
    .B(_12617_),
    .Y(_12618_));
 sky130_as_sc_hs__nor2b_2 _43381_ (.A(_05533_),
    .Y(_12622_),
    .B(_12570_));
 sky130_as_sc_hs__or2_2 _43382_ (.A(_05526_),
    .B(_12622_),
    .Y(_12623_));
 sky130_as_sc_hs__nand3_2 _43383_ (.A(_05917_),
    .B(_06527_),
    .C(_12623_),
    .Y(_12624_));
 sky130_as_sc_hs__nand3_2 _43384_ (.A(net119),
    .B(_12621_),
    .C(_12624_),
    .Y(_12625_));
 sky130_as_sc_hs__nor2_2 _43385_ (.A(_05498_),
    .B(_05505_),
    .Y(_12626_));
 sky130_as_sc_hs__nor2_2 _43386_ (.A(_12539_),
    .B(_12626_),
    .Y(_12627_));
 sky130_as_sc_hs__or2_2 _43387_ (.A(_05496_),
    .B(_12627_),
    .Y(_12628_));
 sky130_as_sc_hs__nand3_2 _43389_ (.A(net139),
    .B(_12628_),
    .C(_12629_),
    .Y(_12630_));
 sky130_as_sc_hs__or2_2 _43390_ (.A(\tholin_riscv.div_shifter[62] ),
    .B(_12548_),
    .Y(_12631_));
 sky130_as_sc_hs__and2_2 _43391_ (.A(_21655_),
    .B(_12631_),
    .Y(_12632_));
 sky130_as_sc_hs__or2_2 _43393_ (.A(\tholin_riscv.div_shifter[63] ),
    .B(_12632_),
    .Y(_12634_));
 sky130_as_sc_hs__nand3_2 _43394_ (.A(net109),
    .B(_12633_),
    .C(_12634_),
    .Y(_12635_));
 sky130_as_sc_hs__or2_2 _43395_ (.A(\tholin_riscv.div_res[30] ),
    .B(_12543_),
    .Y(_12636_));
 sky130_as_sc_hs__and2_2 _43396_ (.A(net415),
    .B(_12636_),
    .Y(_12637_));
 sky130_as_sc_hs__or2_2 _43398_ (.A(\tholin_riscv.div_res[31] ),
    .B(_12637_),
    .Y(_12639_));
 sky130_as_sc_hs__nand3_2 _43399_ (.A(net111),
    .B(_12638_),
    .C(_12639_),
    .Y(_12640_));
 sky130_as_sc_hs__and2_2 _43400_ (.A(_05965_),
    .B(_05968_),
    .Y(_12641_));
 sky130_as_sc_hs__or2_2 _43402_ (.A(_05526_),
    .B(_06539_),
    .Y(_12643_));
 sky130_as_sc_hs__nor2_2 _43403_ (.A(_05524_),
    .B(_06158_),
    .Y(_12644_));
 sky130_as_sc_hs__nand3_2 _43407_ (.A(net413),
    .B(_12646_),
    .C(_12647_),
    .Y(_12648_));
 sky130_as_sc_hs__nor2_2 _43408_ (.A(_12644_),
    .B(_12648_),
    .Y(_12649_));
 sky130_as_sc_hs__nand3_2 _43409_ (.A(_12643_),
    .B(_12645_),
    .C(_12649_),
    .Y(_12650_));
 sky130_as_sc_hs__nor2_2 _43410_ (.A(_12641_),
    .B(_12650_),
    .Y(_12651_));
 sky130_as_sc_hs__and2_2 _43411_ (.A(_12642_),
    .B(_12651_),
    .Y(_12652_));
 sky130_as_sc_hs__and2_2 _43412_ (.A(_12640_),
    .B(_12652_),
    .Y(_12653_));
 sky130_as_sc_hs__and2_2 _43413_ (.A(_12635_),
    .B(_12653_),
    .Y(_12654_));
 sky130_as_sc_hs__and2_2 _43414_ (.A(_12630_),
    .B(_12654_),
    .Y(_12655_));
 sky130_as_sc_hs__nand3_2 _43415_ (.A(_12616_),
    .B(_12625_),
    .C(_12655_),
    .Y(_12656_));
 sky130_as_sc_hs__and2_2 _43417_ (.A(_12583_),
    .B(_12657_),
    .Y(_12658_));
 sky130_as_sc_hs__or2_2 _43418_ (.A(\tholin_riscv.PC[31] ),
    .B(net334),
    .Y(_12659_));
 sky130_as_sc_hs__and2_2 _43420_ (.A(_12659_),
    .B(_12660_),
    .Y(_12661_));
 sky130_as_sc_hs__and2_2 _43421_ (.A(_12658_),
    .B(_12661_),
    .Y(_12662_));
 sky130_as_sc_hs__or2_2 _43422_ (.A(_12658_),
    .B(_12661_),
    .Y(_12663_));
 sky130_as_sc_hs__or2_2 _43424_ (.A(_12662_),
    .B(_12664_),
    .Y(_12665_));
 sky130_as_sc_hs__or2_2 _43425_ (.A(net334),
    .B(_21590_),
    .Y(_12666_));
 sky130_as_sc_hs__or2_2 _43426_ (.A(\tholin_riscv.PC[31] ),
    .B(_12589_),
    .Y(_12667_));
 sky130_as_sc_hs__and2_2 _43428_ (.A(_12667_),
    .B(_12668_),
    .Y(_12669_));
 sky130_as_sc_hs__or2_2 _43429_ (.A(_21572_),
    .B(_12669_),
    .Y(_12670_));
 sky130_as_sc_hs__nand3_2 _43430_ (.A(_12665_),
    .B(_12666_),
    .C(_12670_),
    .Y(_12671_));
 sky130_as_sc_hs__nand3_2 _43432_ (.A(_21546_),
    .B(_12656_),
    .C(_12672_),
    .Y(_12673_));
 sky130_as_sc_hs__and2_2 _43437_ (.A(_21549_),
    .B(_21554_),
    .Y(_12677_));
 sky130_as_sc_hs__and2_2 _43438_ (.A(_21559_),
    .B(_12677_),
    .Y(_12678_));
 sky130_as_sc_hs__and2_2 _43439_ (.A(_21576_),
    .B(_21579_),
    .Y(_12679_));
 sky130_as_sc_hs__and2_2 _43440_ (.A(_21584_),
    .B(_12679_),
    .Y(_12680_));
 sky130_as_sc_hs__and2_2 _43441_ (.A(_12678_),
    .B(_12680_),
    .Y(_12681_));
 sky130_as_sc_hs__or2_2 _43444_ (.A(net711),
    .B(_12681_),
    .Y(_12684_));
 sky130_as_sc_hs__and2_2 _43445_ (.A(_12683_),
    .B(net712),
    .Y(_00053_));
 sky130_as_sc_hs__and2_2 _43539_ (.A(_21550_),
    .B(_21553_),
    .Y(_12747_));
 sky130_as_sc_hs__and2_2 _43540_ (.A(_21558_),
    .B(_12747_),
    .Y(_12748_));
 sky130_as_sc_hs__and2_2 _43541_ (.A(_21580_),
    .B(_21584_),
    .Y(_12749_));
 sky130_as_sc_hs__and2_2 _43542_ (.A(_12748_),
    .B(_12749_),
    .Y(_12750_));
 sky130_as_sc_hs__or2_2 _43545_ (.A(net738),
    .B(_12750_),
    .Y(_12753_));
 sky130_as_sc_hs__and2_2 _43546_ (.A(_12752_),
    .B(net739),
    .Y(_00085_));
 sky130_as_sc_hs__and2_2 _43640_ (.A(_21559_),
    .B(_12747_),
    .Y(_12816_));
 sky130_as_sc_hs__and2_2 _43641_ (.A(_21585_),
    .B(_12816_),
    .Y(_12817_));
 sky130_as_sc_hs__or2_2 _43644_ (.A(net690),
    .B(_12817_),
    .Y(_12820_));
 sky130_as_sc_hs__and2_2 _43645_ (.A(_12819_),
    .B(net691),
    .Y(_00117_));
 sky130_as_sc_hs__and2_2 _43739_ (.A(_12680_),
    .B(_12816_),
    .Y(_12883_));
 sky130_as_sc_hs__or2_2 _43742_ (.A(net702),
    .B(_12883_),
    .Y(_12886_));
 sky130_as_sc_hs__and2_2 _43743_ (.A(_12885_),
    .B(net703),
    .Y(_00149_));
 sky130_as_sc_hs__and2_2 _43837_ (.A(_21558_),
    .B(_12677_),
    .Y(_12949_));
 sky130_as_sc_hs__and2_2 _43838_ (.A(_12680_),
    .B(_12949_),
    .Y(_12950_));
 sky130_as_sc_hs__or2_2 _43841_ (.A(net654),
    .B(_12950_),
    .Y(_12953_));
 sky130_as_sc_hs__and2_2 _43842_ (.A(_12952_),
    .B(net655),
    .Y(_00181_));
 sky130_as_sc_hs__nand3_2 _43937_ (.A(_19486_),
    .B(_05917_),
    .C(_05918_),
    .Y(_13017_));
 sky130_as_sc_hs__and2_2 _43938_ (.A(_13016_),
    .B(_13017_),
    .Y(_13018_));
 sky130_as_sc_hs__or2_2 _43939_ (.A(\tholin_riscv.Jimm[12] ),
    .B(_13018_),
    .Y(_13019_));
 sky130_as_sc_hs__nand3_2 _43941_ (.A(net411),
    .B(_13019_),
    .C(_13020_),
    .Y(_13021_));
 sky130_as_sc_hs__nor2_2 _43942_ (.A(_05914_),
    .B(_06155_),
    .Y(_13022_));
 sky130_as_sc_hs__nand3_2 _43943_ (.A(_05824_),
    .B(_05836_),
    .C(_13022_),
    .Y(_13023_));
 sky130_as_sc_hs__and2_2 _43944_ (.A(_05795_),
    .B(_05810_),
    .Y(_13024_));
 sky130_as_sc_hs__and2_2 _43945_ (.A(_05757_),
    .B(_05768_),
    .Y(_13025_));
 sky130_as_sc_hs__nand3_2 _43946_ (.A(_05726_),
    .B(_05738_),
    .C(_13025_),
    .Y(_13026_));
 sky130_as_sc_hs__nand3_2 _43947_ (.A(_05780_),
    .B(_05865_),
    .C(_05901_),
    .Y(_13027_));
 sky130_as_sc_hs__nor2_2 _43948_ (.A(_13026_),
    .B(_13027_),
    .Y(_13028_));
 sky130_as_sc_hs__and2_2 _43949_ (.A(_13024_),
    .B(_13028_),
    .Y(_13029_));
 sky130_as_sc_hs__and2_2 _43950_ (.A(_05565_),
    .B(_05574_),
    .Y(_13030_));
 sky130_as_sc_hs__nand3_2 _43951_ (.A(_05583_),
    .B(_05599_),
    .C(_13030_),
    .Y(_13031_));
 sky130_as_sc_hs__and2_2 _43952_ (.A(_05609_),
    .B(_05619_),
    .Y(_13032_));
 sky130_as_sc_hs__nand3_2 _43953_ (.A(_05629_),
    .B(_05639_),
    .C(_13032_),
    .Y(_13033_));
 sky130_as_sc_hs__nor2_2 _43954_ (.A(_13031_),
    .B(_13033_),
    .Y(_13034_));
 sky130_as_sc_hs__and2_2 _43955_ (.A(_05686_),
    .B(_05696_),
    .Y(_13035_));
 sky130_as_sc_hs__nand3_2 _43956_ (.A(_05706_),
    .B(_05715_),
    .C(_13035_),
    .Y(_13036_));
 sky130_as_sc_hs__and2_2 _43957_ (.A(_05666_),
    .B(_05676_),
    .Y(_13037_));
 sky130_as_sc_hs__nand3_2 _43958_ (.A(_05649_),
    .B(_05658_),
    .C(_13037_),
    .Y(_13038_));
 sky130_as_sc_hs__nor2_2 _43959_ (.A(_13036_),
    .B(_13038_),
    .Y(_13039_));
 sky130_as_sc_hs__nand3_2 _43960_ (.A(_13029_),
    .B(_13034_),
    .C(_13039_),
    .Y(_13040_));
 sky130_as_sc_hs__nor2_2 _43961_ (.A(_13023_),
    .B(_13040_),
    .Y(_13041_));
 sky130_as_sc_hs__or2_2 _43962_ (.A(_23602_),
    .B(_13041_),
    .Y(_13042_));
 sky130_as_sc_hs__nand2b_2 _43963_ (.B(_13041_),
    .Y(_13043_),
    .A(_23605_));
 sky130_as_sc_hs__nand3_2 _43964_ (.A(_13021_),
    .B(_13042_),
    .C(_13043_),
    .Y(_13044_));
 sky130_as_sc_hs__or2_2 _43968_ (.A(\tholin_riscv.Bimm[1] ),
    .B(net127),
    .Y(_13048_));
 sky130_as_sc_hs__and2_2 _43969_ (.A(_13047_),
    .B(_13048_),
    .Y(_13049_));
 sky130_as_sc_hs__or2_2 _43970_ (.A(\tholin_riscv.PC[1] ),
    .B(_13049_),
    .Y(_13050_));
 sky130_as_sc_hs__nand3_2 _43972_ (.A(_13046_),
    .B(_13050_),
    .C(_13051_),
    .Y(_13052_));
 sky130_as_sc_hs__and2_2 _43973_ (.A(_19477_),
    .B(\tholin_riscv.Bimm[6] ),
    .Y(_13053_));
 sky130_as_sc_hs__and2_2 _43974_ (.A(\tholin_riscv.Bimm[5] ),
    .B(_19478_),
    .Y(_13054_));
 sky130_as_sc_hs__and2_2 _43975_ (.A(_13053_),
    .B(_13054_),
    .Y(_13055_));
 sky130_as_sc_hs__nand3_2 _43976_ (.A(\tholin_riscv.Bimm[9] ),
    .B(_19476_),
    .C(_19981_),
    .Y(_13056_));
 sky130_as_sc_hs__and2_2 _43977_ (.A(\tholin_riscv.Iimm[2] ),
    .B(\tholin_riscv.Iimm[0] ),
    .Y(_13057_));
 sky130_as_sc_hs__and2_2 _43978_ (.A(\tholin_riscv.Iimm[3] ),
    .B(_19480_),
    .Y(_13058_));
 sky130_as_sc_hs__nor2_2 _43980_ (.A(_13056_),
    .B(_13059_),
    .Y(_13060_));
 sky130_as_sc_hs__and2_2 _43981_ (.A(_13055_),
    .B(_13060_),
    .Y(_13061_));
 sky130_as_sc_hs__nand3_2 _43983_ (.A(\tholin_riscv.PCE[1] ),
    .B(net135),
    .C(net125),
    .Y(_13063_));
 sky130_as_sc_hs__nor2_2 _43984_ (.A(\tholin_riscv.instr[3] ),
    .B(_19948_),
    .Y(_13064_));
 sky130_as_sc_hs__or2_2 _43985_ (.A(\tholin_riscv.instr[3] ),
    .B(_19948_),
    .Y(_13065_));
 sky130_as_sc_hs__or2_2 _43986_ (.A(_06526_),
    .B(_13065_),
    .Y(_13066_));
 sky130_as_sc_hs__nand3_2 _43987_ (.A(_13052_),
    .B(_13063_),
    .C(_13066_),
    .Y(_13067_));
 sky130_as_sc_hs__nand3_2 _43989_ (.A(_19942_),
    .B(_19991_),
    .C(_13062_),
    .Y(_13069_));
 sky130_as_sc_hs__and2_2 _43990_ (.A(_19944_),
    .B(_13069_),
    .Y(_13070_));
 sky130_as_sc_hs__or2_2 _43991_ (.A(\tholin_riscv.instr[4] ),
    .B(_13044_),
    .Y(_13071_));
 sky130_as_sc_hs__nor2_2 _43993_ (.A(_19949_),
    .B(_19987_),
    .Y(_13073_));
 sky130_as_sc_hs__and2_2 _43995_ (.A(_13070_),
    .B(_13074_),
    .Y(_13075_));
 sky130_as_sc_hs__nand3_2 _43997_ (.A(_13068_),
    .B(_13075_),
    .C(_13076_),
    .Y(_13077_));
 sky130_as_sc_hs__or2_2 _43998_ (.A(net1642),
    .B(_13075_),
    .Y(_13078_));
 sky130_as_sc_hs__and2_2 _43999_ (.A(net502),
    .B(net1643),
    .Y(_13079_));
 sky130_as_sc_hs__and2_2 _44000_ (.A(_13077_),
    .B(_13079_),
    .Y(_00213_));
 sky130_as_sc_hs__and2_2 _44001_ (.A(_12678_),
    .B(_12749_),
    .Y(_13080_));
 sky130_as_sc_hs__or2_2 _44004_ (.A(net729),
    .B(_13080_),
    .Y(_13083_));
 sky130_as_sc_hs__and2_2 _44005_ (.A(_13082_),
    .B(net730),
    .Y(_00214_));
 sky130_as_sc_hs__and2_2 _44099_ (.A(_21583_),
    .B(_12679_),
    .Y(_13146_));
 sky130_as_sc_hs__and2_2 _44100_ (.A(_12678_),
    .B(_13146_),
    .Y(_13147_));
 sky130_as_sc_hs__or2_2 _44103_ (.A(net666),
    .B(_13147_),
    .Y(_13150_));
 sky130_as_sc_hs__and2_2 _44104_ (.A(_13149_),
    .B(net667),
    .Y(_00246_));
 sky130_as_sc_hs__and2_2 _44198_ (.A(_21585_),
    .B(_12748_),
    .Y(_13213_));
 sky130_as_sc_hs__or2_2 _44201_ (.A(net687),
    .B(_13213_),
    .Y(_13216_));
 sky130_as_sc_hs__and2_2 _44202_ (.A(_13215_),
    .B(net688),
    .Y(_00278_));
 sky130_as_sc_hs__and2_2 _44296_ (.A(_12748_),
    .B(_13146_),
    .Y(_13279_));
 sky130_as_sc_hs__or2_2 _44299_ (.A(net651),
    .B(_13279_),
    .Y(_13282_));
 sky130_as_sc_hs__and2_2 _44300_ (.A(_13281_),
    .B(net652),
    .Y(_00310_));
 sky130_as_sc_hs__and2_2 _44394_ (.A(_12680_),
    .B(_12748_),
    .Y(_13345_));
 sky130_as_sc_hs__or2_2 _44397_ (.A(net696),
    .B(_13345_),
    .Y(_13348_));
 sky130_as_sc_hs__and2_2 _44398_ (.A(_13347_),
    .B(net697),
    .Y(_00342_));
 sky130_as_sc_hs__and2_2 _44492_ (.A(_12749_),
    .B(_12816_),
    .Y(_13411_));
 sky130_as_sc_hs__or2_2 _44495_ (.A(net705),
    .B(_13411_),
    .Y(_13414_));
 sky130_as_sc_hs__and2_2 _44496_ (.A(_13413_),
    .B(net706),
    .Y(_00374_));
 sky130_as_sc_hs__and2_2 _44590_ (.A(_21550_),
    .B(_21554_),
    .Y(_13477_));
 sky130_as_sc_hs__and2_2 _44591_ (.A(_21559_),
    .B(_13477_),
    .Y(_13478_));
 sky130_as_sc_hs__and2_2 _44592_ (.A(_12680_),
    .B(_13478_),
    .Y(_13479_));
 sky130_as_sc_hs__and2_2 _44593_ (.A(_06178_),
    .B(net77),
    .Y(_00406_));
 sky130_as_sc_hs__and2_2 _44594_ (.A(_06580_),
    .B(net77),
    .Y(_00407_));
 sky130_as_sc_hs__and2_2 _44595_ (.A(_06920_),
    .B(net77),
    .Y(_00408_));
 sky130_as_sc_hs__and2_2 _44596_ (.A(_07253_),
    .B(net77),
    .Y(_00409_));
 sky130_as_sc_hs__and2_2 _44597_ (.A(_07562_),
    .B(net77),
    .Y(_00410_));
 sky130_as_sc_hs__and2_2 _44598_ (.A(_07854_),
    .B(net77),
    .Y(_00411_));
 sky130_as_sc_hs__and2_2 _44599_ (.A(_08145_),
    .B(net77),
    .Y(_00412_));
 sky130_as_sc_hs__and2_2 _44600_ (.A(_08423_),
    .B(net76),
    .Y(_00413_));
 sky130_as_sc_hs__and2_2 _44601_ (.A(_08697_),
    .B(net76),
    .Y(_00414_));
 sky130_as_sc_hs__and2_2 _44602_ (.A(_08948_),
    .B(net76),
    .Y(_00415_));
 sky130_as_sc_hs__and2_2 _44603_ (.A(_09202_),
    .B(net76),
    .Y(_00416_));
 sky130_as_sc_hs__and2_2 _44604_ (.A(_09442_),
    .B(net76),
    .Y(_00417_));
 sky130_as_sc_hs__and2_2 _44605_ (.A(_09682_),
    .B(net76),
    .Y(_00418_));
 sky130_as_sc_hs__and2_2 _44606_ (.A(_09909_),
    .B(net76),
    .Y(_00419_));
 sky130_as_sc_hs__and2_2 _44607_ (.A(_10135_),
    .B(net77),
    .Y(_00420_));
 sky130_as_sc_hs__and2_2 _44608_ (.A(_10348_),
    .B(net77),
    .Y(_00421_));
 sky130_as_sc_hs__and2_2 _44609_ (.A(_10563_),
    .B(net76),
    .Y(_00422_));
 sky130_as_sc_hs__and2_2 _44610_ (.A(_10754_),
    .B(net76),
    .Y(_00423_));
 sky130_as_sc_hs__and2_2 _44611_ (.A(_10944_),
    .B(net76),
    .Y(_00424_));
 sky130_as_sc_hs__and2_2 _44612_ (.A(_11125_),
    .B(net77),
    .Y(_00425_));
 sky130_as_sc_hs__and2_2 _44613_ (.A(_11302_),
    .B(net77),
    .Y(_00426_));
 sky130_as_sc_hs__and2_2 _44614_ (.A(_11463_),
    .B(net76),
    .Y(_00427_));
 sky130_as_sc_hs__and2_2 _44615_ (.A(_11621_),
    .B(_13479_),
    .Y(_00428_));
 sky130_as_sc_hs__and2_2 _44616_ (.A(_11770_),
    .B(net77),
    .Y(_00429_));
 sky130_as_sc_hs__and2_2 _44617_ (.A(_11916_),
    .B(net76),
    .Y(_00430_));
 sky130_as_sc_hs__and2_2 _44618_ (.A(_12048_),
    .B(net77),
    .Y(_00431_));
 sky130_as_sc_hs__and2_2 _44619_ (.A(_12175_),
    .B(net76),
    .Y(_00432_));
 sky130_as_sc_hs__and2_2 _44620_ (.A(_12297_),
    .B(net76),
    .Y(_00433_));
 sky130_as_sc_hs__and2_2 _44621_ (.A(_12409_),
    .B(net76),
    .Y(_00434_));
 sky130_as_sc_hs__and2_2 _44622_ (.A(_12508_),
    .B(net76),
    .Y(_00435_));
 sky130_as_sc_hs__and2_2 _44623_ (.A(_12600_),
    .B(net77),
    .Y(_00436_));
 sky130_as_sc_hs__and2_2 _44624_ (.A(_12674_),
    .B(net77),
    .Y(_00437_));
 sky130_as_sc_hs__and2_2 _44625_ (.A(_21558_),
    .B(_13477_),
    .Y(_13480_));
 sky130_as_sc_hs__and2_2 _44626_ (.A(_21585_),
    .B(_13480_),
    .Y(_13481_));
 sky130_as_sc_hs__or2_2 _44629_ (.A(net681),
    .B(_13481_),
    .Y(_13484_));
 sky130_as_sc_hs__and2_2 _44630_ (.A(_13483_),
    .B(net682),
    .Y(_00438_));
 sky130_as_sc_hs__nand3_2 _44725_ (.A(\tholin_riscv.PCE[0] ),
    .B(net136),
    .C(net125),
    .Y(_13548_));
 sky130_as_sc_hs__or2_2 _44729_ (.A(_19991_),
    .B(_13551_),
    .Y(_13552_));
 sky130_as_sc_hs__and2_2 _44730_ (.A(_13070_),
    .B(_13552_),
    .Y(_13553_));
 sky130_as_sc_hs__nand3_2 _44732_ (.A(_13550_),
    .B(_13553_),
    .C(_13554_),
    .Y(_13555_));
 sky130_as_sc_hs__or2_2 _44733_ (.A(net1630),
    .B(_13553_),
    .Y(_13556_));
 sky130_as_sc_hs__and2_2 _44734_ (.A(net502),
    .B(net1631),
    .Y(_13557_));
 sky130_as_sc_hs__and2_2 _44735_ (.A(_13555_),
    .B(_13557_),
    .Y(_00470_));
 sky130_as_sc_hs__and2_2 _44736_ (.A(_12749_),
    .B(_13480_),
    .Y(_13558_));
 sky130_as_sc_hs__or2_2 _44739_ (.A(net693),
    .B(_13558_),
    .Y(_13561_));
 sky130_as_sc_hs__and2_2 _44740_ (.A(_13560_),
    .B(net694),
    .Y(_00471_));
 sky130_as_sc_hs__and2_2 _44834_ (.A(_21560_),
    .B(_12749_),
    .Y(_13624_));
 sky130_as_sc_hs__or2_2 _44837_ (.A(net684),
    .B(_13624_),
    .Y(_13627_));
 sky130_as_sc_hs__and2_2 _44838_ (.A(_13626_),
    .B(net685),
    .Y(_00503_));
 sky130_as_sc_hs__and2_2 _44932_ (.A(_12749_),
    .B(_13478_),
    .Y(_13690_));
 sky130_as_sc_hs__or2_2 _44935_ (.A(net708),
    .B(_13690_),
    .Y(_13693_));
 sky130_as_sc_hs__and2_2 _44936_ (.A(_13692_),
    .B(net709),
    .Y(_00535_));
 sky130_as_sc_hs__and2_2 _45030_ (.A(_21560_),
    .B(_12680_),
    .Y(_13756_));
 sky130_as_sc_hs__or2_2 _45033_ (.A(net660),
    .B(_13756_),
    .Y(_13759_));
 sky130_as_sc_hs__and2_2 _45034_ (.A(_13758_),
    .B(net661),
    .Y(_00567_));
 sky130_as_sc_hs__and2_2 _45128_ (.A(_21555_),
    .B(_21559_),
    .Y(_13822_));
 sky130_as_sc_hs__and2_2 _45129_ (.A(_21585_),
    .B(_13822_),
    .Y(_13823_));
 sky130_as_sc_hs__or2_2 _45132_ (.A(net741),
    .B(_13823_),
    .Y(_13826_));
 sky130_as_sc_hs__and2_2 _45133_ (.A(_13825_),
    .B(net742),
    .Y(_00599_));
 sky130_as_sc_hs__and2_2 _45227_ (.A(_12749_),
    .B(_13822_),
    .Y(_13889_));
 sky130_as_sc_hs__or2_2 _45230_ (.A(net732),
    .B(_13889_),
    .Y(_13892_));
 sky130_as_sc_hs__and2_2 _45231_ (.A(_13891_),
    .B(net733),
    .Y(_00631_));
 sky130_as_sc_hs__and2_2 _45325_ (.A(_13146_),
    .B(_13822_),
    .Y(_13955_));
 sky130_as_sc_hs__or2_2 _45328_ (.A(net657),
    .B(_13955_),
    .Y(_13958_));
 sky130_as_sc_hs__and2_2 _45329_ (.A(_13957_),
    .B(net658),
    .Y(_00663_));
 sky130_as_sc_hs__and2_2 _45423_ (.A(_12680_),
    .B(_13822_),
    .Y(_14021_));
 sky130_as_sc_hs__or2_2 _45426_ (.A(net663),
    .B(_14021_),
    .Y(_14024_));
 sky130_as_sc_hs__and2_2 _45427_ (.A(_14023_),
    .B(net664),
    .Y(_00695_));
 sky130_as_sc_hs__and2_2 _45521_ (.A(_21585_),
    .B(_12949_),
    .Y(_14087_));
 sky130_as_sc_hs__or2_2 _45524_ (.A(net714),
    .B(_14087_),
    .Y(_14090_));
 sky130_as_sc_hs__and2_2 _45525_ (.A(_14089_),
    .B(net715),
    .Y(_00727_));
 sky130_as_sc_hs__and2_2 _45619_ (.A(_12749_),
    .B(_12949_),
    .Y(_14153_));
 sky130_as_sc_hs__or2_2 _45622_ (.A(net699),
    .B(_14153_),
    .Y(_14156_));
 sky130_as_sc_hs__and2_2 _45623_ (.A(_14155_),
    .B(net700),
    .Y(_00759_));
 sky130_as_sc_hs__and2_2 _45717_ (.A(_12949_),
    .B(_13146_),
    .Y(_14219_));
 sky130_as_sc_hs__or2_2 _45720_ (.A(net672),
    .B(_14219_),
    .Y(_14222_));
 sky130_as_sc_hs__and2_2 _45721_ (.A(_14221_),
    .B(net673),
    .Y(_00791_));
 sky130_as_sc_hs__and2_2 _45815_ (.A(_13146_),
    .B(_13480_),
    .Y(_14285_));
 sky130_as_sc_hs__or2_2 _45818_ (.A(net720),
    .B(_14285_),
    .Y(_14288_));
 sky130_as_sc_hs__and2_2 _45819_ (.A(_14287_),
    .B(net721),
    .Y(_00823_));
 sky130_as_sc_hs__and2_2 _45913_ (.A(_21585_),
    .B(_12678_),
    .Y(_14351_));
 sky130_as_sc_hs__or2_2 _45916_ (.A(net726),
    .B(_14351_),
    .Y(_14354_));
 sky130_as_sc_hs__and2_2 _45917_ (.A(_14353_),
    .B(net727),
    .Y(_00855_));
 sky130_as_sc_hs__and2_2 _46011_ (.A(_12680_),
    .B(_13480_),
    .Y(_14417_));
 sky130_as_sc_hs__or2_2 _46014_ (.A(net744),
    .B(_14417_),
    .Y(_14420_));
 sky130_as_sc_hs__and2_2 _46015_ (.A(_14419_),
    .B(net745),
    .Y(_00887_));
 sky130_as_sc_hs__and2_2 _46109_ (.A(_21585_),
    .B(_13478_),
    .Y(_14483_));
 sky130_as_sc_hs__or2_2 _46112_ (.A(net675),
    .B(_14483_),
    .Y(_14486_));
 sky130_as_sc_hs__and2_2 _46113_ (.A(_14485_),
    .B(net676),
    .Y(_00919_));
 sky130_as_sc_hs__or2_2 _46214_ (.A(_19513_),
    .B(\tholin_riscv.uart.receive_div_counter[3] ),
    .Y(_14556_));
 sky130_as_sc_hs__nor2_2 _46215_ (.A(_19514_),
    .B(\tholin_riscv.uart.receive_div_counter[2] ),
    .Y(_14557_));
 sky130_as_sc_hs__or2_2 _46216_ (.A(_19506_),
    .B(\tholin_riscv.uart.receive_div_counter[10] ),
    .Y(_14558_));
 sky130_as_sc_hs__or2_2 _46219_ (.A(_19505_),
    .B(\tholin_riscv.uart.receive_div_counter[12] ),
    .Y(_14561_));
 sky130_as_sc_hs__or2_2 _46220_ (.A(_19512_),
    .B(\tholin_riscv.uart.receive_div_counter[4] ),
    .Y(_14562_));
 sky130_as_sc_hs__nor2_2 _46223_ (.A(_19511_),
    .B(\tholin_riscv.uart.receive_div_counter[5] ),
    .Y(_14565_));
 sky130_as_sc_hs__nor2_2 _46224_ (.A(_19503_),
    .B(\tholin_riscv.uart.receive_div_counter[14] ),
    .Y(_14566_));
 sky130_as_sc_hs__nor2_2 _46225_ (.A(_14565_),
    .B(_14566_),
    .Y(_14567_));
 sky130_as_sc_hs__or2_2 _46228_ (.A(\tholin_riscv.uart.divisor[11] ),
    .B(\tholin_riscv.uart.receive_div_counter[11] ),
    .Y(_14570_));
 sky130_as_sc_hs__and2_2 _46233_ (.A(_14573_),
    .B(_14574_),
    .Y(_14575_));
 sky130_as_sc_hs__or2_2 _46234_ (.A(_19507_),
    .B(\tholin_riscv.uart.receive_div_counter[9] ),
    .Y(_14576_));
 sky130_as_sc_hs__or2_2 _46236_ (.A(_19509_),
    .B(\tholin_riscv.uart.receive_div_counter[7] ),
    .Y(_14578_));
 sky130_as_sc_hs__nor2_2 _46237_ (.A(_19508_),
    .B(\tholin_riscv.uart.receive_div_counter[8] ),
    .Y(_14579_));
 sky130_as_sc_hs__nor2_2 _46239_ (.A(_19510_),
    .B(\tholin_riscv.uart.receive_div_counter[6] ),
    .Y(_14581_));
 sky130_as_sc_hs__nand3_2 _46240_ (.A(_14553_),
    .B(_14567_),
    .C(_14576_),
    .Y(_14582_));
 sky130_as_sc_hs__and2_2 _46241_ (.A(_14555_),
    .B(_14577_),
    .Y(_14583_));
 sky130_as_sc_hs__nand3_2 _46242_ (.A(_14564_),
    .B(_14580_),
    .C(_14583_),
    .Y(_14584_));
 sky130_as_sc_hs__nor2_2 _46243_ (.A(_14582_),
    .B(_14584_),
    .Y(_14585_));
 sky130_as_sc_hs__nor2_2 _46244_ (.A(_14579_),
    .B(_14581_),
    .Y(_14586_));
 sky130_as_sc_hs__and2_2 _46245_ (.A(_14549_),
    .B(_14578_),
    .Y(_14587_));
 sky130_as_sc_hs__and2_2 _46247_ (.A(_14561_),
    .B(_14588_),
    .Y(_14589_));
 sky130_as_sc_hs__nor2_2 _46248_ (.A(_19504_),
    .B(\tholin_riscv.uart.receive_div_counter[13] ),
    .Y(_14590_));
 sky130_as_sc_hs__nor2_2 _46249_ (.A(_14557_),
    .B(_14590_),
    .Y(_14591_));
 sky130_as_sc_hs__nand3_2 _46250_ (.A(_14559_),
    .B(_14562_),
    .C(_14589_),
    .Y(_14592_));
 sky130_as_sc_hs__nand3_2 _46251_ (.A(_14551_),
    .B(_14563_),
    .C(_14591_),
    .Y(_14593_));
 sky130_as_sc_hs__nor2_2 _46252_ (.A(_14592_),
    .B(_14593_),
    .Y(_14594_));
 sky130_as_sc_hs__nand3_2 _46253_ (.A(_14558_),
    .B(_14560_),
    .C(_14575_),
    .Y(_14595_));
 sky130_as_sc_hs__nand3_2 _46254_ (.A(_14550_),
    .B(_14568_),
    .C(_14587_),
    .Y(_14596_));
 sky130_as_sc_hs__nor2_2 _46255_ (.A(_14595_),
    .B(_14596_),
    .Y(_14597_));
 sky130_as_sc_hs__and2_2 _46256_ (.A(_14594_),
    .B(_14597_),
    .Y(_14598_));
 sky130_as_sc_hs__nand3_2 _46257_ (.A(_14554_),
    .B(_14556_),
    .C(_14586_),
    .Y(_14599_));
 sky130_as_sc_hs__nand3_2 _46258_ (.A(_14552_),
    .B(_14569_),
    .C(_14572_),
    .Y(_14600_));
 sky130_as_sc_hs__nor2_2 _46259_ (.A(_14599_),
    .B(_14600_),
    .Y(_14601_));
 sky130_as_sc_hs__nand3_2 _46260_ (.A(_14585_),
    .B(_14598_),
    .C(_14601_),
    .Y(_14602_));
 sky130_as_sc_hs__nor2_2 _46261_ (.A(_19531_),
    .B(_14602_),
    .Y(_14603_));
 sky130_as_sc_hs__or2_2 _46263_ (.A(\tholin_riscv.uart.receiving ),
    .B(net12),
    .Y(_14605_));
 sky130_as_sc_hs__or2_2 _46265_ (.A(_14603_),
    .B(_14606_),
    .Y(_14607_));
 sky130_as_sc_hs__and2_2 _46267_ (.A(net521),
    .B(_14608_),
    .Y(_00951_));
 sky130_as_sc_hs__or2_2 _46270_ (.A(_14604_),
    .B(_14609_),
    .Y(_14611_));
 sky130_as_sc_hs__and2_2 _46271_ (.A(net521),
    .B(_14610_),
    .Y(_14612_));
 sky130_as_sc_hs__and2_2 _46272_ (.A(_14611_),
    .B(_14612_),
    .Y(_00952_));
 sky130_as_sc_hs__nor2_2 _46273_ (.A(\tholin_riscv.uart.receive_counter[0] ),
    .B(\tholin_riscv.uart.receive_counter[1] ),
    .Y(_14613_));
 sky130_as_sc_hs__or2_2 _46277_ (.A(_14614_),
    .B(_14615_),
    .Y(_14617_));
 sky130_as_sc_hs__and2_2 _46278_ (.A(net525),
    .B(_14616_),
    .Y(_14618_));
 sky130_as_sc_hs__and2_2 _46279_ (.A(_14617_),
    .B(_14618_),
    .Y(_00953_));
 sky130_as_sc_hs__nor2_2 _46280_ (.A(net1699),
    .B(_14614_),
    .Y(_14619_));
 sky130_as_sc_hs__or2_2 _46283_ (.A(_14619_),
    .B(_14620_),
    .Y(_14622_));
 sky130_as_sc_hs__and2_2 _46284_ (.A(net525),
    .B(_14622_),
    .Y(_14623_));
 sky130_as_sc_hs__and2_2 _46285_ (.A(_14621_),
    .B(_14623_),
    .Y(_00954_));
 sky130_as_sc_hs__or2_2 _46286_ (.A(\tholin_riscv.uart.counter[1] ),
    .B(\tholin_riscv.uart.counter[0] ),
    .Y(_14624_));
 sky130_as_sc_hs__or2_2 _46287_ (.A(net621),
    .B(\tholin_riscv.uart.counter[2] ),
    .Y(_14625_));
 sky130_as_sc_hs__or2_2 _46288_ (.A(_14624_),
    .B(_14625_),
    .Y(_14626_));
 sky130_as_sc_hs__nor2_2 _46289_ (.A(\tholin_riscv.requested_addr[1] ),
    .B(\tholin_riscv.requested_addr[0] ),
    .Y(_14627_));
 sky130_as_sc_hs__and2_2 _46290_ (.A(_19901_),
    .B(_14627_),
    .Y(_14628_));
 sky130_as_sc_hs__and2_2 _46291_ (.A(_20731_),
    .B(_14628_),
    .Y(_14629_));
 sky130_as_sc_hs__nor2_2 _46293_ (.A(_14626_),
    .B(_14629_),
    .Y(_14631_));
 sky130_as_sc_hs__and2_2 _46294_ (.A(net1647),
    .B(_14631_),
    .Y(_14632_));
 sky130_as_sc_hs__or2_2 _46296_ (.A(_19502_),
    .B(\tholin_riscv.uart.div_counter[15] ),
    .Y(_14634_));
 sky130_as_sc_hs__or2_2 _46302_ (.A(_19513_),
    .B(\tholin_riscv.uart.div_counter[3] ),
    .Y(_14640_));
 sky130_as_sc_hs__nor2_2 _46303_ (.A(_19514_),
    .B(\tholin_riscv.uart.div_counter[2] ),
    .Y(_14641_));
 sky130_as_sc_hs__or2_2 _46304_ (.A(_19506_),
    .B(\tholin_riscv.uart.div_counter[10] ),
    .Y(_14642_));
 sky130_as_sc_hs__or2_2 _46307_ (.A(_19505_),
    .B(\tholin_riscv.uart.div_counter[12] ),
    .Y(_14645_));
 sky130_as_sc_hs__or2_2 _46308_ (.A(_19512_),
    .B(\tholin_riscv.uart.div_counter[4] ),
    .Y(_14646_));
 sky130_as_sc_hs__nor2_2 _46311_ (.A(_19511_),
    .B(\tholin_riscv.uart.div_counter[5] ),
    .Y(_14649_));
 sky130_as_sc_hs__nor2_2 _46312_ (.A(_19503_),
    .B(\tholin_riscv.uart.div_counter[14] ),
    .Y(_14650_));
 sky130_as_sc_hs__nor2_2 _46313_ (.A(_14649_),
    .B(_14650_),
    .Y(_14651_));
 sky130_as_sc_hs__or2_2 _46316_ (.A(\tholin_riscv.uart.divisor[11] ),
    .B(\tholin_riscv.uart.div_counter[11] ),
    .Y(_14654_));
 sky130_as_sc_hs__and2_2 _46321_ (.A(_14657_),
    .B(_14658_),
    .Y(_14659_));
 sky130_as_sc_hs__or2_2 _46322_ (.A(_19507_),
    .B(\tholin_riscv.uart.div_counter[9] ),
    .Y(_14660_));
 sky130_as_sc_hs__or2_2 _46324_ (.A(_19509_),
    .B(\tholin_riscv.uart.div_counter[7] ),
    .Y(_14662_));
 sky130_as_sc_hs__nor2_2 _46325_ (.A(_19508_),
    .B(\tholin_riscv.uart.div_counter[8] ),
    .Y(_14663_));
 sky130_as_sc_hs__or2_2 _46326_ (.A(_19516_),
    .B(\tholin_riscv.uart.div_counter[0] ),
    .Y(_14664_));
 sky130_as_sc_hs__nor2_2 _46327_ (.A(_19510_),
    .B(\tholin_riscv.uart.div_counter[6] ),
    .Y(_14665_));
 sky130_as_sc_hs__nand3_2 _46328_ (.A(_14637_),
    .B(_14651_),
    .C(_14660_),
    .Y(_14666_));
 sky130_as_sc_hs__and2_2 _46329_ (.A(_14639_),
    .B(_14661_),
    .Y(_14667_));
 sky130_as_sc_hs__nand3_2 _46330_ (.A(_14648_),
    .B(_14664_),
    .C(_14667_),
    .Y(_14668_));
 sky130_as_sc_hs__nor2_2 _46331_ (.A(_14666_),
    .B(_14668_),
    .Y(_14669_));
 sky130_as_sc_hs__nor2_2 _46332_ (.A(_14663_),
    .B(_14665_),
    .Y(_14670_));
 sky130_as_sc_hs__and2_2 _46333_ (.A(_14633_),
    .B(_14662_),
    .Y(_14671_));
 sky130_as_sc_hs__and2_2 _46335_ (.A(_14645_),
    .B(_14672_),
    .Y(_14673_));
 sky130_as_sc_hs__nor2_2 _46336_ (.A(_19504_),
    .B(\tholin_riscv.uart.div_counter[13] ),
    .Y(_14674_));
 sky130_as_sc_hs__nor2_2 _46337_ (.A(_14641_),
    .B(_14674_),
    .Y(_14675_));
 sky130_as_sc_hs__nand3_2 _46338_ (.A(_14643_),
    .B(_14646_),
    .C(_14673_),
    .Y(_14676_));
 sky130_as_sc_hs__nand3_2 _46339_ (.A(_14635_),
    .B(_14647_),
    .C(_14675_),
    .Y(_14677_));
 sky130_as_sc_hs__nor2_2 _46340_ (.A(_14676_),
    .B(_14677_),
    .Y(_14678_));
 sky130_as_sc_hs__nand3_2 _46341_ (.A(_14642_),
    .B(_14644_),
    .C(_14659_),
    .Y(_14679_));
 sky130_as_sc_hs__nand3_2 _46342_ (.A(_14634_),
    .B(_14652_),
    .C(_14671_),
    .Y(_14680_));
 sky130_as_sc_hs__nor2_2 _46343_ (.A(_14679_),
    .B(_14680_),
    .Y(_14681_));
 sky130_as_sc_hs__and2_2 _46344_ (.A(_14678_),
    .B(_14681_),
    .Y(_14682_));
 sky130_as_sc_hs__nand3_2 _46345_ (.A(_14638_),
    .B(_14640_),
    .C(_14670_),
    .Y(_14683_));
 sky130_as_sc_hs__nand3_2 _46346_ (.A(_14636_),
    .B(_14653_),
    .C(_14656_),
    .Y(_14684_));
 sky130_as_sc_hs__nor2_2 _46347_ (.A(_14683_),
    .B(_14684_),
    .Y(_14685_));
 sky130_as_sc_hs__and2_2 _46348_ (.A(_14669_),
    .B(_14685_),
    .Y(_14686_));
 sky130_as_sc_hs__and2_2 _46349_ (.A(_14682_),
    .B(_14686_),
    .Y(_14687_));
 sky130_as_sc_hs__inv_2 _46350_ (.Y(_14688_),
    .A(_14687_));
 sky130_as_sc_hs__nor2_2 _46352_ (.A(net1647),
    .B(_14689_),
    .Y(_14690_));
 sky130_as_sc_hs__or2_2 _46353_ (.A(net1648),
    .B(_14690_),
    .Y(_14691_));
 sky130_as_sc_hs__and2_2 _46354_ (.A(net518),
    .B(net1649),
    .Y(_00955_));
 sky130_as_sc_hs__or2_2 _46355_ (.A(_14631_),
    .B(_14690_),
    .Y(_14692_));
 sky130_as_sc_hs__or2_2 _46358_ (.A(_14689_),
    .B(_14694_),
    .Y(_14695_));
 sky130_as_sc_hs__and2_2 _46360_ (.A(net518),
    .B(_14696_),
    .Y(_00956_));
 sky130_as_sc_hs__and2_2 _46362_ (.A(\tholin_riscv.uart.div_counter[1] ),
    .B(\tholin_riscv.uart.div_counter[0] ),
    .Y(_14698_));
 sky130_as_sc_hs__and2_2 _46363_ (.A(\tholin_riscv.uart.div_counter[2] ),
    .B(_14698_),
    .Y(_14699_));
 sky130_as_sc_hs__nor2_2 _46364_ (.A(\tholin_riscv.uart.div_counter[2] ),
    .B(_14698_),
    .Y(_14700_));
 sky130_as_sc_hs__or2_2 _46365_ (.A(_14699_),
    .B(_14700_),
    .Y(_14701_));
 sky130_as_sc_hs__or2_2 _46366_ (.A(_14689_),
    .B(_14701_),
    .Y(_14702_));
 sky130_as_sc_hs__and2_2 _46368_ (.A(net521),
    .B(_14703_),
    .Y(_00957_));
 sky130_as_sc_hs__nor2_2 _46370_ (.A(\tholin_riscv.uart.div_counter[3] ),
    .B(_14699_),
    .Y(_14705_));
 sky130_as_sc_hs__and2_2 _46371_ (.A(\tholin_riscv.uart.div_counter[3] ),
    .B(_14699_),
    .Y(_14706_));
 sky130_as_sc_hs__or2_2 _46372_ (.A(_14705_),
    .B(_14706_),
    .Y(_14707_));
 sky130_as_sc_hs__or2_2 _46373_ (.A(_14689_),
    .B(_14707_),
    .Y(_14708_));
 sky130_as_sc_hs__and2_2 _46375_ (.A(net521),
    .B(_14709_),
    .Y(_00958_));
 sky130_as_sc_hs__and2_2 _46377_ (.A(\tholin_riscv.uart.div_counter[4] ),
    .B(_14706_),
    .Y(_14711_));
 sky130_as_sc_hs__nor2_2 _46378_ (.A(\tholin_riscv.uart.div_counter[4] ),
    .B(_14706_),
    .Y(_14712_));
 sky130_as_sc_hs__or2_2 _46379_ (.A(_14711_),
    .B(_14712_),
    .Y(_14713_));
 sky130_as_sc_hs__or2_2 _46380_ (.A(_14689_),
    .B(_14713_),
    .Y(_14714_));
 sky130_as_sc_hs__and2_2 _46382_ (.A(net521),
    .B(_14715_),
    .Y(_00959_));
 sky130_as_sc_hs__and2_2 _46384_ (.A(\tholin_riscv.uart.div_counter[5] ),
    .B(_14711_),
    .Y(_14717_));
 sky130_as_sc_hs__nor2_2 _46385_ (.A(\tholin_riscv.uart.div_counter[5] ),
    .B(_14711_),
    .Y(_14718_));
 sky130_as_sc_hs__or2_2 _46386_ (.A(_14717_),
    .B(_14718_),
    .Y(_14719_));
 sky130_as_sc_hs__or2_2 _46387_ (.A(_14689_),
    .B(_14719_),
    .Y(_14720_));
 sky130_as_sc_hs__and2_2 _46389_ (.A(net521),
    .B(_14721_),
    .Y(_00960_));
 sky130_as_sc_hs__and2_2 _46391_ (.A(\tholin_riscv.uart.div_counter[6] ),
    .B(_14717_),
    .Y(_14723_));
 sky130_as_sc_hs__nor2_2 _46392_ (.A(\tholin_riscv.uart.div_counter[6] ),
    .B(_14717_),
    .Y(_14724_));
 sky130_as_sc_hs__or2_2 _46393_ (.A(_14723_),
    .B(_14724_),
    .Y(_14725_));
 sky130_as_sc_hs__or2_2 _46394_ (.A(_14689_),
    .B(_14725_),
    .Y(_14726_));
 sky130_as_sc_hs__and2_2 _46396_ (.A(net521),
    .B(_14727_),
    .Y(_00961_));
 sky130_as_sc_hs__and2_2 _46397_ (.A(\tholin_riscv.uart.div_counter[7] ),
    .B(_14723_),
    .Y(_14728_));
 sky130_as_sc_hs__nor2_2 _46398_ (.A(_14689_),
    .B(_14728_),
    .Y(_14729_));
 sky130_as_sc_hs__or2_2 _46399_ (.A(_14631_),
    .B(_14729_),
    .Y(_14730_));
 sky130_as_sc_hs__and2_2 _46403_ (.A(net519),
    .B(_14733_),
    .Y(_00962_));
 sky130_as_sc_hs__nor2_2 _46405_ (.A(\tholin_riscv.uart.div_counter[8] ),
    .B(_14689_),
    .Y(_14735_));
 sky130_as_sc_hs__and2_2 _46408_ (.A(net521),
    .B(_14737_),
    .Y(_00963_));
 sky130_as_sc_hs__and2_2 _46410_ (.A(\tholin_riscv.uart.div_counter[8] ),
    .B(_14728_),
    .Y(_14739_));
 sky130_as_sc_hs__and2_2 _46411_ (.A(\tholin_riscv.uart.div_counter[9] ),
    .B(_14739_),
    .Y(_14740_));
 sky130_as_sc_hs__or2_2 _46412_ (.A(_14689_),
    .B(_14740_),
    .Y(_14741_));
 sky130_as_sc_hs__or2_2 _46414_ (.A(net1626),
    .B(_14739_),
    .Y(_14743_));
 sky130_as_sc_hs__and2_2 _46415_ (.A(net519),
    .B(net1627),
    .Y(_14744_));
 sky130_as_sc_hs__and2_2 _46416_ (.A(_14742_),
    .B(_14744_),
    .Y(_00964_));
 sky130_as_sc_hs__and2_2 _46418_ (.A(\tholin_riscv.uart.div_counter[10] ),
    .B(_14740_),
    .Y(_14746_));
 sky130_as_sc_hs__or2_2 _46419_ (.A(_14689_),
    .B(_14746_),
    .Y(_14747_));
 sky130_as_sc_hs__or2_2 _46421_ (.A(net1624),
    .B(_14740_),
    .Y(_14749_));
 sky130_as_sc_hs__and2_2 _46422_ (.A(net519),
    .B(net1625),
    .Y(_14750_));
 sky130_as_sc_hs__and2_2 _46423_ (.A(_14748_),
    .B(_14750_),
    .Y(_00965_));
 sky130_as_sc_hs__and2_2 _46425_ (.A(\tholin_riscv.uart.div_counter[11] ),
    .B(_14746_),
    .Y(_14752_));
 sky130_as_sc_hs__or2_2 _46426_ (.A(_14689_),
    .B(_14752_),
    .Y(_14753_));
 sky130_as_sc_hs__or2_2 _46428_ (.A(net1620),
    .B(_14746_),
    .Y(_14755_));
 sky130_as_sc_hs__and2_2 _46429_ (.A(net519),
    .B(net1621),
    .Y(_14756_));
 sky130_as_sc_hs__and2_2 _46430_ (.A(_14754_),
    .B(_14756_),
    .Y(_00966_));
 sky130_as_sc_hs__and2_2 _46432_ (.A(net1607),
    .B(_14752_),
    .Y(_14758_));
 sky130_as_sc_hs__or2_2 _46433_ (.A(_14689_),
    .B(_14758_),
    .Y(_14759_));
 sky130_as_sc_hs__or2_2 _46435_ (.A(net1607),
    .B(_14752_),
    .Y(_14761_));
 sky130_as_sc_hs__and2_2 _46436_ (.A(net519),
    .B(net1608),
    .Y(_14762_));
 sky130_as_sc_hs__and2_2 _46437_ (.A(_14760_),
    .B(_14762_),
    .Y(_00967_));
 sky130_as_sc_hs__and2_2 _46439_ (.A(\tholin_riscv.uart.div_counter[13] ),
    .B(_14758_),
    .Y(_14764_));
 sky130_as_sc_hs__or2_2 _46440_ (.A(_14689_),
    .B(_14764_),
    .Y(_14765_));
 sky130_as_sc_hs__or2_2 _46442_ (.A(net1636),
    .B(_14758_),
    .Y(_14767_));
 sky130_as_sc_hs__and2_2 _46443_ (.A(net519),
    .B(net1637),
    .Y(_14768_));
 sky130_as_sc_hs__and2_2 _46444_ (.A(_14766_),
    .B(_14768_),
    .Y(_00968_));
 sky130_as_sc_hs__and2_2 _46445_ (.A(\tholin_riscv.uart.div_counter[14] ),
    .B(_14764_),
    .Y(_14769_));
 sky130_as_sc_hs__nor2_2 _46446_ (.A(_14689_),
    .B(_14769_),
    .Y(_14770_));
 sky130_as_sc_hs__or2_2 _46447_ (.A(_14631_),
    .B(_14770_),
    .Y(_14771_));
 sky130_as_sc_hs__and2_2 _46451_ (.A(net519),
    .B(_14774_),
    .Y(_00969_));
 sky130_as_sc_hs__nor2_2 _46453_ (.A(\tholin_riscv.uart.div_counter[15] ),
    .B(_14689_),
    .Y(_14776_));
 sky130_as_sc_hs__and2_2 _46456_ (.A(net516),
    .B(_14778_),
    .Y(_00970_));
 sky130_as_sc_hs__nor2_2 _46457_ (.A(\tholin_riscv.uart.receive_counter[3] ),
    .B(\tholin_riscv.uart.receive_counter[2] ),
    .Y(_14779_));
 sky130_as_sc_hs__and2_2 _46458_ (.A(_14613_),
    .B(_14779_),
    .Y(_14780_));
 sky130_as_sc_hs__and2_2 _46459_ (.A(_14603_),
    .B(_14780_),
    .Y(_14781_));
 sky130_as_sc_hs__or2_2 _46461_ (.A(net1750),
    .B(_14781_),
    .Y(_14783_));
 sky130_as_sc_hs__or2_2 _46462_ (.A(net605),
    .B(_14782_),
    .Y(_14784_));
 sky130_as_sc_hs__and2_2 _46463_ (.A(net525),
    .B(net1751),
    .Y(_14785_));
 sky130_as_sc_hs__and2_2 _46464_ (.A(net606),
    .B(_14785_),
    .Y(_00971_));
 sky130_as_sc_hs__or2_2 _46465_ (.A(net1759),
    .B(_14781_),
    .Y(_14786_));
 sky130_as_sc_hs__or2_2 _46466_ (.A(net593),
    .B(_14782_),
    .Y(_14787_));
 sky130_as_sc_hs__and2_2 _46467_ (.A(net525),
    .B(net1760),
    .Y(_14788_));
 sky130_as_sc_hs__and2_2 _46468_ (.A(net594),
    .B(_14788_),
    .Y(_00972_));
 sky130_as_sc_hs__or2_2 _46469_ (.A(net1753),
    .B(_14781_),
    .Y(_14789_));
 sky130_as_sc_hs__or2_2 _46470_ (.A(net587),
    .B(_14782_),
    .Y(_14790_));
 sky130_as_sc_hs__and2_2 _46471_ (.A(net525),
    .B(net1754),
    .Y(_14791_));
 sky130_as_sc_hs__and2_2 _46472_ (.A(net588),
    .B(_14791_),
    .Y(_00973_));
 sky130_as_sc_hs__or2_2 _46473_ (.A(net1747),
    .B(_14781_),
    .Y(_14792_));
 sky130_as_sc_hs__or2_2 _46474_ (.A(net575),
    .B(_14782_),
    .Y(_14793_));
 sky130_as_sc_hs__and2_2 _46475_ (.A(net525),
    .B(net1748),
    .Y(_14794_));
 sky130_as_sc_hs__and2_2 _46476_ (.A(net576),
    .B(_14794_),
    .Y(_00974_));
 sky130_as_sc_hs__or2_2 _46477_ (.A(\tholin_riscv.uart.dout[4] ),
    .B(_14781_),
    .Y(_14795_));
 sky130_as_sc_hs__or2_2 _46478_ (.A(net1724),
    .B(_14782_),
    .Y(_14796_));
 sky130_as_sc_hs__and2_2 _46479_ (.A(net525),
    .B(_14795_),
    .Y(_14797_));
 sky130_as_sc_hs__and2_2 _46480_ (.A(net555),
    .B(_14797_),
    .Y(_00975_));
 sky130_as_sc_hs__or2_2 _46481_ (.A(net1744),
    .B(_14781_),
    .Y(_14798_));
 sky130_as_sc_hs__or2_2 _46482_ (.A(net590),
    .B(_14782_),
    .Y(_14799_));
 sky130_as_sc_hs__and2_2 _46483_ (.A(net525),
    .B(net1745),
    .Y(_14800_));
 sky130_as_sc_hs__and2_2 _46484_ (.A(net591),
    .B(_14800_),
    .Y(_00976_));
 sky130_as_sc_hs__or2_2 _46485_ (.A(net1756),
    .B(_14781_),
    .Y(_14801_));
 sky130_as_sc_hs__or2_2 _46486_ (.A(net584),
    .B(_14782_),
    .Y(_14802_));
 sky130_as_sc_hs__and2_2 _46487_ (.A(net525),
    .B(net1757),
    .Y(_14803_));
 sky130_as_sc_hs__and2_2 _46488_ (.A(net585),
    .B(_14803_),
    .Y(_00977_));
 sky130_as_sc_hs__or2_2 _46489_ (.A(net1735),
    .B(_14781_),
    .Y(_14804_));
 sky130_as_sc_hs__or2_2 _46490_ (.A(net615),
    .B(_14782_),
    .Y(_14805_));
 sky130_as_sc_hs__and2_2 _46491_ (.A(net525),
    .B(net1736),
    .Y(_14806_));
 sky130_as_sc_hs__and2_2 _46492_ (.A(net567),
    .B(_14806_),
    .Y(_00978_));
 sky130_as_sc_hs__nand3_2 _46494_ (.A(\tholin_riscv.spi.counter[3] ),
    .B(\tholin_riscv.spi.counter[2] ),
    .C(\tholin_riscv.spi.counter[4] ),
    .Y(_14808_));
 sky130_as_sc_hs__nor2_2 _46495_ (.A(_14807_),
    .B(_14808_),
    .Y(_14809_));
 sky130_as_sc_hs__or2_2 _46496_ (.A(_14807_),
    .B(_14808_),
    .Y(_14810_));
 sky130_as_sc_hs__nand2b_2 _46497_ (.B(\tholin_riscv.spi.divisor[6] ),
    .Y(_14811_),
    .A(\tholin_riscv.spi.div_counter[6] ));
 sky130_as_sc_hs__nand2b_2 _46498_ (.B(\tholin_riscv.spi.div_counter[6] ),
    .Y(_14812_),
    .A(\tholin_riscv.spi.divisor[6] ));
 sky130_as_sc_hs__and2_2 _46499_ (.A(_14811_),
    .B(_14812_),
    .Y(_14813_));
 sky130_as_sc_hs__or2_2 _46501_ (.A(\tholin_riscv.spi.divisor[2] ),
    .B(_19520_),
    .Y(_14815_));
 sky130_as_sc_hs__nand3_2 _46502_ (.A(_14813_),
    .B(_14814_),
    .C(_14815_),
    .Y(_14816_));
 sky130_as_sc_hs__or2_2 _46503_ (.A(\tholin_riscv.spi.divisor[0] ),
    .B(_19522_),
    .Y(_14817_));
 sky130_as_sc_hs__nor2b_2 _46505_ (.A(\tholin_riscv.spi.divisor[3] ),
    .Y(_14819_),
    .B(\tholin_riscv.spi.div_counter[3] ));
 sky130_as_sc_hs__nand2b_2 _46506_ (.B(\tholin_riscv.spi.divisor[3] ),
    .Y(_14820_),
    .A(\tholin_riscv.spi.div_counter[3] ));
 sky130_as_sc_hs__or2_2 _46507_ (.A(\tholin_riscv.spi.divisor[5] ),
    .B(\tholin_riscv.spi.div_counter[5] ),
    .Y(_14821_));
 sky130_as_sc_hs__or2_2 _46510_ (.A(\tholin_riscv.spi.divisor[7] ),
    .B(\tholin_riscv.spi.div_counter[7] ),
    .Y(_14824_));
 sky130_as_sc_hs__or2_2 _46514_ (.A(\tholin_riscv.spi.divisor[1] ),
    .B(_19521_),
    .Y(_14828_));
 sky130_as_sc_hs__nor2_2 _46515_ (.A(\tholin_riscv.spi.divisor[4] ),
    .B(_19519_),
    .Y(_14829_));
 sky130_as_sc_hs__nand3_2 _46517_ (.A(_14823_),
    .B(_14827_),
    .C(_14828_),
    .Y(_14831_));
 sky130_as_sc_hs__nand3_2 _46518_ (.A(_14817_),
    .B(_14818_),
    .C(_14826_),
    .Y(_14832_));
 sky130_as_sc_hs__nor2_2 _46519_ (.A(_14831_),
    .B(_14832_),
    .Y(_14833_));
 sky130_as_sc_hs__nor2_2 _46520_ (.A(_14819_),
    .B(_14829_),
    .Y(_14834_));
 sky130_as_sc_hs__nand3_2 _46521_ (.A(_14820_),
    .B(_14830_),
    .C(_14834_),
    .Y(_14835_));
 sky130_as_sc_hs__nor2_2 _46522_ (.A(_14816_),
    .B(_14835_),
    .Y(_14836_));
 sky130_as_sc_hs__nor2_2 _46524_ (.A(_14809_),
    .B(_14837_),
    .Y(_14838_));
 sky130_as_sc_hs__and2_2 _46525_ (.A(\tholin_riscv.spi.counter[0] ),
    .B(_14838_),
    .Y(_14839_));
 sky130_as_sc_hs__and2_2 _46526_ (.A(_20738_),
    .B(_14628_),
    .Y(_14840_));
 sky130_as_sc_hs__nor2_2 _46528_ (.A(_14839_),
    .B(_14840_),
    .Y(_14842_));
 sky130_as_sc_hs__and2_2 _46531_ (.A(net526),
    .B(_14844_),
    .Y(_14845_));
 sky130_as_sc_hs__and2_2 _46532_ (.A(_14843_),
    .B(_14845_),
    .Y(_00979_));
 sky130_as_sc_hs__and2_2 _46536_ (.A(net504),
    .B(_14848_),
    .Y(_00980_));
 sky130_as_sc_hs__and2_2 _46540_ (.A(net504),
    .B(_14851_),
    .Y(_00981_));
 sky130_as_sc_hs__and2_2 _46544_ (.A(net516),
    .B(_14854_),
    .Y(_00982_));
 sky130_as_sc_hs__and2_2 _46548_ (.A(net516),
    .B(_14857_),
    .Y(_00983_));
 sky130_as_sc_hs__and2_2 _46552_ (.A(net500),
    .B(_14860_),
    .Y(_00984_));
 sky130_as_sc_hs__and2_2 _46556_ (.A(net519),
    .B(_14863_),
    .Y(_00985_));
 sky130_as_sc_hs__and2_2 _46560_ (.A(net519),
    .B(_14866_),
    .Y(_00986_));
 sky130_as_sc_hs__and2_2 _46561_ (.A(net518),
    .B(_14626_),
    .Y(_00988_));
 sky130_as_sc_hs__nand3_2 _46564_ (.A(_00988_),
    .B(_14867_),
    .C(_14868_),
    .Y(_00987_));
 sky130_as_sc_hs__and2_2 _46568_ (.A(net500),
    .B(_14871_),
    .Y(_00989_));
 sky130_as_sc_hs__and2_2 _46569_ (.A(_14626_),
    .B(_14687_),
    .Y(_14872_));
 sky130_as_sc_hs__inv_4 _46570_ (.Y(_14873_),
    .A(_14872_));
 sky130_as_sc_hs__nand3_2 _46572_ (.A(\tholin_riscv.uart.data_buff[0] ),
    .B(_14630_),
    .C(_14873_),
    .Y(_14875_));
 sky130_as_sc_hs__and2_2 _46574_ (.A(net516),
    .B(_14876_),
    .Y(_00990_));
 sky130_as_sc_hs__or2_2 _46575_ (.A(\tholin_riscv.uart.data_buff[1] ),
    .B(_14629_),
    .Y(_14877_));
 sky130_as_sc_hs__or2_2 _46576_ (.A(\tholin_riscv.instr[0] ),
    .B(_14630_),
    .Y(_14878_));
 sky130_as_sc_hs__nand3_2 _46577_ (.A(_14873_),
    .B(_14877_),
    .C(_14878_),
    .Y(_14879_));
 sky130_as_sc_hs__and2_2 _46580_ (.A(net516),
    .B(_14881_),
    .Y(_00991_));
 sky130_as_sc_hs__or2_2 _46581_ (.A(\tholin_riscv.uart.data_buff[2] ),
    .B(_14629_),
    .Y(_14882_));
 sky130_as_sc_hs__or2_2 _46582_ (.A(\tholin_riscv.instr[1] ),
    .B(_14630_),
    .Y(_14883_));
 sky130_as_sc_hs__nand3_2 _46583_ (.A(_14873_),
    .B(_14882_),
    .C(_14883_),
    .Y(_14884_));
 sky130_as_sc_hs__and2_2 _46586_ (.A(net516),
    .B(_14886_),
    .Y(_00992_));
 sky130_as_sc_hs__or2_2 _46587_ (.A(\tholin_riscv.uart.data_buff[3] ),
    .B(_14629_),
    .Y(_14887_));
 sky130_as_sc_hs__nand3_2 _46589_ (.A(_14873_),
    .B(_14887_),
    .C(_14888_),
    .Y(_14889_));
 sky130_as_sc_hs__and2_2 _46592_ (.A(net515),
    .B(_14891_),
    .Y(_00993_));
 sky130_as_sc_hs__or2_2 _46593_ (.A(\tholin_riscv.uart.data_buff[4] ),
    .B(_14629_),
    .Y(_14892_));
 sky130_as_sc_hs__nand3_2 _46595_ (.A(_14873_),
    .B(_14892_),
    .C(_14893_),
    .Y(_14894_));
 sky130_as_sc_hs__and2_2 _46598_ (.A(net515),
    .B(_14896_),
    .Y(_00994_));
 sky130_as_sc_hs__or2_2 _46599_ (.A(\tholin_riscv.uart.data_buff[5] ),
    .B(_14629_),
    .Y(_14897_));
 sky130_as_sc_hs__nand3_2 _46601_ (.A(_14873_),
    .B(_14897_),
    .C(_14898_),
    .Y(_14899_));
 sky130_as_sc_hs__and2_2 _46604_ (.A(net515),
    .B(_14901_),
    .Y(_00995_));
 sky130_as_sc_hs__or2_2 _46605_ (.A(\tholin_riscv.uart.data_buff[6] ),
    .B(_14629_),
    .Y(_14902_));
 sky130_as_sc_hs__nand3_2 _46607_ (.A(_14873_),
    .B(_14902_),
    .C(_14903_),
    .Y(_14904_));
 sky130_as_sc_hs__and2_2 _46610_ (.A(net515),
    .B(_14906_),
    .Y(_00996_));
 sky130_as_sc_hs__or2_2 _46611_ (.A(\tholin_riscv.uart.data_buff[7] ),
    .B(_14629_),
    .Y(_14907_));
 sky130_as_sc_hs__nand3_2 _46613_ (.A(_14873_),
    .B(_14907_),
    .C(_14908_),
    .Y(_14909_));
 sky130_as_sc_hs__and2_2 _46616_ (.A(net515),
    .B(_14911_),
    .Y(_00997_));
 sky130_as_sc_hs__or2_2 _46617_ (.A(\tholin_riscv.uart.data_buff[8] ),
    .B(_14629_),
    .Y(_14912_));
 sky130_as_sc_hs__or2_2 _46618_ (.A(\tholin_riscv.Bimm[11] ),
    .B(_14630_),
    .Y(_14913_));
 sky130_as_sc_hs__nand3_2 _46619_ (.A(_14873_),
    .B(_14912_),
    .C(_14913_),
    .Y(_14914_));
 sky130_as_sc_hs__and2_2 _46622_ (.A(net516),
    .B(_14916_),
    .Y(_00998_));
 sky130_as_sc_hs__or2_2 _46623_ (.A(net581),
    .B(_14629_),
    .Y(_14917_));
 sky130_as_sc_hs__nor2_2 _46624_ (.A(_19528_),
    .B(_14872_),
    .Y(_14918_));
 sky130_as_sc_hs__and2_2 _46625_ (.A(net582),
    .B(_14918_),
    .Y(_00999_));
 sky130_as_sc_hs__and2_2 _46628_ (.A(net1694),
    .B(_14687_),
    .Y(_14921_));
 sky130_as_sc_hs__inv_2 _46629_ (.Y(_14922_),
    .A(_14921_));
 sky130_as_sc_hs__and2_2 _46630_ (.A(_00988_),
    .B(_14922_),
    .Y(_14923_));
 sky130_as_sc_hs__and2_2 _46631_ (.A(_14920_),
    .B(_14923_),
    .Y(_01000_));
 sky130_as_sc_hs__and2_2 _46634_ (.A(_14922_),
    .B(_14925_),
    .Y(_14926_));
 sky130_as_sc_hs__or2_2 _46635_ (.A(net754),
    .B(_14926_),
    .Y(_14927_));
 sky130_as_sc_hs__nand3_2 _46636_ (.A(net754),
    .B(_19530_),
    .C(_14687_),
    .Y(_14928_));
 sky130_as_sc_hs__and2_2 _46637_ (.A(net518),
    .B(_14928_),
    .Y(_14929_));
 sky130_as_sc_hs__and2_2 _46638_ (.A(net755),
    .B(_14929_),
    .Y(_01001_));
 sky130_as_sc_hs__or2_2 _46639_ (.A(\tholin_riscv.uart.counter[2] ),
    .B(_14624_),
    .Y(_14930_));
 sky130_as_sc_hs__nand3_2 _46643_ (.A(\tholin_riscv.uart.counter[2] ),
    .B(_14630_),
    .C(_14688_),
    .Y(_14934_));
 sky130_as_sc_hs__and2_2 _46645_ (.A(_00988_),
    .B(_14935_),
    .Y(_01002_));
 sky130_as_sc_hs__or2_2 _46646_ (.A(net621),
    .B(_14629_),
    .Y(_14936_));
 sky130_as_sc_hs__and2_2 _46649_ (.A(net517),
    .B(_14938_),
    .Y(_14939_));
 sky130_as_sc_hs__and2_2 _46650_ (.A(net622),
    .B(_14939_),
    .Y(_01003_));
 sky130_as_sc_hs__and2_2 _46651_ (.A(_19531_),
    .B(net12),
    .Y(_14940_));
 sky130_as_sc_hs__nor2_2 _46652_ (.A(_19528_),
    .B(_14940_),
    .Y(_14941_));
 sky130_as_sc_hs__and2_2 _46653_ (.A(_14782_),
    .B(_14941_),
    .Y(_01004_));
 sky130_as_sc_hs__nor2_2 _46654_ (.A(_14602_),
    .B(_14780_),
    .Y(_14942_));
 sky130_as_sc_hs__and2_2 _46655_ (.A(\tholin_riscv.uart.receiving ),
    .B(_14942_),
    .Y(_14943_));
 sky130_as_sc_hs__nor2_2 _46657_ (.A(_19531_),
    .B(_14942_),
    .Y(_14945_));
 sky130_as_sc_hs__or2_2 _46658_ (.A(_14940_),
    .B(_14945_),
    .Y(_14946_));
 sky130_as_sc_hs__and2_2 _46661_ (.A(net525),
    .B(_14948_),
    .Y(_01005_));
 sky130_as_sc_hs__and2_2 _46665_ (.A(net526),
    .B(_14951_),
    .Y(_01006_));
 sky130_as_sc_hs__and2_2 _46669_ (.A(net525),
    .B(_14954_),
    .Y(_01007_));
 sky130_as_sc_hs__and2_2 _46673_ (.A(net525),
    .B(_14957_),
    .Y(_01008_));
 sky130_as_sc_hs__and2_2 _46677_ (.A(net526),
    .B(_14960_),
    .Y(_01009_));
 sky130_as_sc_hs__and2_2 _46681_ (.A(net525),
    .B(_14963_),
    .Y(_01010_));
 sky130_as_sc_hs__and2_2 _46685_ (.A(net525),
    .B(_14966_),
    .Y(_01011_));
 sky130_as_sc_hs__or2_2 _46686_ (.A(net615),
    .B(_14943_),
    .Y(_14967_));
 sky130_as_sc_hs__or2_2 _46687_ (.A(net12),
    .B(_14945_),
    .Y(_14968_));
 sky130_as_sc_hs__and2_2 _46688_ (.A(net525),
    .B(_14968_),
    .Y(_14969_));
 sky130_as_sc_hs__and2_2 _46689_ (.A(net616),
    .B(_14969_),
    .Y(_01012_));
 sky130_as_sc_hs__and2_2 _46690_ (.A(net1665),
    .B(_14940_),
    .Y(_14970_));
 sky130_as_sc_hs__and2_2 _46691_ (.A(\tholin_riscv.uart.receiving ),
    .B(_14602_),
    .Y(_14971_));
 sky130_as_sc_hs__and2_2 _46692_ (.A(_19525_),
    .B(_14971_),
    .Y(_14972_));
 sky130_as_sc_hs__or2_2 _46693_ (.A(net1666),
    .B(_14972_),
    .Y(_14973_));
 sky130_as_sc_hs__and2_2 _46694_ (.A(net521),
    .B(_14973_),
    .Y(_01013_));
 sky130_as_sc_hs__or2_2 _46695_ (.A(_14940_),
    .B(_14972_),
    .Y(_14974_));
 sky130_as_sc_hs__nand3_2 _46697_ (.A(_19524_),
    .B(\tholin_riscv.uart.receive_div_counter[0] ),
    .C(_14971_),
    .Y(_14976_));
 sky130_as_sc_hs__and2_2 _46699_ (.A(net521),
    .B(_14977_),
    .Y(_01014_));
 sky130_as_sc_hs__and2_2 _46701_ (.A(\tholin_riscv.uart.receive_div_counter[1] ),
    .B(\tholin_riscv.uart.receive_div_counter[0] ),
    .Y(_14979_));
 sky130_as_sc_hs__and2_2 _46702_ (.A(\tholin_riscv.uart.receive_div_counter[2] ),
    .B(_14979_),
    .Y(_14980_));
 sky130_as_sc_hs__nor2_2 _46703_ (.A(\tholin_riscv.uart.receive_div_counter[2] ),
    .B(_14979_),
    .Y(_14981_));
 sky130_as_sc_hs__nor2_2 _46704_ (.A(_14980_),
    .B(_14981_),
    .Y(_14982_));
 sky130_as_sc_hs__and2_2 _46707_ (.A(net521),
    .B(_14984_),
    .Y(_01015_));
 sky130_as_sc_hs__and2_2 _46709_ (.A(\tholin_riscv.uart.receive_div_counter[3] ),
    .B(_14980_),
    .Y(_14986_));
 sky130_as_sc_hs__nor2_2 _46710_ (.A(\tholin_riscv.uart.receive_div_counter[3] ),
    .B(_14980_),
    .Y(_14987_));
 sky130_as_sc_hs__nor2_2 _46711_ (.A(_14986_),
    .B(_14987_),
    .Y(_14988_));
 sky130_as_sc_hs__and2_2 _46714_ (.A(net521),
    .B(_14990_),
    .Y(_01016_));
 sky130_as_sc_hs__and2_2 _46716_ (.A(\tholin_riscv.uart.receive_div_counter[4] ),
    .B(_14986_),
    .Y(_14992_));
 sky130_as_sc_hs__nor2_2 _46717_ (.A(\tholin_riscv.uart.receive_div_counter[4] ),
    .B(_14986_),
    .Y(_14993_));
 sky130_as_sc_hs__nor2_2 _46718_ (.A(_14992_),
    .B(_14993_),
    .Y(_14994_));
 sky130_as_sc_hs__and2_2 _46721_ (.A(net521),
    .B(_14996_),
    .Y(_01017_));
 sky130_as_sc_hs__and2_2 _46723_ (.A(\tholin_riscv.uart.receive_div_counter[5] ),
    .B(_14992_),
    .Y(_14998_));
 sky130_as_sc_hs__nor2_2 _46724_ (.A(\tholin_riscv.uart.receive_div_counter[5] ),
    .B(_14992_),
    .Y(_14999_));
 sky130_as_sc_hs__nor2_2 _46725_ (.A(_14998_),
    .B(_14999_),
    .Y(_15000_));
 sky130_as_sc_hs__and2_2 _46728_ (.A(net522),
    .B(_15002_),
    .Y(_01018_));
 sky130_as_sc_hs__and2_2 _46730_ (.A(\tholin_riscv.uart.receive_div_counter[6] ),
    .B(_14998_),
    .Y(_15004_));
 sky130_as_sc_hs__nor2_2 _46731_ (.A(\tholin_riscv.uart.receive_div_counter[6] ),
    .B(_14998_),
    .Y(_15005_));
 sky130_as_sc_hs__nor2_2 _46732_ (.A(_15004_),
    .B(_15005_),
    .Y(_15006_));
 sky130_as_sc_hs__and2_2 _46735_ (.A(net521),
    .B(_15008_),
    .Y(_01019_));
 sky130_as_sc_hs__and2_2 _46737_ (.A(\tholin_riscv.uart.receive_div_counter[7] ),
    .B(_15004_),
    .Y(_15010_));
 sky130_as_sc_hs__or2_2 _46738_ (.A(\tholin_riscv.uart.receive_div_counter[7] ),
    .B(_15004_),
    .Y(_15011_));
 sky130_as_sc_hs__or2_2 _46740_ (.A(_15010_),
    .B(_15012_),
    .Y(_15013_));
 sky130_as_sc_hs__and2_2 _46742_ (.A(net520),
    .B(_15014_),
    .Y(_01020_));
 sky130_as_sc_hs__and2_2 _46744_ (.A(\tholin_riscv.uart.receive_div_counter[8] ),
    .B(_15010_),
    .Y(_15016_));
 sky130_as_sc_hs__or2_2 _46745_ (.A(\tholin_riscv.uart.receive_div_counter[8] ),
    .B(_15010_),
    .Y(_15017_));
 sky130_as_sc_hs__or2_2 _46747_ (.A(_15016_),
    .B(_15018_),
    .Y(_15019_));
 sky130_as_sc_hs__and2_2 _46749_ (.A(net521),
    .B(_15020_),
    .Y(_01021_));
 sky130_as_sc_hs__or2_2 _46751_ (.A(\tholin_riscv.uart.receive_div_counter[9] ),
    .B(_15016_),
    .Y(_15022_));
 sky130_as_sc_hs__and2_2 _46752_ (.A(\tholin_riscv.uart.receive_div_counter[9] ),
    .B(_15016_),
    .Y(_15023_));
 sky130_as_sc_hs__or2_2 _46754_ (.A(_15023_),
    .B(_15024_),
    .Y(_15025_));
 sky130_as_sc_hs__and2_2 _46756_ (.A(net520),
    .B(_15026_),
    .Y(_01022_));
 sky130_as_sc_hs__or2_2 _46758_ (.A(\tholin_riscv.uart.receive_div_counter[10] ),
    .B(_15023_),
    .Y(_15028_));
 sky130_as_sc_hs__and2_2 _46759_ (.A(\tholin_riscv.uart.receive_div_counter[10] ),
    .B(_15023_),
    .Y(_15029_));
 sky130_as_sc_hs__or2_2 _46761_ (.A(_15029_),
    .B(_15030_),
    .Y(_15031_));
 sky130_as_sc_hs__and2_2 _46763_ (.A(net520),
    .B(_15032_),
    .Y(_01023_));
 sky130_as_sc_hs__and2_2 _46765_ (.A(\tholin_riscv.uart.receive_div_counter[11] ),
    .B(_15029_),
    .Y(_15034_));
 sky130_as_sc_hs__or2_2 _46766_ (.A(\tholin_riscv.uart.receive_div_counter[11] ),
    .B(_15029_),
    .Y(_15035_));
 sky130_as_sc_hs__or2_2 _46768_ (.A(_15034_),
    .B(_15036_),
    .Y(_15037_));
 sky130_as_sc_hs__and2_2 _46770_ (.A(net519),
    .B(_15038_),
    .Y(_01024_));
 sky130_as_sc_hs__or2_2 _46772_ (.A(\tholin_riscv.uart.receive_div_counter[12] ),
    .B(_15034_),
    .Y(_15040_));
 sky130_as_sc_hs__and2_2 _46773_ (.A(\tholin_riscv.uart.receive_div_counter[12] ),
    .B(_15034_),
    .Y(_15041_));
 sky130_as_sc_hs__or2_2 _46775_ (.A(_15041_),
    .B(_15042_),
    .Y(_15043_));
 sky130_as_sc_hs__and2_2 _46777_ (.A(net520),
    .B(_15044_),
    .Y(_01025_));
 sky130_as_sc_hs__and2_2 _46779_ (.A(\tholin_riscv.uart.receive_div_counter[13] ),
    .B(_15041_),
    .Y(_15046_));
 sky130_as_sc_hs__or2_2 _46780_ (.A(\tholin_riscv.uart.receive_div_counter[13] ),
    .B(_15041_),
    .Y(_15047_));
 sky130_as_sc_hs__or2_2 _46782_ (.A(_15046_),
    .B(_15048_),
    .Y(_15049_));
 sky130_as_sc_hs__and2_2 _46784_ (.A(net520),
    .B(_15050_),
    .Y(_01026_));
 sky130_as_sc_hs__and2_2 _46785_ (.A(\tholin_riscv.uart.receive_div_counter[14] ),
    .B(_15046_),
    .Y(_15051_));
 sky130_as_sc_hs__nor2b_2 _46786_ (.A(_15051_),
    .Y(_15052_),
    .B(_14971_));
 sky130_as_sc_hs__or2_2 _46787_ (.A(_14940_),
    .B(_15052_),
    .Y(_15053_));
 sky130_as_sc_hs__and2_2 _46791_ (.A(net520),
    .B(_15056_),
    .Y(_01027_));
 sky130_as_sc_hs__nand3_2 _46793_ (.A(_19523_),
    .B(_14971_),
    .C(_15051_),
    .Y(_15058_));
 sky130_as_sc_hs__and2_2 _46795_ (.A(net520),
    .B(_15059_),
    .Y(_01028_));
 sky130_as_sc_hs__and2_2 _46796_ (.A(_14810_),
    .B(_14837_),
    .Y(_15060_));
 sky130_as_sc_hs__and2_2 _46797_ (.A(_19522_),
    .B(_15060_),
    .Y(_15061_));
 sky130_as_sc_hs__and2_2 _46798_ (.A(_14809_),
    .B(_14841_),
    .Y(_15062_));
 sky130_as_sc_hs__and2_2 _46799_ (.A(net1682),
    .B(_15062_),
    .Y(_15063_));
 sky130_as_sc_hs__or2_2 _46800_ (.A(_15061_),
    .B(_15063_),
    .Y(_15064_));
 sky130_as_sc_hs__and2_2 _46801_ (.A(net515),
    .B(_15064_),
    .Y(_01029_));
 sky130_as_sc_hs__or2_2 _46802_ (.A(_15061_),
    .B(_15062_),
    .Y(_15065_));
 sky130_as_sc_hs__nand3_2 _46804_ (.A(_19521_),
    .B(\tholin_riscv.spi.div_counter[0] ),
    .C(_15060_),
    .Y(_15067_));
 sky130_as_sc_hs__and2_2 _46806_ (.A(net515),
    .B(_15068_),
    .Y(_01030_));
 sky130_as_sc_hs__and2_2 _46808_ (.A(\tholin_riscv.spi.div_counter[1] ),
    .B(\tholin_riscv.spi.div_counter[0] ),
    .Y(_15070_));
 sky130_as_sc_hs__and2_2 _46809_ (.A(\tholin_riscv.spi.div_counter[2] ),
    .B(_15070_),
    .Y(_15071_));
 sky130_as_sc_hs__nor2_2 _46810_ (.A(\tholin_riscv.spi.div_counter[2] ),
    .B(_15070_),
    .Y(_15072_));
 sky130_as_sc_hs__nor2_2 _46811_ (.A(_15071_),
    .B(_15072_),
    .Y(_15073_));
 sky130_as_sc_hs__and2_2 _46814_ (.A(net511),
    .B(_15075_),
    .Y(_01031_));
 sky130_as_sc_hs__nor2_2 _46816_ (.A(\tholin_riscv.spi.div_counter[3] ),
    .B(_15071_),
    .Y(_15077_));
 sky130_as_sc_hs__and2_2 _46817_ (.A(\tholin_riscv.spi.div_counter[3] ),
    .B(_15071_),
    .Y(_15078_));
 sky130_as_sc_hs__nor2_2 _46818_ (.A(_15077_),
    .B(_15078_),
    .Y(_15079_));
 sky130_as_sc_hs__and2_2 _46821_ (.A(net511),
    .B(_15081_),
    .Y(_01032_));
 sky130_as_sc_hs__and2_2 _46823_ (.A(\tholin_riscv.spi.div_counter[4] ),
    .B(_15078_),
    .Y(_15083_));
 sky130_as_sc_hs__nor2_2 _46824_ (.A(\tholin_riscv.spi.div_counter[4] ),
    .B(_15078_),
    .Y(_15084_));
 sky130_as_sc_hs__nor2_2 _46825_ (.A(_15083_),
    .B(_15084_),
    .Y(_15085_));
 sky130_as_sc_hs__and2_2 _46828_ (.A(net515),
    .B(_15087_),
    .Y(_01033_));
 sky130_as_sc_hs__and2_2 _46830_ (.A(\tholin_riscv.spi.div_counter[5] ),
    .B(_15083_),
    .Y(_15089_));
 sky130_as_sc_hs__nor2_2 _46831_ (.A(\tholin_riscv.spi.div_counter[5] ),
    .B(_15083_),
    .Y(_15090_));
 sky130_as_sc_hs__nor2_2 _46832_ (.A(_15089_),
    .B(_15090_),
    .Y(_15091_));
 sky130_as_sc_hs__and2_2 _46835_ (.A(net515),
    .B(_15093_),
    .Y(_01034_));
 sky130_as_sc_hs__and2_2 _46837_ (.A(_15060_),
    .B(_15094_),
    .Y(_15095_));
 sky130_as_sc_hs__or2_2 _46838_ (.A(_15062_),
    .B(_15095_),
    .Y(_15096_));
 sky130_as_sc_hs__and2_2 _46842_ (.A(net511),
    .B(_15099_),
    .Y(_01035_));
 sky130_as_sc_hs__or2_2 _46845_ (.A(_15094_),
    .B(_15101_),
    .Y(_15102_));
 sky130_as_sc_hs__and2_2 _46847_ (.A(net515),
    .B(_15103_),
    .Y(_01036_));
 sky130_as_sc_hs__or2_2 _46848_ (.A(net1238),
    .B(_14809_),
    .Y(_15104_));
 sky130_as_sc_hs__and2_2 _46850_ (.A(net519),
    .B(net1239),
    .Y(_15106_));
 sky130_as_sc_hs__and2_2 _46851_ (.A(_15105_),
    .B(net1240),
    .Y(_01037_));
 sky130_as_sc_hs__or2_2 _46852_ (.A(net1765),
    .B(_14809_),
    .Y(_15107_));
 sky130_as_sc_hs__or2_2 _46853_ (.A(net569),
    .B(_14810_),
    .Y(_15108_));
 sky130_as_sc_hs__and2_2 _46854_ (.A(net519),
    .B(net1766),
    .Y(_15109_));
 sky130_as_sc_hs__and2_2 _46855_ (.A(net570),
    .B(_15109_),
    .Y(_01038_));
 sky130_as_sc_hs__or2_2 _46856_ (.A(net1737),
    .B(_14809_),
    .Y(_15110_));
 sky130_as_sc_hs__or2_2 _46857_ (.A(net572),
    .B(_14810_),
    .Y(_15111_));
 sky130_as_sc_hs__and2_2 _46858_ (.A(net519),
    .B(net1738),
    .Y(_15112_));
 sky130_as_sc_hs__and2_2 _46859_ (.A(net573),
    .B(_15112_),
    .Y(_01039_));
 sky130_as_sc_hs__or2_2 _46860_ (.A(\tholin_riscv.spi.dout[3] ),
    .B(_14809_),
    .Y(_15113_));
 sky130_as_sc_hs__or2_2 _46861_ (.A(net1732),
    .B(_14810_),
    .Y(_15114_));
 sky130_as_sc_hs__and2_2 _46862_ (.A(net516),
    .B(_15113_),
    .Y(_15115_));
 sky130_as_sc_hs__and2_2 _46863_ (.A(net561),
    .B(_15115_),
    .Y(_01040_));
 sky130_as_sc_hs__or2_2 _46864_ (.A(net1762),
    .B(_14809_),
    .Y(_15116_));
 sky130_as_sc_hs__or2_2 _46865_ (.A(net578),
    .B(_14810_),
    .Y(_15117_));
 sky130_as_sc_hs__and2_2 _46866_ (.A(net516),
    .B(net1763),
    .Y(_15118_));
 sky130_as_sc_hs__and2_2 _46867_ (.A(net579),
    .B(_15118_),
    .Y(_01041_));
 sky130_as_sc_hs__or2_2 _46868_ (.A(net1740),
    .B(_14809_),
    .Y(_15119_));
 sky130_as_sc_hs__or2_2 _46869_ (.A(net563),
    .B(_14810_),
    .Y(_15120_));
 sky130_as_sc_hs__and2_2 _46870_ (.A(net516),
    .B(net1741),
    .Y(_15121_));
 sky130_as_sc_hs__and2_2 _46871_ (.A(net564),
    .B(_15121_),
    .Y(_01042_));
 sky130_as_sc_hs__or2_2 _46872_ (.A(net1768),
    .B(_14809_),
    .Y(_15122_));
 sky130_as_sc_hs__or2_2 _46873_ (.A(net599),
    .B(_14810_),
    .Y(_15123_));
 sky130_as_sc_hs__and2_2 _46874_ (.A(net519),
    .B(net1769),
    .Y(_15124_));
 sky130_as_sc_hs__and2_2 _46875_ (.A(net600),
    .B(_15124_),
    .Y(_01043_));
 sky130_as_sc_hs__or2_2 _46876_ (.A(\tholin_riscv.spi.dout[7] ),
    .B(_14809_),
    .Y(_15125_));
 sky130_as_sc_hs__or2_2 _46877_ (.A(net1728),
    .B(_14810_),
    .Y(_15126_));
 sky130_as_sc_hs__and2_2 _46878_ (.A(net519),
    .B(_15125_),
    .Y(_15127_));
 sky130_as_sc_hs__and2_2 _46879_ (.A(net558),
    .B(_15127_),
    .Y(_01044_));
 sky130_as_sc_hs__nor2_2 _46880_ (.A(\tholin_riscv.spi.counter[0] ),
    .B(_14837_),
    .Y(_15128_));
 sky130_as_sc_hs__inv_4 _46881_ (.Y(_15129_),
    .A(_15128_));
 sky130_as_sc_hs__or2_2 _46882_ (.A(_14809_),
    .B(_15128_),
    .Y(_15130_));
 sky130_as_sc_hs__and2_2 _46885_ (.A(net516),
    .B(_14810_),
    .Y(_15133_));
 sky130_as_sc_hs__nand3_2 _46886_ (.A(\tholin_riscv.spi.data_out_buff[7] ),
    .B(_15128_),
    .C(_15133_),
    .Y(_15134_));
 sky130_as_sc_hs__nand3_2 _46891_ (.A(net516),
    .B(_14839_),
    .C(_15135_),
    .Y(_15138_));
 sky130_as_sc_hs__and2_2 _46893_ (.A(_19528_),
    .B(net608),
    .Y(_15139_));
 sky130_as_sc_hs__or2_2 _46894_ (.A(_15133_),
    .B(net609),
    .Y(_01047_));
 sky130_as_sc_hs__nor2_2 _46895_ (.A(_14838_),
    .B(_14840_),
    .Y(_15140_));
 sky130_as_sc_hs__nor2_2 _46897_ (.A(_19528_),
    .B(_15128_),
    .Y(_15142_));
 sky130_as_sc_hs__or2_2 _46900_ (.A(\tholin_riscv.spi.counter[0] ),
    .B(\tholin_riscv.spi.counter[1] ),
    .Y(_15144_));
 sky130_as_sc_hs__nand3_2 _46903_ (.A(net501),
    .B(_15143_),
    .C(_15146_),
    .Y(_01049_));
 sky130_as_sc_hs__or2_2 _46906_ (.A(\tholin_riscv.spi.counter[2] ),
    .B(_15144_),
    .Y(_15149_));
 sky130_as_sc_hs__nand3_2 _46909_ (.A(net501),
    .B(_15147_),
    .C(_15151_),
    .Y(_01050_));
 sky130_as_sc_hs__and2_2 _46911_ (.A(\tholin_riscv.spi.counter[3] ),
    .B(_15149_),
    .Y(_15153_));
 sky130_as_sc_hs__nor2_2 _46912_ (.A(\tholin_riscv.spi.counter[3] ),
    .B(_15149_),
    .Y(_15154_));
 sky130_as_sc_hs__or2_2 _46913_ (.A(_15153_),
    .B(_15154_),
    .Y(_15155_));
 sky130_as_sc_hs__nand3_2 _46915_ (.A(net516),
    .B(_15152_),
    .C(_15156_),
    .Y(_01051_));
 sky130_as_sc_hs__nor2b_2 _46917_ (.A(_14837_),
    .Y(_15158_),
    .B(_15154_));
 sky130_as_sc_hs__or2_2 _46919_ (.A(net718),
    .B(_15158_),
    .Y(_15160_));
 sky130_as_sc_hs__and2_2 _46920_ (.A(net516),
    .B(_15159_),
    .Y(_15161_));
 sky130_as_sc_hs__nand3_2 _46921_ (.A(_15157_),
    .B(net719),
    .C(_15161_),
    .Y(_01052_));
 sky130_as_sc_hs__or2_2 _46922_ (.A(net1319),
    .B(_14840_),
    .Y(_15162_));
 sky130_as_sc_hs__or2_2 _46923_ (.A(\tholin_riscv.instr[0] ),
    .B(_14841_),
    .Y(_15163_));
 sky130_as_sc_hs__and2_2 _46924_ (.A(_15142_),
    .B(net1320),
    .Y(_15164_));
 sky130_as_sc_hs__and2_2 _46925_ (.A(_15163_),
    .B(net1321),
    .Y(_01053_));
 sky130_as_sc_hs__or2_2 _46926_ (.A(\tholin_riscv.spi.data_out_buff[1] ),
    .B(_14840_),
    .Y(_15165_));
 sky130_as_sc_hs__or2_2 _46927_ (.A(\tholin_riscv.instr[1] ),
    .B(_14841_),
    .Y(_15166_));
 sky130_as_sc_hs__nand3_2 _46928_ (.A(_15129_),
    .B(_15165_),
    .C(_15166_),
    .Y(_15167_));
 sky130_as_sc_hs__and2_2 _46931_ (.A(net515),
    .B(_15169_),
    .Y(_01054_));
 sky130_as_sc_hs__or2_2 _46932_ (.A(\tholin_riscv.spi.data_out_buff[2] ),
    .B(_14840_),
    .Y(_15170_));
 sky130_as_sc_hs__nand3_2 _46934_ (.A(_15129_),
    .B(_15170_),
    .C(_15171_),
    .Y(_15172_));
 sky130_as_sc_hs__and2_2 _46937_ (.A(net500),
    .B(_15174_),
    .Y(_01055_));
 sky130_as_sc_hs__or2_2 _46938_ (.A(\tholin_riscv.spi.data_out_buff[3] ),
    .B(_14840_),
    .Y(_15175_));
 sky130_as_sc_hs__nand3_2 _46940_ (.A(_15129_),
    .B(_15175_),
    .C(_15176_),
    .Y(_15177_));
 sky130_as_sc_hs__and2_2 _46943_ (.A(net500),
    .B(_15179_),
    .Y(_01056_));
 sky130_as_sc_hs__or2_2 _46944_ (.A(\tholin_riscv.spi.data_out_buff[4] ),
    .B(_14840_),
    .Y(_15180_));
 sky130_as_sc_hs__nand3_2 _46946_ (.A(_15129_),
    .B(_15180_),
    .C(_15181_),
    .Y(_15182_));
 sky130_as_sc_hs__and2_2 _46949_ (.A(net515),
    .B(_15184_),
    .Y(_01057_));
 sky130_as_sc_hs__or2_2 _46950_ (.A(\tholin_riscv.spi.data_out_buff[5] ),
    .B(_14840_),
    .Y(_15185_));
 sky130_as_sc_hs__nand3_2 _46952_ (.A(_15129_),
    .B(_15185_),
    .C(_15186_),
    .Y(_15187_));
 sky130_as_sc_hs__and2_2 _46955_ (.A(net501),
    .B(_15189_),
    .Y(_01058_));
 sky130_as_sc_hs__or2_2 _46956_ (.A(\tholin_riscv.spi.data_out_buff[6] ),
    .B(_14840_),
    .Y(_15190_));
 sky130_as_sc_hs__nand3_2 _46958_ (.A(_15129_),
    .B(_15190_),
    .C(_15191_),
    .Y(_15192_));
 sky130_as_sc_hs__and2_2 _46961_ (.A(net501),
    .B(_15194_),
    .Y(_01059_));
 sky130_as_sc_hs__or2_2 _46962_ (.A(\tholin_riscv.spi.data_out_buff[7] ),
    .B(_14840_),
    .Y(_15195_));
 sky130_as_sc_hs__or2_2 _46963_ (.A(\tholin_riscv.Bimm[11] ),
    .B(_14841_),
    .Y(_15196_));
 sky130_as_sc_hs__nand3_2 _46964_ (.A(_15129_),
    .B(_15195_),
    .C(_15196_),
    .Y(_15197_));
 sky130_as_sc_hs__and2_2 _46967_ (.A(net515),
    .B(_15199_),
    .Y(_01060_));
 sky130_as_sc_hs__and2_2 _46968_ (.A(_19901_),
    .B(_20733_),
    .Y(_15200_));
 sky130_as_sc_hs__nand3_2 _46972_ (.A(net518),
    .B(_15202_),
    .C(_15203_),
    .Y(_01061_));
 sky130_as_sc_hs__or2_2 _46974_ (.A(net1685),
    .B(_15201_),
    .Y(_15205_));
 sky130_as_sc_hs__and2_2 _46975_ (.A(net517),
    .B(_15204_),
    .Y(_15206_));
 sky130_as_sc_hs__and2_2 _46976_ (.A(_15205_),
    .B(_15206_),
    .Y(_01062_));
 sky130_as_sc_hs__and2_2 _46979_ (.A(net522),
    .B(_15207_),
    .Y(_15209_));
 sky130_as_sc_hs__and2_2 _46980_ (.A(_15208_),
    .B(_15209_),
    .Y(_01063_));
 sky130_as_sc_hs__and2_2 _46983_ (.A(net522),
    .B(_15210_),
    .Y(_15212_));
 sky130_as_sc_hs__and2_2 _46984_ (.A(_15211_),
    .B(_15212_),
    .Y(_01064_));
 sky130_as_sc_hs__and2_2 _46987_ (.A(net522),
    .B(_15213_),
    .Y(_15215_));
 sky130_as_sc_hs__and2_2 _46988_ (.A(_15214_),
    .B(_15215_),
    .Y(_01065_));
 sky130_as_sc_hs__and2_2 _46991_ (.A(net520),
    .B(_15216_),
    .Y(_15218_));
 sky130_as_sc_hs__and2_2 _46992_ (.A(_15217_),
    .B(_15218_),
    .Y(_01066_));
 sky130_as_sc_hs__and2_2 _46995_ (.A(net521),
    .B(_15219_),
    .Y(_15221_));
 sky130_as_sc_hs__and2_2 _46996_ (.A(_15220_),
    .B(_15221_),
    .Y(_01067_));
 sky130_as_sc_hs__or2_2 _46998_ (.A(net1688),
    .B(_15201_),
    .Y(_15223_));
 sky130_as_sc_hs__and2_2 _46999_ (.A(net517),
    .B(_15222_),
    .Y(_15224_));
 sky130_as_sc_hs__and2_2 _47000_ (.A(_15223_),
    .B(_15224_),
    .Y(_01068_));
 sky130_as_sc_hs__nand3_2 _47003_ (.A(net519),
    .B(_15225_),
    .C(_15226_),
    .Y(_01069_));
 sky130_as_sc_hs__or2_2 _47005_ (.A(net1168),
    .B(_15201_),
    .Y(_15228_));
 sky130_as_sc_hs__and2_2 _47006_ (.A(net517),
    .B(_15227_),
    .Y(_15229_));
 sky130_as_sc_hs__and2_2 _47007_ (.A(net1169),
    .B(_15229_),
    .Y(_01070_));
 sky130_as_sc_hs__or2_2 _47009_ (.A(net1374),
    .B(_15201_),
    .Y(_15231_));
 sky130_as_sc_hs__and2_2 _47010_ (.A(net520),
    .B(_15230_),
    .Y(_15232_));
 sky130_as_sc_hs__and2_2 _47011_ (.A(net1375),
    .B(_15232_),
    .Y(_01071_));
 sky130_as_sc_hs__or2_2 _47012_ (.A(net1830),
    .B(_15200_),
    .Y(_15233_));
 sky130_as_sc_hs__or2_2 _47013_ (.A(net1343),
    .B(_15201_),
    .Y(_15234_));
 sky130_as_sc_hs__and2_2 _47014_ (.A(net516),
    .B(_15233_),
    .Y(_15235_));
 sky130_as_sc_hs__and2_2 _47015_ (.A(net1344),
    .B(_15235_),
    .Y(_01072_));
 sky130_as_sc_hs__and2_2 _47018_ (.A(net520),
    .B(_15236_),
    .Y(_15238_));
 sky130_as_sc_hs__and2_2 _47019_ (.A(_15237_),
    .B(_15238_),
    .Y(_01073_));
 sky130_as_sc_hs__and2_2 _47022_ (.A(net520),
    .B(_15239_),
    .Y(_15241_));
 sky130_as_sc_hs__and2_2 _47023_ (.A(_15240_),
    .B(_15241_),
    .Y(_01074_));
 sky130_as_sc_hs__or2_2 _47025_ (.A(net1032),
    .B(_15201_),
    .Y(_15243_));
 sky130_as_sc_hs__and2_2 _47026_ (.A(net516),
    .B(_15242_),
    .Y(_15244_));
 sky130_as_sc_hs__and2_2 _47027_ (.A(net1033),
    .B(_15244_),
    .Y(_01075_));
 sky130_as_sc_hs__and2_2 _47030_ (.A(net517),
    .B(_15245_),
    .Y(_15247_));
 sky130_as_sc_hs__and2_2 _47031_ (.A(_15246_),
    .B(_15247_),
    .Y(_01076_));
 sky130_as_sc_hs__nor2_2 _47033_ (.A(_19899_),
    .B(_15248_),
    .Y(_15249_));
 sky130_as_sc_hs__or2_2 _47034_ (.A(net627),
    .B(_15249_),
    .Y(_15250_));
 sky130_as_sc_hs__and2_2 _47036_ (.A(net515),
    .B(_15251_),
    .Y(_15252_));
 sky130_as_sc_hs__and2_2 _47037_ (.A(net628),
    .B(_15252_),
    .Y(_01077_));
 sky130_as_sc_hs__or2_2 _47038_ (.A(net611),
    .B(_15249_),
    .Y(_15253_));
 sky130_as_sc_hs__and2_2 _47040_ (.A(net515),
    .B(_15254_),
    .Y(_15255_));
 sky130_as_sc_hs__and2_2 _47041_ (.A(net612),
    .B(_15255_),
    .Y(_01078_));
 sky130_as_sc_hs__or2_2 _47042_ (.A(net618),
    .B(_15249_),
    .Y(_15256_));
 sky130_as_sc_hs__and2_2 _47044_ (.A(net511),
    .B(_15257_),
    .Y(_15258_));
 sky130_as_sc_hs__and2_2 _47045_ (.A(net619),
    .B(_15258_),
    .Y(_01079_));
 sky130_as_sc_hs__or2_2 _47046_ (.A(net772),
    .B(_15249_),
    .Y(_15259_));
 sky130_as_sc_hs__and2_2 _47048_ (.A(net511),
    .B(_15260_),
    .Y(_15261_));
 sky130_as_sc_hs__and2_2 _47049_ (.A(net773),
    .B(_15261_),
    .Y(_01080_));
 sky130_as_sc_hs__or2_2 _47050_ (.A(net648),
    .B(_15249_),
    .Y(_15262_));
 sky130_as_sc_hs__and2_2 _47052_ (.A(net511),
    .B(_15263_),
    .Y(_15264_));
 sky130_as_sc_hs__and2_2 _47053_ (.A(net649),
    .B(_15264_),
    .Y(_01081_));
 sky130_as_sc_hs__or2_2 _47054_ (.A(net624),
    .B(_15249_),
    .Y(_15265_));
 sky130_as_sc_hs__and2_2 _47056_ (.A(net515),
    .B(_15266_),
    .Y(_15267_));
 sky130_as_sc_hs__and2_2 _47057_ (.A(net625),
    .B(_15267_),
    .Y(_01082_));
 sky130_as_sc_hs__or2_2 _47058_ (.A(net751),
    .B(_15249_),
    .Y(_15268_));
 sky130_as_sc_hs__and2_2 _47060_ (.A(net511),
    .B(_15269_),
    .Y(_15270_));
 sky130_as_sc_hs__and2_2 _47061_ (.A(net752),
    .B(_15270_),
    .Y(_01083_));
 sky130_as_sc_hs__or2_2 _47062_ (.A(\tholin_riscv.spi.divisor[7] ),
    .B(_15249_),
    .Y(_15271_));
 sky130_as_sc_hs__nand3_2 _47063_ (.A(_21468_),
    .B(_21469_),
    .C(_15249_),
    .Y(_15272_));
 sky130_as_sc_hs__nor2_2 _47066_ (.A(_19935_),
    .B(_19972_),
    .Y(_15274_));
 sky130_as_sc_hs__and2_2 _47067_ (.A(net501),
    .B(_15274_),
    .Y(_15275_));
 sky130_as_sc_hs__or2_2 _47069_ (.A(\tholin_riscv.Bimm[11] ),
    .B(_15276_),
    .Y(_15277_));
 sky130_as_sc_hs__or2_2 _47070_ (.A(net645),
    .B(_15275_),
    .Y(_15278_));
 sky130_as_sc_hs__and2_2 _47071_ (.A(_15277_),
    .B(net646),
    .Y(_01085_));
 sky130_as_sc_hs__or2_2 _47072_ (.A(net1710),
    .B(_15276_),
    .Y(_15279_));
 sky130_as_sc_hs__or2_2 _47073_ (.A(net630),
    .B(_15275_),
    .Y(_15280_));
 sky130_as_sc_hs__and2_2 _47074_ (.A(_15279_),
    .B(net631),
    .Y(_01086_));
 sky130_as_sc_hs__or2_2 _47075_ (.A(net1168),
    .B(_15276_),
    .Y(_15281_));
 sky130_as_sc_hs__or2_2 _47076_ (.A(net642),
    .B(_15275_),
    .Y(_15282_));
 sky130_as_sc_hs__and2_2 _47077_ (.A(_15281_),
    .B(net643),
    .Y(_01087_));
 sky130_as_sc_hs__or2_2 _47078_ (.A(net1374),
    .B(_15276_),
    .Y(_15283_));
 sky130_as_sc_hs__or2_2 _47079_ (.A(net636),
    .B(_15275_),
    .Y(_15284_));
 sky130_as_sc_hs__and2_2 _47080_ (.A(_15283_),
    .B(net637),
    .Y(_01088_));
 sky130_as_sc_hs__or2_2 _47081_ (.A(net1794),
    .B(_15276_),
    .Y(_15285_));
 sky130_as_sc_hs__or2_2 _47082_ (.A(net633),
    .B(_15275_),
    .Y(_15286_));
 sky130_as_sc_hs__and2_2 _47083_ (.A(_15285_),
    .B(net634),
    .Y(_01089_));
 sky130_as_sc_hs__and2_2 _47084_ (.A(_19749_),
    .B(_21561_),
    .Y(_15287_));
 sky130_as_sc_hs__or2_2 _47085_ (.A(net145),
    .B(net134),
    .Y(_15288_));
 sky130_as_sc_hs__or2_2 _47086_ (.A(_19935_),
    .B(_06165_),
    .Y(_15289_));
 sky130_as_sc_hs__and2_2 _47087_ (.A(_15288_),
    .B(_15289_),
    .Y(_15290_));
 sky130_as_sc_hs__nand3_2 _47089_ (.A(\tholin_riscv.cycle[3] ),
    .B(_19501_),
    .C(net134),
    .Y(_15292_));
 sky130_as_sc_hs__and2_2 _47092_ (.A(net494),
    .B(_15294_),
    .Y(_01090_));
 sky130_as_sc_hs__nor2_2 _47094_ (.A(\tholin_riscv.div_counter[1] ),
    .B(\tholin_riscv.div_counter[0] ),
    .Y(_15296_));
 sky130_as_sc_hs__and2_2 _47095_ (.A(\tholin_riscv.div_counter[1] ),
    .B(\tholin_riscv.div_counter[0] ),
    .Y(_15297_));
 sky130_as_sc_hs__nor2_2 _47096_ (.A(_15296_),
    .B(_15297_),
    .Y(_15298_));
 sky130_as_sc_hs__and2_2 _47099_ (.A(net494),
    .B(_15300_),
    .Y(_01091_));
 sky130_as_sc_hs__and2_2 _47101_ (.A(\tholin_riscv.div_counter[2] ),
    .B(_15297_),
    .Y(_15302_));
 sky130_as_sc_hs__or2_2 _47102_ (.A(\tholin_riscv.div_counter[2] ),
    .B(_15297_),
    .Y(_15303_));
 sky130_as_sc_hs__or2_2 _47104_ (.A(_15302_),
    .B(_15304_),
    .Y(_15305_));
 sky130_as_sc_hs__and2_2 _47106_ (.A(net494),
    .B(_15306_),
    .Y(_01092_));
 sky130_as_sc_hs__or2_2 _47108_ (.A(\tholin_riscv.div_counter[3] ),
    .B(_15302_),
    .Y(_15308_));
 sky130_as_sc_hs__and2_2 _47109_ (.A(\tholin_riscv.div_counter[3] ),
    .B(_15302_),
    .Y(_15309_));
 sky130_as_sc_hs__or2_2 _47111_ (.A(_15309_),
    .B(_15310_),
    .Y(_15311_));
 sky130_as_sc_hs__and2_2 _47113_ (.A(net494),
    .B(_15312_),
    .Y(_01093_));
 sky130_as_sc_hs__and2_2 _47115_ (.A(\tholin_riscv.div_counter[4] ),
    .B(_15309_),
    .Y(_15314_));
 sky130_as_sc_hs__or2_2 _47116_ (.A(\tholin_riscv.div_counter[4] ),
    .B(_15309_),
    .Y(_15315_));
 sky130_as_sc_hs__or2_2 _47118_ (.A(_15314_),
    .B(_15316_),
    .Y(_15317_));
 sky130_as_sc_hs__and2_2 _47120_ (.A(net494),
    .B(_15318_),
    .Y(_01094_));
 sky130_as_sc_hs__or2_2 _47123_ (.A(_02381_),
    .B(_06546_),
    .Y(_15321_));
 sky130_as_sc_hs__or2_2 _47125_ (.A(\tholin_riscv.div_shifter[61] ),
    .B(_15322_),
    .Y(_15323_));
 sky130_as_sc_hs__and2_2 _47127_ (.A(_15323_),
    .B(_15324_),
    .Y(_15325_));
 sky130_as_sc_hs__or2_2 _47130_ (.A(\tholin_riscv.div_shifter[62] ),
    .B(_15327_),
    .Y(_15328_));
 sky130_as_sc_hs__or2_2 _47137_ (.A(\tholin_riscv.div_shifter[58] ),
    .B(_15333_),
    .Y(_15335_));
 sky130_as_sc_hs__or2_2 _47142_ (.A(\tholin_riscv.div_shifter[55] ),
    .B(_15339_),
    .Y(_15340_));
 sky130_as_sc_hs__and2_2 _47144_ (.A(_15340_),
    .B(_15341_),
    .Y(_15342_));
 sky130_as_sc_hs__or2_2 _47149_ (.A(\tholin_riscv.div_shifter[56] ),
    .B(_15345_),
    .Y(_15347_));
 sky130_as_sc_hs__and2_2 _47150_ (.A(_15346_),
    .B(_15347_),
    .Y(_15348_));
 sky130_as_sc_hs__inv_2 _47151_ (.Y(_15349_),
    .A(_15348_));
 sky130_as_sc_hs__or2_2 _47156_ (.A(\tholin_riscv.div_shifter[57] ),
    .B(_15352_),
    .Y(_15354_));
 sky130_as_sc_hs__and2_2 _47157_ (.A(_15353_),
    .B(_15354_),
    .Y(_15355_));
 sky130_as_sc_hs__nand3_2 _47158_ (.A(_15342_),
    .B(_15348_),
    .C(_15355_),
    .Y(_15356_));
 sky130_as_sc_hs__or2_2 _47159_ (.A(_15336_),
    .B(_15356_),
    .Y(_15357_));
 sky130_as_sc_hs__nor2_2 _47160_ (.A(_15330_),
    .B(_15357_),
    .Y(_15358_));
 sky130_as_sc_hs__or2_2 _47164_ (.A(\tholin_riscv.div_shifter[59] ),
    .B(_15361_),
    .Y(_15362_));
 sky130_as_sc_hs__and2_2 _47166_ (.A(_15362_),
    .B(_15363_),
    .Y(_15364_));
 sky130_as_sc_hs__or2_2 _47170_ (.A(\tholin_riscv.div_shifter[60] ),
    .B(_15367_),
    .Y(_15368_));
 sky130_as_sc_hs__and2_2 _47172_ (.A(_15368_),
    .B(_15369_),
    .Y(_15370_));
 sky130_as_sc_hs__and2_2 _47173_ (.A(_15364_),
    .B(_15370_),
    .Y(_15371_));
 sky130_as_sc_hs__and2_2 _47174_ (.A(_15325_),
    .B(_15371_),
    .Y(_15372_));
 sky130_as_sc_hs__and2_2 _47175_ (.A(_15358_),
    .B(_15372_),
    .Y(_15373_));
 sky130_as_sc_hs__or2_2 _47180_ (.A(\tholin_riscv.div_shifter[44] ),
    .B(_15376_),
    .Y(_15378_));
 sky130_as_sc_hs__and2_2 _47181_ (.A(_15377_),
    .B(_15378_),
    .Y(_15379_));
 sky130_as_sc_hs__or2_2 _47185_ (.A(\tholin_riscv.div_shifter[43] ),
    .B(_15382_),
    .Y(_15383_));
 sky130_as_sc_hs__and2_2 _47187_ (.A(_15383_),
    .B(_15384_),
    .Y(_15385_));
 sky130_as_sc_hs__or2_2 _47191_ (.A(\tholin_riscv.div_shifter[42] ),
    .B(_15388_),
    .Y(_15389_));
 sky130_as_sc_hs__and2_2 _47193_ (.A(_15389_),
    .B(_15390_),
    .Y(_15391_));
 sky130_as_sc_hs__or2_2 _47197_ (.A(\tholin_riscv.div_shifter[41] ),
    .B(_15394_),
    .Y(_15395_));
 sky130_as_sc_hs__and2_2 _47199_ (.A(_15395_),
    .B(_15396_),
    .Y(_15397_));
 sky130_as_sc_hs__and2_2 _47202_ (.A(_15398_),
    .B(_15399_),
    .Y(_15400_));
 sky130_as_sc_hs__or2_2 _47203_ (.A(\tholin_riscv.div_shifter[40] ),
    .B(_15400_),
    .Y(_15401_));
 sky130_as_sc_hs__and2_2 _47205_ (.A(_15401_),
    .B(_15402_),
    .Y(_15403_));
 sky130_as_sc_hs__and2_2 _47208_ (.A(_15404_),
    .B(_15405_),
    .Y(_15406_));
 sky130_as_sc_hs__or2_2 _47209_ (.A(\tholin_riscv.div_shifter[39] ),
    .B(_15406_),
    .Y(_15407_));
 sky130_as_sc_hs__and2_2 _47211_ (.A(_15407_),
    .B(_15408_),
    .Y(_15409_));
 sky130_as_sc_hs__nand3_2 _47212_ (.A(_15385_),
    .B(_15403_),
    .C(_15409_),
    .Y(_15410_));
 sky130_as_sc_hs__nor2_2 _47214_ (.A(_15410_),
    .B(_15411_),
    .Y(_15412_));
 sky130_as_sc_hs__and2_2 _47215_ (.A(_15391_),
    .B(_15412_),
    .Y(_15413_));
 sky130_as_sc_hs__and2_2 _47218_ (.A(_15414_),
    .B(_15415_),
    .Y(_15416_));
 sky130_as_sc_hs__and2_2 _47222_ (.A(_15418_),
    .B(_15419_),
    .Y(_15420_));
 sky130_as_sc_hs__or2_2 _47223_ (.A(\tholin_riscv.div_shifter[34] ),
    .B(_15420_),
    .Y(_15421_));
 sky130_as_sc_hs__and2_2 _47226_ (.A(_15422_),
    .B(_15423_),
    .Y(_15424_));
 sky130_as_sc_hs__or2_2 _47231_ (.A(_19499_),
    .B(_15428_),
    .Y(_15429_));
 sky130_as_sc_hs__and2_2 _47232_ (.A(_19500_),
    .B(net116),
    .Y(_15430_));
 sky130_as_sc_hs__or2_2 _47235_ (.A(_15430_),
    .B(_15432_),
    .Y(_15433_));
 sky130_as_sc_hs__or2_2 _47237_ (.A(\tholin_riscv.div_shifter[33] ),
    .B(_15424_),
    .Y(_15435_));
 sky130_as_sc_hs__and2_2 _47238_ (.A(_15425_),
    .B(_15435_),
    .Y(_15436_));
 sky130_as_sc_hs__and2_2 _47242_ (.A(\tholin_riscv.div_shifter[31] ),
    .B(_20826_),
    .Y(_15440_));
 sky130_as_sc_hs__nor2_2 _47243_ (.A(_15433_),
    .B(_15440_),
    .Y(_15441_));
 sky130_as_sc_hs__and2_2 _47244_ (.A(_15425_),
    .B(_15441_),
    .Y(_15442_));
 sky130_as_sc_hs__or2_2 _47245_ (.A(_15439_),
    .B(_15442_),
    .Y(_15443_));
 sky130_as_sc_hs__or2_2 _47246_ (.A(_21242_),
    .B(_06546_),
    .Y(_15444_));
 sky130_as_sc_hs__and2_2 _47248_ (.A(_15444_),
    .B(_15445_),
    .Y(_15446_));
 sky130_as_sc_hs__nand3_2 _47251_ (.A(_15443_),
    .B(_15447_),
    .C(_15448_),
    .Y(_15449_));
 sky130_as_sc_hs__or2_2 _47252_ (.A(\tholin_riscv.div_shifter[35] ),
    .B(_15446_),
    .Y(_15450_));
 sky130_as_sc_hs__and2_2 _47255_ (.A(_15451_),
    .B(_15452_),
    .Y(_15453_));
 sky130_as_sc_hs__or2_2 _47256_ (.A(\tholin_riscv.div_shifter[36] ),
    .B(_15453_),
    .Y(_15454_));
 sky130_as_sc_hs__nand3_2 _47257_ (.A(_15449_),
    .B(_15450_),
    .C(_15454_),
    .Y(_15455_));
 sky130_as_sc_hs__and2_2 _47261_ (.A(_15457_),
    .B(_15458_),
    .Y(_15459_));
 sky130_as_sc_hs__nand3_2 _47263_ (.A(_15455_),
    .B(_15456_),
    .C(_15460_),
    .Y(_15461_));
 sky130_as_sc_hs__or2_2 _47264_ (.A(\tholin_riscv.div_shifter[38] ),
    .B(_15416_),
    .Y(_15462_));
 sky130_as_sc_hs__or2_2 _47265_ (.A(\tholin_riscv.div_shifter[37] ),
    .B(_15459_),
    .Y(_15463_));
 sky130_as_sc_hs__nand3_2 _47266_ (.A(_15461_),
    .B(_15462_),
    .C(_15463_),
    .Y(_15464_));
 sky130_as_sc_hs__nand3_2 _47267_ (.A(_15413_),
    .B(_15417_),
    .C(_15464_),
    .Y(_15465_));
 sky130_as_sc_hs__nand2b_2 _47268_ (.B(_15402_),
    .Y(_15466_),
    .A(_15407_));
 sky130_as_sc_hs__nand3_2 _47269_ (.A(_15395_),
    .B(_15401_),
    .C(_15466_),
    .Y(_15467_));
 sky130_as_sc_hs__nand3_2 _47270_ (.A(_15390_),
    .B(_15396_),
    .C(_15467_),
    .Y(_15468_));
 sky130_as_sc_hs__nand3_2 _47271_ (.A(_15383_),
    .B(_15389_),
    .C(_15468_),
    .Y(_15469_));
 sky130_as_sc_hs__nand3_2 _47272_ (.A(_15377_),
    .B(_15384_),
    .C(_15469_),
    .Y(_15470_));
 sky130_as_sc_hs__nand3_2 _47273_ (.A(_15378_),
    .B(_15465_),
    .C(_15470_),
    .Y(_15471_));
 sky130_as_sc_hs__or2_2 _47275_ (.A(_20622_),
    .B(_06546_),
    .Y(_15473_));
 sky130_as_sc_hs__or2_2 _47280_ (.A(_20707_),
    .B(_06546_),
    .Y(_15478_));
 sky130_as_sc_hs__or2_2 _47282_ (.A(\tholin_riscv.div_shifter[46] ),
    .B(_15479_),
    .Y(_15480_));
 sky130_as_sc_hs__or2_2 _47283_ (.A(\tholin_riscv.div_shifter[45] ),
    .B(_15474_),
    .Y(_15481_));
 sky130_as_sc_hs__nand3_2 _47284_ (.A(_15476_),
    .B(_15480_),
    .C(_15481_),
    .Y(_15482_));
 sky130_as_sc_hs__or2_2 _47289_ (.A(\tholin_riscv.div_shifter[54] ),
    .B(_15485_),
    .Y(_15487_));
 sky130_as_sc_hs__and2_2 _47290_ (.A(_15486_),
    .B(_15487_),
    .Y(_15488_));
 sky130_as_sc_hs__inv_2 _47291_ (.Y(_15489_),
    .A(_15488_));
 sky130_as_sc_hs__or2_2 _47295_ (.A(\tholin_riscv.div_shifter[53] ),
    .B(_15492_),
    .Y(_15493_));
 sky130_as_sc_hs__or2_2 _47302_ (.A(\tholin_riscv.div_shifter[52] ),
    .B(_15498_),
    .Y(_15500_));
 sky130_as_sc_hs__and2_2 _47303_ (.A(_15499_),
    .B(_15500_),
    .Y(_15501_));
 sky130_as_sc_hs__or2_2 _47307_ (.A(\tholin_riscv.div_shifter[51] ),
    .B(_15504_),
    .Y(_15505_));
 sky130_as_sc_hs__and2_2 _47309_ (.A(_15505_),
    .B(_15506_),
    .Y(_15507_));
 sky130_as_sc_hs__or2_2 _47314_ (.A(\tholin_riscv.div_shifter[50] ),
    .B(_15510_),
    .Y(_15512_));
 sky130_as_sc_hs__and2_2 _47315_ (.A(_15511_),
    .B(_15512_),
    .Y(_15513_));
 sky130_as_sc_hs__or2_2 _47319_ (.A(\tholin_riscv.div_shifter[49] ),
    .B(_15516_),
    .Y(_15517_));
 sky130_as_sc_hs__and2_2 _47321_ (.A(_15517_),
    .B(_15518_),
    .Y(_15519_));
 sky130_as_sc_hs__or2_2 _47325_ (.A(\tholin_riscv.div_shifter[48] ),
    .B(_15522_),
    .Y(_15523_));
 sky130_as_sc_hs__and2_2 _47327_ (.A(_15523_),
    .B(_15524_),
    .Y(_15525_));
 sky130_as_sc_hs__inv_2 _47328_ (.Y(_15526_),
    .A(_15525_));
 sky130_as_sc_hs__or2_2 _47329_ (.A(_24037_),
    .B(_06546_),
    .Y(_15527_));
 sky130_as_sc_hs__and2_2 _47331_ (.A(_15527_),
    .B(_15528_),
    .Y(_15529_));
 sky130_as_sc_hs__or2_2 _47332_ (.A(\tholin_riscv.div_shifter[47] ),
    .B(_15529_),
    .Y(_15530_));
 sky130_as_sc_hs__inv_2 _47333_ (.Y(_15531_),
    .A(_15530_));
 sky130_as_sc_hs__and2_2 _47335_ (.A(_15530_),
    .B(_15532_),
    .Y(_15533_));
 sky130_as_sc_hs__and2_2 _47336_ (.A(_15525_),
    .B(_15533_),
    .Y(_15534_));
 sky130_as_sc_hs__and2_2 _47337_ (.A(_15519_),
    .B(_15534_),
    .Y(_15535_));
 sky130_as_sc_hs__and2_2 _47338_ (.A(_15513_),
    .B(_15535_),
    .Y(_15536_));
 sky130_as_sc_hs__nand3_2 _47339_ (.A(_15501_),
    .B(_15507_),
    .C(_15536_),
    .Y(_15537_));
 sky130_as_sc_hs__nor2_2 _47340_ (.A(_15495_),
    .B(_15537_),
    .Y(_15538_));
 sky130_as_sc_hs__and2_2 _47341_ (.A(_15488_),
    .B(_15538_),
    .Y(_15539_));
 sky130_as_sc_hs__and2_2 _47344_ (.A(_15475_),
    .B(_15481_),
    .Y(_15542_));
 sky130_as_sc_hs__nand3_2 _47345_ (.A(_15482_),
    .B(_15539_),
    .C(_15540_),
    .Y(_15543_));
 sky130_as_sc_hs__nand3_2 _47347_ (.A(_15517_),
    .B(_15523_),
    .C(_15544_),
    .Y(_15545_));
 sky130_as_sc_hs__nand3_2 _47348_ (.A(_15511_),
    .B(_15518_),
    .C(_15545_),
    .Y(_15546_));
 sky130_as_sc_hs__nand3_2 _47349_ (.A(_15505_),
    .B(_15512_),
    .C(_15546_),
    .Y(_15547_));
 sky130_as_sc_hs__nand3_2 _47350_ (.A(_15499_),
    .B(_15506_),
    .C(_15547_),
    .Y(_15548_));
 sky130_as_sc_hs__nand3_2 _47351_ (.A(_15493_),
    .B(_15500_),
    .C(_15548_),
    .Y(_15549_));
 sky130_as_sc_hs__nand3_2 _47352_ (.A(_15486_),
    .B(_15494_),
    .C(_15549_),
    .Y(_15550_));
 sky130_as_sc_hs__nand3_2 _47353_ (.A(_15487_),
    .B(_15543_),
    .C(_15550_),
    .Y(_15551_));
 sky130_as_sc_hs__nand3_2 _47356_ (.A(_15346_),
    .B(_15353_),
    .C(_15553_),
    .Y(_15554_));
 sky130_as_sc_hs__nand3_2 _47357_ (.A(_15335_),
    .B(_15354_),
    .C(_15554_),
    .Y(_15555_));
 sky130_as_sc_hs__nand3_2 _47358_ (.A(_15334_),
    .B(_15371_),
    .C(_15555_),
    .Y(_15556_));
 sky130_as_sc_hs__nand2b_2 _47359_ (.B(_15369_),
    .Y(_15557_),
    .A(_15362_));
 sky130_as_sc_hs__and2_2 _47360_ (.A(_15368_),
    .B(_15557_),
    .Y(_15558_));
 sky130_as_sc_hs__nand3_2 _47361_ (.A(_15323_),
    .B(_15556_),
    .C(_15558_),
    .Y(_15559_));
 sky130_as_sc_hs__nand3_2 _47362_ (.A(_15324_),
    .B(_15329_),
    .C(_15559_),
    .Y(_15560_));
 sky130_as_sc_hs__nand3_2 _47363_ (.A(_15328_),
    .B(_15552_),
    .C(_15560_),
    .Y(_15561_));
 sky130_as_sc_hs__and2_2 _47365_ (.A(_15460_),
    .B(_15463_),
    .Y(_15563_));
 sky130_as_sc_hs__and2_2 _47366_ (.A(_15454_),
    .B(_15456_),
    .Y(_15564_));
 sky130_as_sc_hs__and2_2 _47368_ (.A(_15421_),
    .B(_15448_),
    .Y(_15566_));
 sky130_as_sc_hs__nand3_2 _47369_ (.A(_15436_),
    .B(_15441_),
    .C(_15566_),
    .Y(_15567_));
 sky130_as_sc_hs__nor2_2 _47370_ (.A(_15565_),
    .B(_15567_),
    .Y(_15568_));
 sky130_as_sc_hs__nand3_2 _47371_ (.A(_15563_),
    .B(_15564_),
    .C(_15568_),
    .Y(_15569_));
 sky130_as_sc_hs__nor2_2 _47372_ (.A(_15562_),
    .B(_15569_),
    .Y(_15570_));
 sky130_as_sc_hs__nand3_2 _47373_ (.A(_15413_),
    .B(_15542_),
    .C(_15570_),
    .Y(_15571_));
 sky130_as_sc_hs__nor2_2 _47374_ (.A(_15541_),
    .B(_15571_),
    .Y(_15572_));
 sky130_as_sc_hs__nand3_2 _47375_ (.A(_15373_),
    .B(_15539_),
    .C(_15572_),
    .Y(_15573_));
 sky130_as_sc_hs__and2_2 _47379_ (.A(net497),
    .B(_15576_),
    .Y(_01095_));
 sky130_as_sc_hs__and2_2 _47383_ (.A(net497),
    .B(_15579_),
    .Y(_01096_));
 sky130_as_sc_hs__and2_2 _47387_ (.A(net487),
    .B(_15582_),
    .Y(_01097_));
 sky130_as_sc_hs__and2_2 _47391_ (.A(net487),
    .B(_15585_),
    .Y(_01098_));
 sky130_as_sc_hs__and2_2 _47395_ (.A(net487),
    .B(_15588_),
    .Y(_01099_));
 sky130_as_sc_hs__and2_2 _47399_ (.A(net487),
    .B(_15591_),
    .Y(_01100_));
 sky130_as_sc_hs__and2_2 _47403_ (.A(net487),
    .B(_15594_),
    .Y(_01101_));
 sky130_as_sc_hs__and2_2 _47407_ (.A(net487),
    .B(_15597_),
    .Y(_01102_));
 sky130_as_sc_hs__and2_2 _47411_ (.A(net487),
    .B(_15600_),
    .Y(_01103_));
 sky130_as_sc_hs__and2_2 _47415_ (.A(net487),
    .B(_15603_),
    .Y(_01104_));
 sky130_as_sc_hs__and2_2 _47419_ (.A(net487),
    .B(_15606_),
    .Y(_01105_));
 sky130_as_sc_hs__and2_2 _47423_ (.A(net496),
    .B(_15609_),
    .Y(_01106_));
 sky130_as_sc_hs__and2_2 _47427_ (.A(net496),
    .B(_15612_),
    .Y(_01107_));
 sky130_as_sc_hs__and2_2 _47431_ (.A(net496),
    .B(_15615_),
    .Y(_01108_));
 sky130_as_sc_hs__and2_2 _47435_ (.A(net486),
    .B(_15618_),
    .Y(_01109_));
 sky130_as_sc_hs__and2_2 _47439_ (.A(net486),
    .B(_15621_),
    .Y(_01110_));
 sky130_as_sc_hs__and2_2 _47443_ (.A(net486),
    .B(_15624_),
    .Y(_01111_));
 sky130_as_sc_hs__and2_2 _47447_ (.A(net486),
    .B(_15627_),
    .Y(_01112_));
 sky130_as_sc_hs__and2_2 _47451_ (.A(net486),
    .B(_15630_),
    .Y(_01113_));
 sky130_as_sc_hs__and2_2 _47455_ (.A(net487),
    .B(_15633_),
    .Y(_01114_));
 sky130_as_sc_hs__and2_2 _47459_ (.A(net487),
    .B(_15636_),
    .Y(_01115_));
 sky130_as_sc_hs__and2_2 _47463_ (.A(net487),
    .B(_15639_),
    .Y(_01116_));
 sky130_as_sc_hs__and2_2 _47467_ (.A(net487),
    .B(_15642_),
    .Y(_01117_));
 sky130_as_sc_hs__and2_2 _47471_ (.A(net484),
    .B(_15645_),
    .Y(_01118_));
 sky130_as_sc_hs__and2_2 _47475_ (.A(net484),
    .B(_15648_),
    .Y(_01119_));
 sky130_as_sc_hs__and2_2 _47479_ (.A(net484),
    .B(_15651_),
    .Y(_01120_));
 sky130_as_sc_hs__and2_2 _47483_ (.A(net484),
    .B(_15654_),
    .Y(_01121_));
 sky130_as_sc_hs__and2_2 _47487_ (.A(net484),
    .B(_15657_),
    .Y(_01122_));
 sky130_as_sc_hs__and2_2 _47491_ (.A(net484),
    .B(_15660_),
    .Y(_01123_));
 sky130_as_sc_hs__and2_2 _47495_ (.A(net484),
    .B(_15663_),
    .Y(_01124_));
 sky130_as_sc_hs__and2_2 _47499_ (.A(net496),
    .B(_15666_),
    .Y(_01125_));
 sky130_as_sc_hs__and2_2 _47503_ (.A(net496),
    .B(_15669_),
    .Y(_01126_));
 sky130_as_sc_hs__nand3_2 _47505_ (.A(net145),
    .B(net113),
    .C(_06165_),
    .Y(_15671_));
 sky130_as_sc_hs__and2_2 _47507_ (.A(net526),
    .B(_15672_),
    .Y(_01127_));
 sky130_as_sc_hs__nand3_2 _47510_ (.A(net143),
    .B(_15673_),
    .C(_15674_),
    .Y(_15675_));
 sky130_as_sc_hs__nand3_2 _47512_ (.A(net102),
    .B(_15675_),
    .C(_15676_),
    .Y(_15677_));
 sky130_as_sc_hs__or2_2 _47513_ (.A(net1214),
    .B(net102),
    .Y(_15678_));
 sky130_as_sc_hs__and2_2 _47514_ (.A(net498),
    .B(net1215),
    .Y(_15679_));
 sky130_as_sc_hs__and2_2 _47515_ (.A(_15677_),
    .B(net1216),
    .Y(_01128_));
 sky130_as_sc_hs__and2_2 _47516_ (.A(_22169_),
    .B(_06548_),
    .Y(_15680_));
 sky130_as_sc_hs__or2_2 _47518_ (.A(_22040_),
    .B(_15680_),
    .Y(_15682_));
 sky130_as_sc_hs__nand3_2 _47519_ (.A(net144),
    .B(_15681_),
    .C(_15682_),
    .Y(_15683_));
 sky130_as_sc_hs__nand3_2 _47521_ (.A(net100),
    .B(_15683_),
    .C(_15684_),
    .Y(_15685_));
 sky130_as_sc_hs__or2_2 _47522_ (.A(net1289),
    .B(net102),
    .Y(_15686_));
 sky130_as_sc_hs__and2_2 _47523_ (.A(net527),
    .B(net1290),
    .Y(_15687_));
 sky130_as_sc_hs__and2_2 _47524_ (.A(_15685_),
    .B(net1291),
    .Y(_01129_));
 sky130_as_sc_hs__or2_2 _47525_ (.A(_24051_),
    .B(_06549_),
    .Y(_15688_));
 sky130_as_sc_hs__or2_2 _47526_ (.A(_21977_),
    .B(_06548_),
    .Y(_15689_));
 sky130_as_sc_hs__nand3_2 _47527_ (.A(net143),
    .B(_15688_),
    .C(_15689_),
    .Y(_15690_));
 sky130_as_sc_hs__nand3_2 _47529_ (.A(net101),
    .B(_15690_),
    .C(_15691_),
    .Y(_15692_));
 sky130_as_sc_hs__or2_2 _47530_ (.A(net1274),
    .B(net101),
    .Y(_15693_));
 sky130_as_sc_hs__and2_2 _47531_ (.A(net498),
    .B(net1275),
    .Y(_15694_));
 sky130_as_sc_hs__and2_2 _47532_ (.A(_15692_),
    .B(net1276),
    .Y(_01130_));
 sky130_as_sc_hs__nand3_2 _47535_ (.A(net143),
    .B(_15695_),
    .C(_15696_),
    .Y(_15697_));
 sky130_as_sc_hs__nand3_2 _47537_ (.A(net102),
    .B(_15697_),
    .C(_15698_),
    .Y(_15699_));
 sky130_as_sc_hs__or2_2 _47538_ (.A(net1248),
    .B(net102),
    .Y(_15700_));
 sky130_as_sc_hs__and2_2 _47539_ (.A(net498),
    .B(net1249),
    .Y(_15701_));
 sky130_as_sc_hs__and2_2 _47540_ (.A(_15699_),
    .B(net1250),
    .Y(_01131_));
 sky130_as_sc_hs__or2_2 _47542_ (.A(_21914_),
    .B(_06548_),
    .Y(_15703_));
 sky130_as_sc_hs__nand3_2 _47543_ (.A(net144),
    .B(_15702_),
    .C(_15703_),
    .Y(_15704_));
 sky130_as_sc_hs__nand3_2 _47545_ (.A(net102),
    .B(_15704_),
    .C(_15705_),
    .Y(_15706_));
 sky130_as_sc_hs__or2_2 _47546_ (.A(net1340),
    .B(net102),
    .Y(_15707_));
 sky130_as_sc_hs__and2_2 _47547_ (.A(net527),
    .B(net1341),
    .Y(_15708_));
 sky130_as_sc_hs__and2_2 _47548_ (.A(_15706_),
    .B(net1342),
    .Y(_01132_));
 sky130_as_sc_hs__nand3_2 _47551_ (.A(net143),
    .B(_15709_),
    .C(_15710_),
    .Y(_15711_));
 sky130_as_sc_hs__nand3_2 _47553_ (.A(net99),
    .B(_15711_),
    .C(_15712_),
    .Y(_15713_));
 sky130_as_sc_hs__or2_2 _47554_ (.A(net1103),
    .B(net99),
    .Y(_15714_));
 sky130_as_sc_hs__and2_2 _47555_ (.A(net498),
    .B(net1104),
    .Y(_15715_));
 sky130_as_sc_hs__and2_2 _47556_ (.A(_15713_),
    .B(net1105),
    .Y(_01133_));
 sky130_as_sc_hs__nand3_2 _47558_ (.A(_22367_),
    .B(_24254_),
    .C(_06548_),
    .Y(_15717_));
 sky130_as_sc_hs__nand3_2 _47562_ (.A(net100),
    .B(_15719_),
    .C(_15720_),
    .Y(_15721_));
 sky130_as_sc_hs__or2_2 _47563_ (.A(net1232),
    .B(net99),
    .Y(_15722_));
 sky130_as_sc_hs__and2_2 _47564_ (.A(net527),
    .B(net1233),
    .Y(_15723_));
 sky130_as_sc_hs__and2_2 _47565_ (.A(_15721_),
    .B(net1234),
    .Y(_01134_));
 sky130_as_sc_hs__or2_2 _47567_ (.A(_22622_),
    .B(_06548_),
    .Y(_15725_));
 sky130_as_sc_hs__nand3_2 _47568_ (.A(net144),
    .B(_15724_),
    .C(_15725_),
    .Y(_15726_));
 sky130_as_sc_hs__nand3_2 _47570_ (.A(net101),
    .B(_15726_),
    .C(_15727_),
    .Y(_15728_));
 sky130_as_sc_hs__or2_2 _47571_ (.A(net1179),
    .B(net101),
    .Y(_15729_));
 sky130_as_sc_hs__and2_2 _47572_ (.A(net527),
    .B(net1180),
    .Y(_15730_));
 sky130_as_sc_hs__and2_2 _47573_ (.A(_15728_),
    .B(net1181),
    .Y(_01135_));
 sky130_as_sc_hs__nand3_2 _47576_ (.A(net143),
    .B(_15731_),
    .C(_15732_),
    .Y(_15733_));
 sky130_as_sc_hs__nand3_2 _47578_ (.A(net100),
    .B(_15733_),
    .C(_15734_),
    .Y(_15735_));
 sky130_as_sc_hs__or2_2 _47579_ (.A(net1135),
    .B(net100),
    .Y(_15736_));
 sky130_as_sc_hs__and2_2 _47580_ (.A(net527),
    .B(net1136),
    .Y(_15737_));
 sky130_as_sc_hs__and2_2 _47581_ (.A(_15735_),
    .B(net1137),
    .Y(_01136_));
 sky130_as_sc_hs__nand3_2 _47584_ (.A(net143),
    .B(_15738_),
    .C(_15739_),
    .Y(_15740_));
 sky130_as_sc_hs__nand3_2 _47586_ (.A(net102),
    .B(_15740_),
    .C(_15741_),
    .Y(_15742_));
 sky130_as_sc_hs__or2_2 _47587_ (.A(net1283),
    .B(net102),
    .Y(_15743_));
 sky130_as_sc_hs__and2_2 _47588_ (.A(net498),
    .B(net1284),
    .Y(_15744_));
 sky130_as_sc_hs__and2_2 _47589_ (.A(_15742_),
    .B(net1285),
    .Y(_01137_));
 sky130_as_sc_hs__or2_2 _47591_ (.A(_22430_),
    .B(_06548_),
    .Y(_15746_));
 sky130_as_sc_hs__nand3_2 _47592_ (.A(net144),
    .B(_15745_),
    .C(_15746_),
    .Y(_15747_));
 sky130_as_sc_hs__nand3_2 _47594_ (.A(net101),
    .B(_15747_),
    .C(_15748_),
    .Y(_15749_));
 sky130_as_sc_hs__or2_2 _47595_ (.A(net1313),
    .B(_15290_),
    .Y(_15750_));
 sky130_as_sc_hs__and2_2 _47596_ (.A(net527),
    .B(net1314),
    .Y(_15751_));
 sky130_as_sc_hs__and2_2 _47597_ (.A(_15749_),
    .B(net1315),
    .Y(_01138_));
 sky130_as_sc_hs__nand3_2 _47600_ (.A(net144),
    .B(_15752_),
    .C(_15753_),
    .Y(_15754_));
 sky130_as_sc_hs__nand3_2 _47602_ (.A(_15290_),
    .B(_15754_),
    .C(_15755_),
    .Y(_15756_));
 sky130_as_sc_hs__or2_2 _47603_ (.A(net1192),
    .B(net101),
    .Y(_15757_));
 sky130_as_sc_hs__and2_2 _47604_ (.A(net527),
    .B(net1193),
    .Y(_15758_));
 sky130_as_sc_hs__and2_2 _47605_ (.A(_15756_),
    .B(net1194),
    .Y(_01139_));
 sky130_as_sc_hs__nand3_2 _47608_ (.A(net143),
    .B(_15759_),
    .C(_15760_),
    .Y(_15761_));
 sky130_as_sc_hs__nand3_2 _47610_ (.A(net102),
    .B(_15761_),
    .C(_15762_),
    .Y(_15763_));
 sky130_as_sc_hs__or2_2 _47611_ (.A(net1201),
    .B(net102),
    .Y(_15764_));
 sky130_as_sc_hs__and2_2 _47612_ (.A(net498),
    .B(net1202),
    .Y(_15765_));
 sky130_as_sc_hs__and2_2 _47613_ (.A(_15763_),
    .B(net1203),
    .Y(_01140_));
 sky130_as_sc_hs__or2_2 _47615_ (.A(_22687_),
    .B(_06548_),
    .Y(_15767_));
 sky130_as_sc_hs__nand3_2 _47616_ (.A(net144),
    .B(_15766_),
    .C(_15767_),
    .Y(_15768_));
 sky130_as_sc_hs__nand3_2 _47618_ (.A(net100),
    .B(_15768_),
    .C(_15769_),
    .Y(_15770_));
 sky130_as_sc_hs__or2_2 _47619_ (.A(net1155),
    .B(net100),
    .Y(_15771_));
 sky130_as_sc_hs__and2_2 _47620_ (.A(net527),
    .B(net1156),
    .Y(_15772_));
 sky130_as_sc_hs__and2_2 _47621_ (.A(_15770_),
    .B(net1157),
    .Y(_01141_));
 sky130_as_sc_hs__nand3_2 _47624_ (.A(net143),
    .B(_15773_),
    .C(_15774_),
    .Y(_15775_));
 sky130_as_sc_hs__nand3_2 _47626_ (.A(net99),
    .B(_15775_),
    .C(_15776_),
    .Y(_15777_));
 sky130_as_sc_hs__or2_2 _47627_ (.A(net1093),
    .B(net99),
    .Y(_15778_));
 sky130_as_sc_hs__and2_2 _47628_ (.A(net498),
    .B(net1094),
    .Y(_15779_));
 sky130_as_sc_hs__and2_2 _47629_ (.A(_15777_),
    .B(net1095),
    .Y(_01142_));
 sky130_as_sc_hs__or2_2 _47630_ (.A(_23672_),
    .B(_06549_),
    .Y(_15780_));
 sky130_as_sc_hs__nand3_2 _47632_ (.A(net143),
    .B(_15780_),
    .C(_15781_),
    .Y(_15782_));
 sky130_as_sc_hs__nand3_2 _47634_ (.A(net99),
    .B(_15782_),
    .C(_15783_),
    .Y(_15784_));
 sky130_as_sc_hs__or2_2 _47635_ (.A(net1079),
    .B(net99),
    .Y(_15785_));
 sky130_as_sc_hs__and2_2 _47636_ (.A(net498),
    .B(net1080),
    .Y(_15786_));
 sky130_as_sc_hs__and2_2 _47637_ (.A(_15784_),
    .B(net1081),
    .Y(_01143_));
 sky130_as_sc_hs__nand3_2 _47640_ (.A(net143),
    .B(_15787_),
    .C(_15788_),
    .Y(_15789_));
 sky130_as_sc_hs__nand3_2 _47642_ (.A(net102),
    .B(_15789_),
    .C(_15790_),
    .Y(_15791_));
 sky130_as_sc_hs__or2_2 _47643_ (.A(net1176),
    .B(net102),
    .Y(_15792_));
 sky130_as_sc_hs__and2_2 _47644_ (.A(net498),
    .B(net1177),
    .Y(_15793_));
 sky130_as_sc_hs__and2_2 _47645_ (.A(_15791_),
    .B(net1178),
    .Y(_01144_));
 sky130_as_sc_hs__nand3_2 _47648_ (.A(net143),
    .B(_15794_),
    .C(_15795_),
    .Y(_15796_));
 sky130_as_sc_hs__nand3_2 _47650_ (.A(net99),
    .B(_15796_),
    .C(_15797_),
    .Y(_15798_));
 sky130_as_sc_hs__or2_2 _47651_ (.A(net1307),
    .B(net99),
    .Y(_15799_));
 sky130_as_sc_hs__and2_2 _47652_ (.A(net498),
    .B(net1308),
    .Y(_15800_));
 sky130_as_sc_hs__and2_2 _47653_ (.A(_15798_),
    .B(net1309),
    .Y(_01145_));
 sky130_as_sc_hs__nand3_2 _47656_ (.A(net144),
    .B(_15801_),
    .C(_15802_),
    .Y(_15803_));
 sky130_as_sc_hs__nand3_2 _47658_ (.A(net101),
    .B(_15803_),
    .C(_15804_),
    .Y(_15805_));
 sky130_as_sc_hs__or2_2 _47659_ (.A(net1292),
    .B(net101),
    .Y(_15806_));
 sky130_as_sc_hs__and2_2 _47660_ (.A(net503),
    .B(net1293),
    .Y(_15807_));
 sky130_as_sc_hs__and2_2 _47661_ (.A(_15805_),
    .B(net1294),
    .Y(_01146_));
 sky130_as_sc_hs__nand3_2 _47664_ (.A(net143),
    .B(_15808_),
    .C(_15809_),
    .Y(_15810_));
 sky130_as_sc_hs__nand3_2 _47666_ (.A(net99),
    .B(_15810_),
    .C(_15811_),
    .Y(_15812_));
 sky130_as_sc_hs__or2_2 _47667_ (.A(net1226),
    .B(net100),
    .Y(_15813_));
 sky130_as_sc_hs__and2_2 _47668_ (.A(net498),
    .B(net1227),
    .Y(_15814_));
 sky130_as_sc_hs__and2_2 _47669_ (.A(_15812_),
    .B(net1228),
    .Y(_01147_));
 sky130_as_sc_hs__nand3_2 _47672_ (.A(net143),
    .B(_15815_),
    .C(_15816_),
    .Y(_15817_));
 sky130_as_sc_hs__nand3_2 _47674_ (.A(net100),
    .B(_15817_),
    .C(_15818_),
    .Y(_15819_));
 sky130_as_sc_hs__or2_2 _47675_ (.A(net1189),
    .B(net100),
    .Y(_15820_));
 sky130_as_sc_hs__and2_2 _47676_ (.A(net527),
    .B(net1190),
    .Y(_15821_));
 sky130_as_sc_hs__and2_2 _47677_ (.A(_15819_),
    .B(net1191),
    .Y(_01148_));
 sky130_as_sc_hs__nand3_2 _47680_ (.A(net144),
    .B(_15822_),
    .C(_15823_),
    .Y(_15824_));
 sky130_as_sc_hs__nand3_2 _47682_ (.A(net101),
    .B(_15824_),
    .C(_15825_),
    .Y(_15826_));
 sky130_as_sc_hs__or2_2 _47683_ (.A(net1298),
    .B(net101),
    .Y(_15827_));
 sky130_as_sc_hs__and2_2 _47684_ (.A(net503),
    .B(net1299),
    .Y(_15828_));
 sky130_as_sc_hs__and2_2 _47685_ (.A(_15826_),
    .B(net1300),
    .Y(_01149_));
 sky130_as_sc_hs__or2_2 _47687_ (.A(_23141_),
    .B(_06548_),
    .Y(_15830_));
 sky130_as_sc_hs__nand3_2 _47688_ (.A(net144),
    .B(_15829_),
    .C(_15830_),
    .Y(_15831_));
 sky130_as_sc_hs__nand3_2 _47690_ (.A(net99),
    .B(_15831_),
    .C(_15832_),
    .Y(_15833_));
 sky130_as_sc_hs__or2_2 _47691_ (.A(net1165),
    .B(net99),
    .Y(_15834_));
 sky130_as_sc_hs__and2_2 _47692_ (.A(net527),
    .B(net1166),
    .Y(_15835_));
 sky130_as_sc_hs__and2_2 _47693_ (.A(_15833_),
    .B(net1167),
    .Y(_01150_));
 sky130_as_sc_hs__nand3_2 _47696_ (.A(net143),
    .B(_15836_),
    .C(_15837_),
    .Y(_15838_));
 sky130_as_sc_hs__nand3_2 _47698_ (.A(net99),
    .B(_15838_),
    .C(_15839_),
    .Y(_15840_));
 sky130_as_sc_hs__or2_2 _47699_ (.A(net1304),
    .B(net99),
    .Y(_15841_));
 sky130_as_sc_hs__and2_2 _47700_ (.A(net498),
    .B(net1305),
    .Y(_15842_));
 sky130_as_sc_hs__and2_2 _47701_ (.A(_15840_),
    .B(net1306),
    .Y(_01151_));
 sky130_as_sc_hs__nand3_2 _47704_ (.A(net143),
    .B(_15843_),
    .C(_15844_),
    .Y(_15845_));
 sky130_as_sc_hs__nand3_2 _47706_ (.A(net102),
    .B(_15845_),
    .C(_15846_),
    .Y(_15847_));
 sky130_as_sc_hs__or2_2 _47707_ (.A(net1138),
    .B(net102),
    .Y(_15848_));
 sky130_as_sc_hs__and2_2 _47708_ (.A(net498),
    .B(net1139),
    .Y(_15849_));
 sky130_as_sc_hs__and2_2 _47709_ (.A(_15847_),
    .B(net1140),
    .Y(_01152_));
 sky130_as_sc_hs__nand3_2 _47712_ (.A(net144),
    .B(_15850_),
    .C(_15851_),
    .Y(_15852_));
 sky130_as_sc_hs__nand3_2 _47714_ (.A(net100),
    .B(_15852_),
    .C(_15853_),
    .Y(_15854_));
 sky130_as_sc_hs__or2_2 _47715_ (.A(net1223),
    .B(net100),
    .Y(_15855_));
 sky130_as_sc_hs__and2_2 _47716_ (.A(net527),
    .B(net1224),
    .Y(_15856_));
 sky130_as_sc_hs__and2_2 _47717_ (.A(_15854_),
    .B(net1225),
    .Y(_01153_));
 sky130_as_sc_hs__or2_2 _47719_ (.A(_23334_),
    .B(_06548_),
    .Y(_15858_));
 sky130_as_sc_hs__nand3_2 _47720_ (.A(net144),
    .B(_15857_),
    .C(_15858_),
    .Y(_15859_));
 sky130_as_sc_hs__nand3_2 _47722_ (.A(net101),
    .B(_15859_),
    .C(_15860_),
    .Y(_15861_));
 sky130_as_sc_hs__or2_2 _47723_ (.A(net1235),
    .B(net101),
    .Y(_15862_));
 sky130_as_sc_hs__and2_2 _47724_ (.A(net527),
    .B(net1236),
    .Y(_15863_));
 sky130_as_sc_hs__and2_2 _47725_ (.A(_15861_),
    .B(net1237),
    .Y(_01154_));
 sky130_as_sc_hs__or2_2 _47727_ (.A(_21723_),
    .B(_06548_),
    .Y(_15865_));
 sky130_as_sc_hs__nand3_2 _47728_ (.A(net143),
    .B(_15864_),
    .C(_15865_),
    .Y(_15866_));
 sky130_as_sc_hs__nand3_2 _47730_ (.A(net99),
    .B(_15866_),
    .C(_15867_),
    .Y(_15868_));
 sky130_as_sc_hs__or2_2 _47731_ (.A(net1208),
    .B(net99),
    .Y(_15869_));
 sky130_as_sc_hs__and2_2 _47732_ (.A(net498),
    .B(net1209),
    .Y(_15870_));
 sky130_as_sc_hs__and2_2 _47733_ (.A(_15868_),
    .B(net1210),
    .Y(_01155_));
 sky130_as_sc_hs__nand3_2 _47736_ (.A(net144),
    .B(_15871_),
    .C(_15872_),
    .Y(_15873_));
 sky130_as_sc_hs__nand3_2 _47738_ (.A(net101),
    .B(_15873_),
    .C(_15874_),
    .Y(_15875_));
 sky130_as_sc_hs__or2_2 _47739_ (.A(net1280),
    .B(net101),
    .Y(_15876_));
 sky130_as_sc_hs__and2_2 _47740_ (.A(net503),
    .B(net1281),
    .Y(_15877_));
 sky130_as_sc_hs__and2_2 _47741_ (.A(_15875_),
    .B(net1282),
    .Y(_01156_));
 sky130_as_sc_hs__nand3_2 _47744_ (.A(net144),
    .B(_15878_),
    .C(_15879_),
    .Y(_15880_));
 sky130_as_sc_hs__nand3_2 _47746_ (.A(net101),
    .B(_15880_),
    .C(_15881_),
    .Y(_15882_));
 sky130_as_sc_hs__or2_2 _47747_ (.A(net1254),
    .B(net101),
    .Y(_15883_));
 sky130_as_sc_hs__and2_2 _47748_ (.A(net503),
    .B(net1255),
    .Y(_15884_));
 sky130_as_sc_hs__and2_2 _47749_ (.A(_15882_),
    .B(net1256),
    .Y(_01157_));
 sky130_as_sc_hs__or2_2 _47750_ (.A(_02476_),
    .B(_06545_),
    .Y(_15885_));
 sky130_as_sc_hs__nand3_2 _47751_ (.A(net145),
    .B(_21655_),
    .C(_15885_),
    .Y(_15886_));
 sky130_as_sc_hs__nand3_2 _47753_ (.A(net102),
    .B(_15886_),
    .C(_15887_),
    .Y(_15888_));
 sky130_as_sc_hs__and2_2 _47755_ (.A(net497),
    .B(_15889_),
    .Y(_15890_));
 sky130_as_sc_hs__and2_2 _47756_ (.A(_15888_),
    .B(_15890_),
    .Y(_01158_));
 sky130_as_sc_hs__and2_2 _47758_ (.A(net116),
    .B(_15574_),
    .Y(_15892_));
 sky130_as_sc_hs__or2_2 _47760_ (.A(\tholin_riscv.div_shifter[31] ),
    .B(_15892_),
    .Y(_15894_));
 sky130_as_sc_hs__nand3_2 _47761_ (.A(net134),
    .B(_15893_),
    .C(_15894_),
    .Y(_15895_));
 sky130_as_sc_hs__and2_2 _47763_ (.A(net495),
    .B(_15896_),
    .Y(_01159_));
 sky130_as_sc_hs__or2_2 _47767_ (.A(\tholin_riscv.div_shifter[32] ),
    .B(_15574_),
    .Y(_15900_));
 sky130_as_sc_hs__nand3_2 _47769_ (.A(net134),
    .B(_15900_),
    .C(_15901_),
    .Y(_15902_));
 sky130_as_sc_hs__and2_2 _47771_ (.A(net495),
    .B(_15903_),
    .Y(_01160_));
 sky130_as_sc_hs__or2_2 _47773_ (.A(_15434_),
    .B(_15436_),
    .Y(_15905_));
 sky130_as_sc_hs__or2_2 _47776_ (.A(\tholin_riscv.div_shifter[33] ),
    .B(_15574_),
    .Y(_15908_));
 sky130_as_sc_hs__nand3_2 _47777_ (.A(net134),
    .B(_15907_),
    .C(_15908_),
    .Y(_15909_));
 sky130_as_sc_hs__and2_2 _47779_ (.A(net495),
    .B(_15910_),
    .Y(_01161_));
 sky130_as_sc_hs__or2_2 _47782_ (.A(_15438_),
    .B(_15566_),
    .Y(_15913_));
 sky130_as_sc_hs__or2_2 _47785_ (.A(\tholin_riscv.div_shifter[34] ),
    .B(_15574_),
    .Y(_15916_));
 sky130_as_sc_hs__nand3_2 _47786_ (.A(net134),
    .B(_15915_),
    .C(_15916_),
    .Y(_15917_));
 sky130_as_sc_hs__and2_2 _47788_ (.A(net495),
    .B(_15918_),
    .Y(_01162_));
 sky130_as_sc_hs__and2_2 _47790_ (.A(_15439_),
    .B(_15448_),
    .Y(_15920_));
 sky130_as_sc_hs__or2_2 _47791_ (.A(_15565_),
    .B(_15920_),
    .Y(_15921_));
 sky130_as_sc_hs__or2_2 _47794_ (.A(\tholin_riscv.div_shifter[35] ),
    .B(_15574_),
    .Y(_15924_));
 sky130_as_sc_hs__nand3_2 _47796_ (.A(net134),
    .B(_15924_),
    .C(_15925_),
    .Y(_15926_));
 sky130_as_sc_hs__and2_2 _47798_ (.A(net495),
    .B(_15927_),
    .Y(_01163_));
 sky130_as_sc_hs__or2_2 _47802_ (.A(_15564_),
    .B(_15929_),
    .Y(_15931_));
 sky130_as_sc_hs__or2_2 _47805_ (.A(\tholin_riscv.div_shifter[36] ),
    .B(_15574_),
    .Y(_15934_));
 sky130_as_sc_hs__nand3_2 _47806_ (.A(net134),
    .B(_15933_),
    .C(_15934_),
    .Y(_15935_));
 sky130_as_sc_hs__and2_2 _47808_ (.A(net495),
    .B(_15936_),
    .Y(_01164_));
 sky130_as_sc_hs__or2_2 _47813_ (.A(_15563_),
    .B(_15939_),
    .Y(_15941_));
 sky130_as_sc_hs__or2_2 _47815_ (.A(\tholin_riscv.div_shifter[37] ),
    .B(_15574_),
    .Y(_15943_));
 sky130_as_sc_hs__nand3_2 _47817_ (.A(net134),
    .B(_15943_),
    .C(_15944_),
    .Y(_15945_));
 sky130_as_sc_hs__and2_2 _47819_ (.A(net495),
    .B(_15946_),
    .Y(_01165_));
 sky130_as_sc_hs__or2_2 _47823_ (.A(_15562_),
    .B(_15948_),
    .Y(_15950_));
 sky130_as_sc_hs__nand3_2 _47824_ (.A(_15574_),
    .B(_15949_),
    .C(_15950_),
    .Y(_15951_));
 sky130_as_sc_hs__or2_2 _47825_ (.A(\tholin_riscv.div_shifter[38] ),
    .B(_15574_),
    .Y(_15952_));
 sky130_as_sc_hs__nand3_2 _47826_ (.A(net134),
    .B(_15951_),
    .C(_15952_),
    .Y(_15953_));
 sky130_as_sc_hs__and2_2 _47828_ (.A(net489),
    .B(_15954_),
    .Y(_01166_));
 sky130_as_sc_hs__or2_2 _47833_ (.A(_15409_),
    .B(_15957_),
    .Y(_15959_));
 sky130_as_sc_hs__or2_2 _47835_ (.A(\tholin_riscv.div_shifter[39] ),
    .B(_15574_),
    .Y(_15961_));
 sky130_as_sc_hs__nand3_2 _47837_ (.A(net133),
    .B(_15961_),
    .C(_15962_),
    .Y(_15963_));
 sky130_as_sc_hs__and2_2 _47839_ (.A(net489),
    .B(_15964_),
    .Y(_01167_));
 sky130_as_sc_hs__or2_2 _47843_ (.A(_15403_),
    .B(_15966_),
    .Y(_15968_));
 sky130_as_sc_hs__or2_2 _47846_ (.A(\tholin_riscv.div_shifter[40] ),
    .B(_15574_),
    .Y(_15971_));
 sky130_as_sc_hs__nand3_2 _47847_ (.A(net133),
    .B(_15970_),
    .C(_15971_),
    .Y(_15972_));
 sky130_as_sc_hs__and2_2 _47849_ (.A(net489),
    .B(_15973_),
    .Y(_01168_));
 sky130_as_sc_hs__or2_2 _47854_ (.A(_15397_),
    .B(_15976_),
    .Y(_15978_));
 sky130_as_sc_hs__or2_2 _47856_ (.A(\tholin_riscv.div_shifter[41] ),
    .B(_15574_),
    .Y(_15980_));
 sky130_as_sc_hs__nand3_2 _47858_ (.A(net133),
    .B(_15980_),
    .C(_15981_),
    .Y(_15982_));
 sky130_as_sc_hs__and2_2 _47860_ (.A(net489),
    .B(_15983_),
    .Y(_01169_));
 sky130_as_sc_hs__and2_2 _47862_ (.A(_15396_),
    .B(_15977_),
    .Y(_15985_));
 sky130_as_sc_hs__or2_2 _47863_ (.A(_15391_),
    .B(_15985_),
    .Y(_15986_));
 sky130_as_sc_hs__nand3_2 _47865_ (.A(_15574_),
    .B(_15986_),
    .C(_15987_),
    .Y(_15988_));
 sky130_as_sc_hs__or2_2 _47866_ (.A(\tholin_riscv.div_shifter[42] ),
    .B(_15574_),
    .Y(_15989_));
 sky130_as_sc_hs__nand3_2 _47867_ (.A(net133),
    .B(_15988_),
    .C(_15989_),
    .Y(_15990_));
 sky130_as_sc_hs__and2_2 _47869_ (.A(net488),
    .B(_15991_),
    .Y(_01170_));
 sky130_as_sc_hs__and2_2 _47872_ (.A(_15389_),
    .B(_15993_),
    .Y(_15994_));
 sky130_as_sc_hs__or2_2 _47873_ (.A(_15385_),
    .B(_15994_),
    .Y(_15995_));
 sky130_as_sc_hs__or2_2 _47877_ (.A(\tholin_riscv.div_shifter[43] ),
    .B(_15574_),
    .Y(_15999_));
 sky130_as_sc_hs__nand3_2 _47878_ (.A(net133),
    .B(_15998_),
    .C(_15999_),
    .Y(_16000_));
 sky130_as_sc_hs__and2_2 _47880_ (.A(net488),
    .B(_16001_),
    .Y(_01171_));
 sky130_as_sc_hs__and2_2 _47882_ (.A(_15384_),
    .B(_15996_),
    .Y(_16003_));
 sky130_as_sc_hs__or2_2 _47884_ (.A(_15379_),
    .B(_16003_),
    .Y(_16005_));
 sky130_as_sc_hs__nand3_2 _47885_ (.A(_15574_),
    .B(_16004_),
    .C(_16005_),
    .Y(_16006_));
 sky130_as_sc_hs__or2_2 _47886_ (.A(\tholin_riscv.div_shifter[44] ),
    .B(_15574_),
    .Y(_16007_));
 sky130_as_sc_hs__nand3_2 _47887_ (.A(net133),
    .B(_16006_),
    .C(_16007_),
    .Y(_16008_));
 sky130_as_sc_hs__and2_2 _47889_ (.A(net488),
    .B(_16009_),
    .Y(_01172_));
 sky130_as_sc_hs__and2_2 _47892_ (.A(_15378_),
    .B(_16011_),
    .Y(_16012_));
 sky130_as_sc_hs__or2_2 _47893_ (.A(_15542_),
    .B(_16012_),
    .Y(_16013_));
 sky130_as_sc_hs__or2_2 _47897_ (.A(\tholin_riscv.div_shifter[45] ),
    .B(_15574_),
    .Y(_16017_));
 sky130_as_sc_hs__nand3_2 _47898_ (.A(net133),
    .B(_16016_),
    .C(_16017_),
    .Y(_16018_));
 sky130_as_sc_hs__and2_2 _47900_ (.A(net488),
    .B(_16019_),
    .Y(_01173_));
 sky130_as_sc_hs__or2_2 _47903_ (.A(_15541_),
    .B(_16021_),
    .Y(_16022_));
 sky130_as_sc_hs__nand3_2 _47905_ (.A(_15574_),
    .B(_16022_),
    .C(_16023_),
    .Y(_16024_));
 sky130_as_sc_hs__or2_2 _47906_ (.A(\tholin_riscv.div_shifter[46] ),
    .B(_15574_),
    .Y(_16025_));
 sky130_as_sc_hs__nand3_2 _47907_ (.A(net133),
    .B(_16024_),
    .C(_16025_),
    .Y(_16026_));
 sky130_as_sc_hs__and2_2 _47909_ (.A(net486),
    .B(_16027_),
    .Y(_01174_));
 sky130_as_sc_hs__or2_2 _47913_ (.A(_15533_),
    .B(_16030_),
    .Y(_16031_));
 sky130_as_sc_hs__or2_2 _47917_ (.A(\tholin_riscv.div_shifter[47] ),
    .B(_15574_),
    .Y(_16035_));
 sky130_as_sc_hs__nand3_2 _47918_ (.A(net132),
    .B(_16034_),
    .C(_16035_),
    .Y(_16036_));
 sky130_as_sc_hs__and2_2 _47920_ (.A(net486),
    .B(_16037_),
    .Y(_01175_));
 sky130_as_sc_hs__nor2_2 _47923_ (.A(_15526_),
    .B(_16039_),
    .Y(_16040_));
 sky130_as_sc_hs__or2_2 _47926_ (.A(_16040_),
    .B(_16042_),
    .Y(_16043_));
 sky130_as_sc_hs__or2_2 _47927_ (.A(\tholin_riscv.div_shifter[48] ),
    .B(_15574_),
    .Y(_16044_));
 sky130_as_sc_hs__nand3_2 _47928_ (.A(net132),
    .B(_16043_),
    .C(_16044_),
    .Y(_16045_));
 sky130_as_sc_hs__and2_2 _47930_ (.A(net486),
    .B(_16046_),
    .Y(_01176_));
 sky130_as_sc_hs__or2_2 _47935_ (.A(_15519_),
    .B(_16049_),
    .Y(_16051_));
 sky130_as_sc_hs__or2_2 _47938_ (.A(\tholin_riscv.div_shifter[49] ),
    .B(_15574_),
    .Y(_16054_));
 sky130_as_sc_hs__nand3_2 _47939_ (.A(net132),
    .B(_16053_),
    .C(_16054_),
    .Y(_16055_));
 sky130_as_sc_hs__and2_2 _47941_ (.A(net486),
    .B(_16056_),
    .Y(_01177_));
 sky130_as_sc_hs__and2_2 _47943_ (.A(_15518_),
    .B(_16050_),
    .Y(_16058_));
 sky130_as_sc_hs__or2_2 _47945_ (.A(_15513_),
    .B(_16058_),
    .Y(_16060_));
 sky130_as_sc_hs__nand3_2 _47946_ (.A(_15574_),
    .B(_16059_),
    .C(_16060_),
    .Y(_16061_));
 sky130_as_sc_hs__or2_2 _47947_ (.A(\tholin_riscv.div_shifter[50] ),
    .B(_15574_),
    .Y(_16062_));
 sky130_as_sc_hs__nand3_2 _47948_ (.A(net132),
    .B(_16061_),
    .C(_16062_),
    .Y(_16063_));
 sky130_as_sc_hs__and2_2 _47950_ (.A(net486),
    .B(_16064_),
    .Y(_01178_));
 sky130_as_sc_hs__and2_2 _47953_ (.A(_15512_),
    .B(_16066_),
    .Y(_16067_));
 sky130_as_sc_hs__or2_2 _47955_ (.A(_15507_),
    .B(_16067_),
    .Y(_16069_));
 sky130_as_sc_hs__or2_2 _47958_ (.A(\tholin_riscv.div_shifter[51] ),
    .B(_15574_),
    .Y(_16072_));
 sky130_as_sc_hs__nand3_2 _47959_ (.A(net132),
    .B(_16071_),
    .C(_16072_),
    .Y(_16073_));
 sky130_as_sc_hs__and2_2 _47961_ (.A(net486),
    .B(_16074_),
    .Y(_01179_));
 sky130_as_sc_hs__and2_2 _47963_ (.A(_15506_),
    .B(_16068_),
    .Y(_16076_));
 sky130_as_sc_hs__or2_2 _47965_ (.A(_15501_),
    .B(_16076_),
    .Y(_16078_));
 sky130_as_sc_hs__nand3_2 _47966_ (.A(_15574_),
    .B(_16077_),
    .C(_16078_),
    .Y(_16079_));
 sky130_as_sc_hs__or2_2 _47967_ (.A(\tholin_riscv.div_shifter[52] ),
    .B(_15574_),
    .Y(_16080_));
 sky130_as_sc_hs__nand3_2 _47968_ (.A(net132),
    .B(_16079_),
    .C(_16080_),
    .Y(_16081_));
 sky130_as_sc_hs__and2_2 _47970_ (.A(net486),
    .B(_16082_),
    .Y(_01180_));
 sky130_as_sc_hs__or2_2 _47974_ (.A(_15495_),
    .B(_16085_),
    .Y(_16086_));
 sky130_as_sc_hs__or2_2 _47978_ (.A(\tholin_riscv.div_shifter[53] ),
    .B(_15574_),
    .Y(_16090_));
 sky130_as_sc_hs__nand3_2 _47979_ (.A(net132),
    .B(_16089_),
    .C(_16090_),
    .Y(_16091_));
 sky130_as_sc_hs__and2_2 _47981_ (.A(net486),
    .B(_16092_),
    .Y(_01181_));
 sky130_as_sc_hs__nor2_2 _47984_ (.A(_15489_),
    .B(_16094_),
    .Y(_16095_));
 sky130_as_sc_hs__or2_2 _47987_ (.A(_16095_),
    .B(_16097_),
    .Y(_16098_));
 sky130_as_sc_hs__or2_2 _47988_ (.A(\tholin_riscv.div_shifter[54] ),
    .B(_15574_),
    .Y(_16099_));
 sky130_as_sc_hs__nand3_2 _47989_ (.A(net132),
    .B(_16098_),
    .C(_16099_),
    .Y(_16100_));
 sky130_as_sc_hs__and2_2 _47991_ (.A(net486),
    .B(_16101_),
    .Y(_01182_));
 sky130_as_sc_hs__or2_2 _47996_ (.A(_15342_),
    .B(_16104_),
    .Y(_16106_));
 sky130_as_sc_hs__or2_2 _47999_ (.A(\tholin_riscv.div_shifter[55] ),
    .B(_15574_),
    .Y(_16109_));
 sky130_as_sc_hs__nand3_2 _48000_ (.A(net132),
    .B(_16108_),
    .C(_16109_),
    .Y(_16110_));
 sky130_as_sc_hs__and2_2 _48002_ (.A(net486),
    .B(_16111_),
    .Y(_01183_));
 sky130_as_sc_hs__nor2_2 _48005_ (.A(_15349_),
    .B(_16113_),
    .Y(_16114_));
 sky130_as_sc_hs__or2_2 _48008_ (.A(_16114_),
    .B(_16116_),
    .Y(_16117_));
 sky130_as_sc_hs__or2_2 _48009_ (.A(\tholin_riscv.div_shifter[56] ),
    .B(_15574_),
    .Y(_16118_));
 sky130_as_sc_hs__nand3_2 _48010_ (.A(net132),
    .B(_16117_),
    .C(_16118_),
    .Y(_16119_));
 sky130_as_sc_hs__and2_2 _48012_ (.A(net486),
    .B(_16120_),
    .Y(_01184_));
 sky130_as_sc_hs__or2_2 _48017_ (.A(_15355_),
    .B(_16123_),
    .Y(_16125_));
 sky130_as_sc_hs__or2_2 _48020_ (.A(\tholin_riscv.div_shifter[57] ),
    .B(_15574_),
    .Y(_16128_));
 sky130_as_sc_hs__nand3_2 _48021_ (.A(net132),
    .B(_16127_),
    .C(_16128_),
    .Y(_16129_));
 sky130_as_sc_hs__and2_2 _48023_ (.A(net485),
    .B(_16130_),
    .Y(_01185_));
 sky130_as_sc_hs__or2_2 _48026_ (.A(_15336_),
    .B(_16132_),
    .Y(_16133_));
 sky130_as_sc_hs__nand3_2 _48028_ (.A(_15574_),
    .B(_16133_),
    .C(_16134_),
    .Y(_16135_));
 sky130_as_sc_hs__or2_2 _48029_ (.A(\tholin_riscv.div_shifter[58] ),
    .B(_15574_),
    .Y(_16136_));
 sky130_as_sc_hs__nand3_2 _48030_ (.A(net132),
    .B(_16135_),
    .C(_16136_),
    .Y(_16137_));
 sky130_as_sc_hs__and2_2 _48032_ (.A(net485),
    .B(_16138_),
    .Y(_01186_));
 sky130_as_sc_hs__or2_2 _48037_ (.A(_15364_),
    .B(_16141_),
    .Y(_16143_));
 sky130_as_sc_hs__or2_2 _48040_ (.A(\tholin_riscv.div_shifter[59] ),
    .B(_15574_),
    .Y(_16146_));
 sky130_as_sc_hs__nand3_2 _48041_ (.A(net132),
    .B(_16145_),
    .C(_16146_),
    .Y(_16147_));
 sky130_as_sc_hs__and2_2 _48043_ (.A(net485),
    .B(_16148_),
    .Y(_01187_));
 sky130_as_sc_hs__or2_2 _48047_ (.A(_15370_),
    .B(_16150_),
    .Y(_16152_));
 sky130_as_sc_hs__or2_2 _48050_ (.A(\tholin_riscv.div_shifter[60] ),
    .B(_15574_),
    .Y(_16155_));
 sky130_as_sc_hs__nand3_2 _48051_ (.A(net132),
    .B(_16154_),
    .C(_16155_),
    .Y(_16156_));
 sky130_as_sc_hs__and2_2 _48053_ (.A(net485),
    .B(_16157_),
    .Y(_01188_));
 sky130_as_sc_hs__or2_2 _48058_ (.A(_15325_),
    .B(_16160_),
    .Y(_16162_));
 sky130_as_sc_hs__or2_2 _48061_ (.A(\tholin_riscv.div_shifter[61] ),
    .B(_15574_),
    .Y(_16165_));
 sky130_as_sc_hs__nand3_2 _48062_ (.A(net132),
    .B(_16164_),
    .C(_16165_),
    .Y(_16166_));
 sky130_as_sc_hs__and2_2 _48064_ (.A(net485),
    .B(_16167_),
    .Y(_01189_));
 sky130_as_sc_hs__or2_2 _48069_ (.A(\tholin_riscv.div_shifter[62] ),
    .B(_15574_),
    .Y(_16172_));
 sky130_as_sc_hs__nand3_2 _48070_ (.A(net132),
    .B(_16171_),
    .C(_16172_),
    .Y(_16173_));
 sky130_as_sc_hs__and2_2 _48072_ (.A(net496),
    .B(_16174_),
    .Y(_01190_));
 sky130_as_sc_hs__or2_2 _48074_ (.A(net639),
    .B(_15275_),
    .Y(_16176_));
 sky130_as_sc_hs__and2_2 _48075_ (.A(_16175_),
    .B(net640),
    .Y(_01191_));
 sky130_as_sc_hs__and2_2 _48076_ (.A(net542),
    .B(net768),
    .Y(_16177_));
 sky130_as_sc_hs__and2_2 _48077_ (.A(net967),
    .B(_16177_),
    .Y(_16178_));
 sky130_as_sc_hs__and2_2 _48078_ (.A(net1020),
    .B(_16178_),
    .Y(_16179_));
 sky130_as_sc_hs__and2_2 _48079_ (.A(net822),
    .B(_16179_),
    .Y(_16180_));
 sky130_as_sc_hs__and2_2 _48080_ (.A(net851),
    .B(_16180_),
    .Y(_16181_));
 sky130_as_sc_hs__and2_2 _48081_ (.A(net1000),
    .B(_16181_),
    .Y(_16182_));
 sky130_as_sc_hs__and2_2 _48082_ (.A(net1024),
    .B(_16182_),
    .Y(_16183_));
 sky130_as_sc_hs__and2_2 _48083_ (.A(net1016),
    .B(_16183_),
    .Y(_16184_));
 sky130_as_sc_hs__and2_2 _48084_ (.A(net947),
    .B(_16184_),
    .Y(_16185_));
 sky130_as_sc_hs__and2_2 _48085_ (.A(net1049),
    .B(_16185_),
    .Y(_16186_));
 sky130_as_sc_hs__and2_2 _48086_ (.A(net1012),
    .B(_16186_),
    .Y(_16187_));
 sky130_as_sc_hs__and2_2 _48087_ (.A(net1123),
    .B(_16187_),
    .Y(_16188_));
 sky130_as_sc_hs__and2_2 _48088_ (.A(net843),
    .B(_16188_),
    .Y(_16189_));
 sky130_as_sc_hs__and2_2 _48089_ (.A(net943),
    .B(_16189_),
    .Y(_16190_));
 sky130_as_sc_hs__and2_2 _48090_ (.A(net907),
    .B(_16190_),
    .Y(_16191_));
 sky130_as_sc_hs__and2_2 _48091_ (.A(net859),
    .B(_16191_),
    .Y(_16192_));
 sky130_as_sc_hs__and2_2 _48092_ (.A(net867),
    .B(_16192_),
    .Y(_16193_));
 sky130_as_sc_hs__and2_2 _48093_ (.A(net895),
    .B(_16193_),
    .Y(_16194_));
 sky130_as_sc_hs__and2_2 _48094_ (.A(net863),
    .B(_16194_),
    .Y(_16195_));
 sky130_as_sc_hs__and2_2 _48095_ (.A(net1045),
    .B(_16195_),
    .Y(_16196_));
 sky130_as_sc_hs__and2_2 _48096_ (.A(net1204),
    .B(_16196_),
    .Y(_16197_));
 sky130_as_sc_hs__and2_2 _48097_ (.A(net903),
    .B(_16197_),
    .Y(_16198_));
 sky130_as_sc_hs__and2_2 _48098_ (.A(net810),
    .B(_16198_),
    .Y(_16199_));
 sky130_as_sc_hs__and2_2 _48099_ (.A(net915),
    .B(_16199_),
    .Y(_16200_));
 sky130_as_sc_hs__and2_2 _48100_ (.A(net764),
    .B(_16200_),
    .Y(_16201_));
 sky130_as_sc_hs__and2_2 _48101_ (.A(net939),
    .B(_16201_),
    .Y(_16202_));
 sky130_as_sc_hs__and2_2 _48102_ (.A(net988),
    .B(_16202_),
    .Y(_16203_));
 sky130_as_sc_hs__and2_2 _48103_ (.A(net1089),
    .B(_16203_),
    .Y(_16204_));
 sky130_as_sc_hs__and2_2 _48104_ (.A(net1061),
    .B(_16204_),
    .Y(_16205_));
 sky130_as_sc_hs__and2_2 _48105_ (.A(net787),
    .B(_16205_),
    .Y(_16206_));
 sky130_as_sc_hs__or2_2 _48106_ (.A(\tholin_riscv.tmr1_pre_ctr[31] ),
    .B(_16206_),
    .Y(_16207_));
 sky130_as_sc_hs__nor2_2 _48110_ (.A(net1045),
    .B(_16195_),
    .Y(_16211_));
 sky130_as_sc_hs__or2_2 _48111_ (.A(_16196_),
    .B(net1046),
    .Y(_16212_));
 sky130_as_sc_hs__nor2_2 _48113_ (.A(net863),
    .B(_16194_),
    .Y(_16214_));
 sky130_as_sc_hs__or2_2 _48114_ (.A(_16195_),
    .B(net864),
    .Y(_16215_));
 sky130_as_sc_hs__or2_2 _48115_ (.A(\tholin_riscv.tmr1_pre[19] ),
    .B(_16215_),
    .Y(_16216_));
 sky130_as_sc_hs__nor2_2 _48116_ (.A(net943),
    .B(_16189_),
    .Y(_16217_));
 sky130_as_sc_hs__or2_2 _48117_ (.A(_16190_),
    .B(net944),
    .Y(_16218_));
 sky130_as_sc_hs__or2_2 _48118_ (.A(\tholin_riscv.tmr1_pre[14] ),
    .B(_16218_),
    .Y(_16219_));
 sky130_as_sc_hs__nor2_2 _48119_ (.A(net843),
    .B(_16188_),
    .Y(_16220_));
 sky130_as_sc_hs__or2_2 _48120_ (.A(_16189_),
    .B(net844),
    .Y(_16221_));
 sky130_as_sc_hs__nor2_2 _48122_ (.A(net1123),
    .B(_16187_),
    .Y(_16223_));
 sky130_as_sc_hs__or2_2 _48123_ (.A(_16188_),
    .B(net1124),
    .Y(_16224_));
 sky130_as_sc_hs__nor2_2 _48125_ (.A(net822),
    .B(_16179_),
    .Y(_16226_));
 sky130_as_sc_hs__or2_2 _48126_ (.A(_16180_),
    .B(net823),
    .Y(_16227_));
 sky130_as_sc_hs__or2_2 _48127_ (.A(\tholin_riscv.tmr1_pre[4] ),
    .B(_16227_),
    .Y(_16228_));
 sky130_as_sc_hs__nor2_2 _48128_ (.A(net1020),
    .B(_16178_),
    .Y(_16229_));
 sky130_as_sc_hs__or2_2 _48129_ (.A(_16179_),
    .B(net1021),
    .Y(_16230_));
 sky130_as_sc_hs__or2_2 _48130_ (.A(\tholin_riscv.tmr1_pre[3] ),
    .B(_16230_),
    .Y(_16231_));
 sky130_as_sc_hs__nor2_2 _48132_ (.A(net967),
    .B(_16177_),
    .Y(_16233_));
 sky130_as_sc_hs__or2_2 _48133_ (.A(_16178_),
    .B(net968),
    .Y(_16234_));
 sky130_as_sc_hs__or2_2 _48134_ (.A(\tholin_riscv.tmr1_pre[2] ),
    .B(_16234_),
    .Y(_16235_));
 sky130_as_sc_hs__nor2_2 _48136_ (.A(net542),
    .B(net768),
    .Y(_16237_));
 sky130_as_sc_hs__or2_2 _48137_ (.A(_16177_),
    .B(net769),
    .Y(_16238_));
 sky130_as_sc_hs__or2_2 _48138_ (.A(\tholin_riscv.tmr1_pre[1] ),
    .B(_16238_),
    .Y(_16239_));
 sky130_as_sc_hs__nand3_2 _48142_ (.A(_16235_),
    .B(_16239_),
    .C(_16242_),
    .Y(_16243_));
 sky130_as_sc_hs__nand3_2 _48143_ (.A(_16232_),
    .B(_16236_),
    .C(_16243_),
    .Y(_16244_));
 sky130_as_sc_hs__nand3_2 _48144_ (.A(_16228_),
    .B(_16231_),
    .C(_16244_),
    .Y(_16245_));
 sky130_as_sc_hs__nor2_2 _48145_ (.A(net851),
    .B(_16180_),
    .Y(_16246_));
 sky130_as_sc_hs__or2_2 _48146_ (.A(_16181_),
    .B(net852),
    .Y(_16247_));
 sky130_as_sc_hs__nand3_2 _48149_ (.A(_16245_),
    .B(_16248_),
    .C(_16249_),
    .Y(_16250_));
 sky130_as_sc_hs__or2_2 _48150_ (.A(\tholin_riscv.tmr1_pre[5] ),
    .B(_16247_),
    .Y(_16251_));
 sky130_as_sc_hs__nor2_2 _48151_ (.A(net1000),
    .B(_16181_),
    .Y(_16252_));
 sky130_as_sc_hs__or2_2 _48152_ (.A(_16182_),
    .B(net1001),
    .Y(_16253_));
 sky130_as_sc_hs__or2_2 _48153_ (.A(\tholin_riscv.tmr1_pre[6] ),
    .B(_16253_),
    .Y(_16254_));
 sky130_as_sc_hs__nand3_2 _48154_ (.A(_16250_),
    .B(_16251_),
    .C(_16254_),
    .Y(_16255_));
 sky130_as_sc_hs__nor2_2 _48156_ (.A(net1024),
    .B(_16182_),
    .Y(_16257_));
 sky130_as_sc_hs__or2_2 _48157_ (.A(_16183_),
    .B(net1025),
    .Y(_16258_));
 sky130_as_sc_hs__nand3_2 _48159_ (.A(_16255_),
    .B(_16256_),
    .C(_16259_),
    .Y(_16260_));
 sky130_as_sc_hs__or2_2 _48160_ (.A(\tholin_riscv.tmr1_pre[7] ),
    .B(_16258_),
    .Y(_16261_));
 sky130_as_sc_hs__nor2_2 _48161_ (.A(net1016),
    .B(_16183_),
    .Y(_16262_));
 sky130_as_sc_hs__or2_2 _48162_ (.A(_16184_),
    .B(net1017),
    .Y(_16263_));
 sky130_as_sc_hs__or2_2 _48163_ (.A(\tholin_riscv.tmr1_pre[8] ),
    .B(_16263_),
    .Y(_16264_));
 sky130_as_sc_hs__nand3_2 _48164_ (.A(_16260_),
    .B(_16261_),
    .C(_16264_),
    .Y(_16265_));
 sky130_as_sc_hs__nor2_2 _48166_ (.A(net947),
    .B(_16184_),
    .Y(_16267_));
 sky130_as_sc_hs__or2_2 _48167_ (.A(_16185_),
    .B(net948),
    .Y(_16268_));
 sky130_as_sc_hs__nand3_2 _48169_ (.A(_16265_),
    .B(_16266_),
    .C(_16269_),
    .Y(_16270_));
 sky130_as_sc_hs__or2_2 _48170_ (.A(\tholin_riscv.tmr1_pre[9] ),
    .B(_16268_),
    .Y(_16271_));
 sky130_as_sc_hs__nor2_2 _48171_ (.A(net1049),
    .B(_16185_),
    .Y(_16272_));
 sky130_as_sc_hs__or2_2 _48172_ (.A(_16186_),
    .B(net1050),
    .Y(_16273_));
 sky130_as_sc_hs__or2_2 _48173_ (.A(\tholin_riscv.tmr1_pre[10] ),
    .B(_16273_),
    .Y(_16274_));
 sky130_as_sc_hs__nand3_2 _48174_ (.A(_16270_),
    .B(_16271_),
    .C(_16274_),
    .Y(_16275_));
 sky130_as_sc_hs__nor2_2 _48176_ (.A(net1012),
    .B(_16186_),
    .Y(_16277_));
 sky130_as_sc_hs__or2_2 _48177_ (.A(_16187_),
    .B(net1013),
    .Y(_16278_));
 sky130_as_sc_hs__nand3_2 _48179_ (.A(_16275_),
    .B(_16276_),
    .C(_16279_),
    .Y(_16280_));
 sky130_as_sc_hs__or2_2 _48180_ (.A(\tholin_riscv.tmr1_pre[12] ),
    .B(_16224_),
    .Y(_16281_));
 sky130_as_sc_hs__or2_2 _48181_ (.A(\tholin_riscv.tmr1_pre[11] ),
    .B(_16278_),
    .Y(_16282_));
 sky130_as_sc_hs__nand3_2 _48182_ (.A(_16280_),
    .B(_16281_),
    .C(_16282_),
    .Y(_16283_));
 sky130_as_sc_hs__or2_2 _48184_ (.A(\tholin_riscv.tmr1_pre[13] ),
    .B(_16221_),
    .Y(_16285_));
 sky130_as_sc_hs__nor2_2 _48188_ (.A(net907),
    .B(_16190_),
    .Y(_16289_));
 sky130_as_sc_hs__or2_2 _48189_ (.A(_16191_),
    .B(net908),
    .Y(_16290_));
 sky130_as_sc_hs__nand3_2 _48192_ (.A(_16288_),
    .B(_16291_),
    .C(_16292_),
    .Y(_16293_));
 sky130_as_sc_hs__or2_2 _48193_ (.A(\tholin_riscv.tmr1_pre[15] ),
    .B(_16290_),
    .Y(_16294_));
 sky130_as_sc_hs__nor2_2 _48194_ (.A(net859),
    .B(_16191_),
    .Y(_16295_));
 sky130_as_sc_hs__or2_2 _48195_ (.A(_16192_),
    .B(net860),
    .Y(_16296_));
 sky130_as_sc_hs__or2_2 _48196_ (.A(\tholin_riscv.tmr1_pre[16] ),
    .B(_16296_),
    .Y(_16297_));
 sky130_as_sc_hs__nand3_2 _48197_ (.A(_16293_),
    .B(_16294_),
    .C(_16297_),
    .Y(_16298_));
 sky130_as_sc_hs__nor2_2 _48199_ (.A(net867),
    .B(_16192_),
    .Y(_16300_));
 sky130_as_sc_hs__or2_2 _48200_ (.A(_16193_),
    .B(net868),
    .Y(_16301_));
 sky130_as_sc_hs__nand3_2 _48202_ (.A(_16298_),
    .B(_16299_),
    .C(_16302_),
    .Y(_16303_));
 sky130_as_sc_hs__nor2_2 _48203_ (.A(net895),
    .B(_16193_),
    .Y(_16304_));
 sky130_as_sc_hs__or2_2 _48204_ (.A(_16194_),
    .B(net896),
    .Y(_16305_));
 sky130_as_sc_hs__or2_2 _48205_ (.A(\tholin_riscv.tmr1_pre[18] ),
    .B(_16305_),
    .Y(_16306_));
 sky130_as_sc_hs__or2_2 _48206_ (.A(\tholin_riscv.tmr1_pre[17] ),
    .B(_16301_),
    .Y(_16307_));
 sky130_as_sc_hs__nand3_2 _48207_ (.A(_16303_),
    .B(_16306_),
    .C(_16307_),
    .Y(_16308_));
 sky130_as_sc_hs__nand3_2 _48210_ (.A(_16308_),
    .B(_16309_),
    .C(_16310_),
    .Y(_16311_));
 sky130_as_sc_hs__nor2_2 _48213_ (.A(net1204),
    .B(_16196_),
    .Y(_16314_));
 sky130_as_sc_hs__or2_2 _48214_ (.A(_16197_),
    .B(net1205),
    .Y(_16315_));
 sky130_as_sc_hs__or2_2 _48215_ (.A(\tholin_riscv.tmr1_pre[21] ),
    .B(_16315_),
    .Y(_16316_));
 sky130_as_sc_hs__or2_2 _48216_ (.A(\tholin_riscv.tmr1_pre[20] ),
    .B(_16212_),
    .Y(_16317_));
 sky130_as_sc_hs__nand3_2 _48217_ (.A(_16313_),
    .B(_16316_),
    .C(_16317_),
    .Y(_16318_));
 sky130_as_sc_hs__nor2_2 _48218_ (.A(net903),
    .B(_16197_),
    .Y(_16319_));
 sky130_as_sc_hs__or2_2 _48219_ (.A(_16198_),
    .B(net904),
    .Y(_16320_));
 sky130_as_sc_hs__nand3_2 _48222_ (.A(_16318_),
    .B(_16321_),
    .C(_16322_),
    .Y(_16323_));
 sky130_as_sc_hs__nor2_2 _48223_ (.A(net810),
    .B(_16198_),
    .Y(_16324_));
 sky130_as_sc_hs__or2_2 _48224_ (.A(_16199_),
    .B(net811),
    .Y(_16325_));
 sky130_as_sc_hs__or2_2 _48225_ (.A(\tholin_riscv.tmr1_pre[23] ),
    .B(_16325_),
    .Y(_16326_));
 sky130_as_sc_hs__or2_2 _48226_ (.A(\tholin_riscv.tmr1_pre[22] ),
    .B(_16320_),
    .Y(_16327_));
 sky130_as_sc_hs__nand3_2 _48227_ (.A(_16323_),
    .B(_16326_),
    .C(_16327_),
    .Y(_16328_));
 sky130_as_sc_hs__nor2_2 _48228_ (.A(net915),
    .B(_16199_),
    .Y(_16329_));
 sky130_as_sc_hs__or2_2 _48229_ (.A(_16200_),
    .B(net916),
    .Y(_16330_));
 sky130_as_sc_hs__or2_2 _48232_ (.A(\tholin_riscv.tmr1_pre[24] ),
    .B(_16330_),
    .Y(_16333_));
 sky130_as_sc_hs__nor2_2 _48233_ (.A(net764),
    .B(_16200_),
    .Y(_16334_));
 sky130_as_sc_hs__nor2_2 _48234_ (.A(_16201_),
    .B(net765),
    .Y(_16335_));
 sky130_as_sc_hs__nor2_2 _48235_ (.A(net939),
    .B(_16201_),
    .Y(_16336_));
 sky130_as_sc_hs__or2_2 _48236_ (.A(_16202_),
    .B(net940),
    .Y(_16337_));
 sky130_as_sc_hs__nor2_2 _48238_ (.A(net988),
    .B(_16202_),
    .Y(_16339_));
 sky130_as_sc_hs__or2_2 _48239_ (.A(_16203_),
    .B(net989),
    .Y(_16340_));
 sky130_as_sc_hs__or2_2 _48240_ (.A(\tholin_riscv.tmr1_pre[27] ),
    .B(_16340_),
    .Y(_16341_));
 sky130_as_sc_hs__or2_2 _48241_ (.A(\tholin_riscv.tmr1_pre[26] ),
    .B(_16337_),
    .Y(_16342_));
 sky130_as_sc_hs__or2_2 _48247_ (.A(\tholin_riscv.tmr1_pre[25] ),
    .B(_16345_),
    .Y(_16348_));
 sky130_as_sc_hs__nand3_2 _48248_ (.A(_16342_),
    .B(_16347_),
    .C(_16348_),
    .Y(_16349_));
 sky130_as_sc_hs__nor2_2 _48251_ (.A(net1089),
    .B(_16203_),
    .Y(_16352_));
 sky130_as_sc_hs__or2_2 _48252_ (.A(_16204_),
    .B(net1090),
    .Y(_16353_));
 sky130_as_sc_hs__nand3_2 _48255_ (.A(_16351_),
    .B(_16354_),
    .C(_16355_),
    .Y(_16356_));
 sky130_as_sc_hs__nor2_2 _48256_ (.A(net1061),
    .B(_16204_),
    .Y(_16357_));
 sky130_as_sc_hs__or2_2 _48257_ (.A(_16205_),
    .B(net1062),
    .Y(_16358_));
 sky130_as_sc_hs__or2_2 _48258_ (.A(\tholin_riscv.tmr1_pre[29] ),
    .B(_16358_),
    .Y(_16359_));
 sky130_as_sc_hs__or2_2 _48259_ (.A(\tholin_riscv.tmr1_pre[28] ),
    .B(_16353_),
    .Y(_16360_));
 sky130_as_sc_hs__nand3_2 _48260_ (.A(_16356_),
    .B(_16359_),
    .C(_16360_),
    .Y(_16361_));
 sky130_as_sc_hs__nor2_2 _48261_ (.A(net787),
    .B(_16205_),
    .Y(_16362_));
 sky130_as_sc_hs__or2_2 _48262_ (.A(net788),
    .B(_16362_),
    .Y(_16363_));
 sky130_as_sc_hs__nand3_2 _48265_ (.A(_16361_),
    .B(_16364_),
    .C(_16365_),
    .Y(_16366_));
 sky130_as_sc_hs__or2_2 _48266_ (.A(\tholin_riscv.tmr1_pre[31] ),
    .B(_16209_),
    .Y(_16367_));
 sky130_as_sc_hs__or2_2 _48267_ (.A(\tholin_riscv.tmr1_pre[30] ),
    .B(_16363_),
    .Y(_16368_));
 sky130_as_sc_hs__nand3_2 _48268_ (.A(_16366_),
    .B(_16367_),
    .C(_16368_),
    .Y(_16369_));
 sky130_as_sc_hs__inv_2 _48271_ (.Y(_16372_),
    .A(_16371_));
 sky130_as_sc_hs__nor2_2 _48272_ (.A(net1711),
    .B(_16371_),
    .Y(_01192_));
 sky130_as_sc_hs__nor2_2 _48273_ (.A(net770),
    .B(_16371_),
    .Y(_01193_));
 sky130_as_sc_hs__nor2_2 _48274_ (.A(net969),
    .B(_16371_),
    .Y(_01194_));
 sky130_as_sc_hs__nor2_2 _48275_ (.A(net1022),
    .B(_16371_),
    .Y(_01195_));
 sky130_as_sc_hs__nor2_2 _48276_ (.A(net824),
    .B(_16371_),
    .Y(_01196_));
 sky130_as_sc_hs__nor2_2 _48277_ (.A(net853),
    .B(_16371_),
    .Y(_01197_));
 sky130_as_sc_hs__nor2_2 _48278_ (.A(net1002),
    .B(_16371_),
    .Y(_01198_));
 sky130_as_sc_hs__nor2_2 _48279_ (.A(net1026),
    .B(_16371_),
    .Y(_01199_));
 sky130_as_sc_hs__nor2_2 _48280_ (.A(net1018),
    .B(_16371_),
    .Y(_01200_));
 sky130_as_sc_hs__nor2_2 _48281_ (.A(net949),
    .B(_16371_),
    .Y(_01201_));
 sky130_as_sc_hs__nor2_2 _48282_ (.A(net1051),
    .B(_16371_),
    .Y(_01202_));
 sky130_as_sc_hs__nor2_2 _48283_ (.A(net1014),
    .B(_16371_),
    .Y(_01203_));
 sky130_as_sc_hs__nor2_2 _48284_ (.A(net1125),
    .B(_16371_),
    .Y(_01204_));
 sky130_as_sc_hs__nor2_2 _48285_ (.A(net845),
    .B(_16371_),
    .Y(_01205_));
 sky130_as_sc_hs__nor2_2 _48286_ (.A(net945),
    .B(_16371_),
    .Y(_01206_));
 sky130_as_sc_hs__nor2_2 _48287_ (.A(net909),
    .B(_16371_),
    .Y(_01207_));
 sky130_as_sc_hs__nor2_2 _48288_ (.A(net861),
    .B(_16371_),
    .Y(_01208_));
 sky130_as_sc_hs__nor2_2 _48289_ (.A(net869),
    .B(_16371_),
    .Y(_01209_));
 sky130_as_sc_hs__nor2_2 _48290_ (.A(net897),
    .B(_16371_),
    .Y(_01210_));
 sky130_as_sc_hs__nor2_2 _48291_ (.A(net865),
    .B(_16371_),
    .Y(_01211_));
 sky130_as_sc_hs__nor2_2 _48292_ (.A(net1047),
    .B(_16371_),
    .Y(_01212_));
 sky130_as_sc_hs__nor2_2 _48293_ (.A(net1206),
    .B(_16371_),
    .Y(_01213_));
 sky130_as_sc_hs__nor2_2 _48294_ (.A(net905),
    .B(_16371_),
    .Y(_01214_));
 sky130_as_sc_hs__nor2_2 _48295_ (.A(net812),
    .B(_16371_),
    .Y(_01215_));
 sky130_as_sc_hs__nor2_2 _48296_ (.A(net917),
    .B(_16371_),
    .Y(_01216_));
 sky130_as_sc_hs__and2_2 _48297_ (.A(net766),
    .B(_16372_),
    .Y(_01217_));
 sky130_as_sc_hs__nor2_2 _48298_ (.A(net941),
    .B(_16371_),
    .Y(_01218_));
 sky130_as_sc_hs__nor2_2 _48299_ (.A(net990),
    .B(_16371_),
    .Y(_01219_));
 sky130_as_sc_hs__nor2_2 _48300_ (.A(net1091),
    .B(_16371_),
    .Y(_01220_));
 sky130_as_sc_hs__nor2_2 _48301_ (.A(net1063),
    .B(_16371_),
    .Y(_01221_));
 sky130_as_sc_hs__nor2_2 _48302_ (.A(net789),
    .B(_16371_),
    .Y(_01222_));
 sky130_as_sc_hs__nor2_2 _48303_ (.A(_16209_),
    .B(_16371_),
    .Y(_01223_));
 sky130_as_sc_hs__nand3_2 _48304_ (.A(_19973_),
    .B(_19977_),
    .C(_20012_),
    .Y(_16373_));
 sky130_as_sc_hs__and2_2 _48305_ (.A(_19749_),
    .B(_15314_),
    .Y(_16374_));
 sky130_as_sc_hs__or2_2 _48306_ (.A(_21563_),
    .B(_16374_),
    .Y(_16375_));
 sky130_as_sc_hs__and2_2 _48309_ (.A(_19942_),
    .B(_16377_),
    .Y(_16378_));
 sky130_as_sc_hs__and2_2 _48310_ (.A(_16373_),
    .B(_16378_),
    .Y(_16379_));
 sky130_as_sc_hs__or2_2 _48311_ (.A(_20009_),
    .B(_05509_),
    .Y(_16380_));
 sky130_as_sc_hs__nor2_2 _48314_ (.A(net371),
    .B(_19755_),
    .Y(_16383_));
 sky130_as_sc_hs__nor2_2 _48315_ (.A(_19750_),
    .B(_16383_),
    .Y(_16384_));
 sky130_as_sc_hs__nand3_2 _48318_ (.A(_16379_),
    .B(_16382_),
    .C(_16386_),
    .Y(_16387_));
 sky130_as_sc_hs__or2_2 _48319_ (.A(net1705),
    .B(_16379_),
    .Y(_16388_));
 sky130_as_sc_hs__and2_2 _48320_ (.A(net494),
    .B(_16388_),
    .Y(_16389_));
 sky130_as_sc_hs__and2_2 _48321_ (.A(_16387_),
    .B(_16389_),
    .Y(_01224_));
 sky130_as_sc_hs__or2_2 _48322_ (.A(_19495_),
    .B(_16384_),
    .Y(_16390_));
 sky130_as_sc_hs__or2_2 _48323_ (.A(\tholin_riscv.ret_cycle[1] ),
    .B(_19899_),
    .Y(_16391_));
 sky130_as_sc_hs__or2_2 _48324_ (.A(_19995_),
    .B(net134),
    .Y(_16392_));
 sky130_as_sc_hs__or2_2 _48326_ (.A(net1644),
    .B(_16379_),
    .Y(_16394_));
 sky130_as_sc_hs__nand3_2 _48327_ (.A(_16379_),
    .B(_16390_),
    .C(_16393_),
    .Y(_16395_));
 sky130_as_sc_hs__and2_2 _48328_ (.A(net494),
    .B(_16395_),
    .Y(_16396_));
 sky130_as_sc_hs__and2_2 _48329_ (.A(net1645),
    .B(_16396_),
    .Y(_01225_));
 sky130_as_sc_hs__and2_2 _48330_ (.A(_19755_),
    .B(_19761_),
    .Y(_16397_));
 sky130_as_sc_hs__and2_2 _48331_ (.A(_19751_),
    .B(_16397_),
    .Y(_16398_));
 sky130_as_sc_hs__or2_2 _48333_ (.A(_16383_),
    .B(_16397_),
    .Y(_16400_));
 sky130_as_sc_hs__or2_2 _48336_ (.A(_19497_),
    .B(_16379_),
    .Y(_16403_));
 sky130_as_sc_hs__and2_2 _48338_ (.A(net495),
    .B(_16404_),
    .Y(_01226_));
 sky130_as_sc_hs__nand3_2 _48339_ (.A(_21565_),
    .B(_15288_),
    .C(_16379_),
    .Y(_16405_));
 sky130_as_sc_hs__and2_2 _48341_ (.A(net494),
    .B(_16406_),
    .Y(_01227_));
 sky130_as_sc_hs__nor2_2 _48342_ (.A(\tholin_riscv.Bimm[5] ),
    .B(\tholin_riscv.Iimm[4] ),
    .Y(_16407_));
 sky130_as_sc_hs__nand3_2 _48343_ (.A(_19983_),
    .B(_19984_),
    .C(_16407_),
    .Y(_16408_));
 sky130_as_sc_hs__nand3_2 _48344_ (.A(_19479_),
    .B(\tholin_riscv.Iimm[1] ),
    .C(_13057_),
    .Y(_16409_));
 sky130_as_sc_hs__nor2_2 _48345_ (.A(\tholin_riscv.Iimm[2] ),
    .B(\tholin_riscv.Iimm[0] ),
    .Y(_16410_));
 sky130_as_sc_hs__and2_2 _48347_ (.A(_16409_),
    .B(_16411_),
    .Y(_16412_));
 sky130_as_sc_hs__or2_2 _48348_ (.A(_16408_),
    .B(_16412_),
    .Y(_16413_));
 sky130_as_sc_hs__nand3_2 _48349_ (.A(net145),
    .B(_13062_),
    .C(_16413_),
    .Y(_16414_));
 sky130_as_sc_hs__nor2_2 _48350_ (.A(_19943_),
    .B(_20010_),
    .Y(_16415_));
 sky130_as_sc_hs__and2_2 _48351_ (.A(_16414_),
    .B(_16415_),
    .Y(_16416_));
 sky130_as_sc_hs__or2_2 _48352_ (.A(net757),
    .B(_16416_),
    .Y(_16417_));
 sky130_as_sc_hs__or2_2 _48353_ (.A(\tholin_riscv.int_enabled ),
    .B(_13062_),
    .Y(_16418_));
 sky130_as_sc_hs__or2_2 _48354_ (.A(_16408_),
    .B(_16409_),
    .Y(_16419_));
 sky130_as_sc_hs__and2_2 _48358_ (.A(net502),
    .B(_16422_),
    .Y(_16423_));
 sky130_as_sc_hs__and2_2 _48359_ (.A(net758),
    .B(_16423_),
    .Y(_01228_));
 sky130_as_sc_hs__or2_2 _48360_ (.A(\tholin_riscv.cycle[2] ),
    .B(\tholin_riscv.cycle[1] ),
    .Y(_16424_));
 sky130_as_sc_hs__and2_2 _48363_ (.A(_19933_),
    .B(_19950_),
    .Y(_16427_));
 sky130_as_sc_hs__and2_2 _48364_ (.A(_16426_),
    .B(_16427_),
    .Y(_16428_));
 sky130_as_sc_hs__and2_2 _48366_ (.A(net1173),
    .B(_16429_),
    .Y(_16430_));
 sky130_as_sc_hs__or2_2 _48367_ (.A(_15274_),
    .B(net1174),
    .Y(_16431_));
 sky130_as_sc_hs__and2_2 _48368_ (.A(net501),
    .B(net1175),
    .Y(_01229_));
 sky130_as_sc_hs__and2_2 _48369_ (.A(_19937_),
    .B(_16428_),
    .Y(_16432_));
 sky130_as_sc_hs__and2_2 _48372_ (.A(net495),
    .B(_16434_),
    .Y(_16435_));
 sky130_as_sc_hs__and2_2 _48373_ (.A(_16433_),
    .B(_16435_),
    .Y(_01230_));
 sky130_as_sc_hs__and2_2 _48377_ (.A(net501),
    .B(_16438_),
    .Y(_01231_));
 sky130_as_sc_hs__and2_2 _48378_ (.A(_19486_),
    .B(_16432_),
    .Y(_16439_));
 sky130_as_sc_hs__or2_2 _48379_ (.A(net371),
    .B(_16428_),
    .Y(_16440_));
 sky130_as_sc_hs__nor2_2 _48381_ (.A(_16439_),
    .B(_16441_),
    .Y(_01232_));
 sky130_as_sc_hs__nand3_2 _48383_ (.A(_19950_),
    .B(_16397_),
    .C(_16442_),
    .Y(_16443_));
 sky130_as_sc_hs__nor2_2 _48384_ (.A(_20016_),
    .B(_16443_),
    .Y(_16444_));
 sky130_as_sc_hs__nand3_2 _48385_ (.A(_20015_),
    .B(_20019_),
    .C(_16444_),
    .Y(_16445_));
 sky130_as_sc_hs__or2_2 _48387_ (.A(net3),
    .B(_19751_),
    .Y(_16447_));
 sky130_as_sc_hs__nand3_2 _48388_ (.A(_19759_),
    .B(_16446_),
    .C(_16447_),
    .Y(_16448_));
 sky130_as_sc_hs__nand3_2 _48393_ (.A(_16450_),
    .B(_16451_),
    .C(_16452_),
    .Y(_16453_));
 sky130_as_sc_hs__and2_2 _48396_ (.A(_16454_),
    .B(_16455_),
    .Y(_16456_));
 sky130_as_sc_hs__nand3_2 _48399_ (.A(_16456_),
    .B(_16457_),
    .C(_16458_),
    .Y(_16459_));
 sky130_as_sc_hs__or2_2 _48400_ (.A(_16453_),
    .B(_16459_),
    .Y(_16460_));
 sky130_as_sc_hs__or2_2 _48401_ (.A(_16449_),
    .B(_16460_),
    .Y(_16461_));
 sky130_as_sc_hs__or2_2 _48402_ (.A(\tholin_riscv.intr_vec[14] ),
    .B(_20005_),
    .Y(_16462_));
 sky130_as_sc_hs__nand3_2 _48403_ (.A(net137),
    .B(_16461_),
    .C(_16462_),
    .Y(_16463_));
 sky130_as_sc_hs__or2_2 _48405_ (.A(_16445_),
    .B(_16464_),
    .Y(_16465_));
 sky130_as_sc_hs__and2_2 _48407_ (.A(net498),
    .B(_16466_),
    .Y(_16467_));
 sky130_as_sc_hs__and2_2 _48408_ (.A(_16465_),
    .B(_16467_),
    .Y(_01233_));
 sky130_as_sc_hs__or2_2 _48410_ (.A(net10),
    .B(_19751_),
    .Y(_16469_));
 sky130_as_sc_hs__nand3_2 _48411_ (.A(_19759_),
    .B(_16468_),
    .C(_16469_),
    .Y(_16470_));
 sky130_as_sc_hs__nand3_2 _48415_ (.A(_16471_),
    .B(_16472_),
    .C(_16473_),
    .Y(_16474_));
 sky130_as_sc_hs__and2_2 _48418_ (.A(_16475_),
    .B(_16476_),
    .Y(_16477_));
 sky130_as_sc_hs__nand3_2 _48421_ (.A(_16477_),
    .B(_16478_),
    .C(_16479_),
    .Y(_16480_));
 sky130_as_sc_hs__nor2_2 _48422_ (.A(_16474_),
    .B(_16480_),
    .Y(_16481_));
 sky130_as_sc_hs__and2_2 _48425_ (.A(net137),
    .B(_16483_),
    .Y(_16484_));
 sky130_as_sc_hs__nor2_2 _48426_ (.A(_16445_),
    .B(_16484_),
    .Y(_16485_));
 sky130_as_sc_hs__and2_2 _48429_ (.A(net526),
    .B(_16487_),
    .Y(_16488_));
 sky130_as_sc_hs__and2_2 _48430_ (.A(_16486_),
    .B(_16488_),
    .Y(_01234_));
 sky130_as_sc_hs__or2_2 _48432_ (.A(net13),
    .B(_19751_),
    .Y(_16490_));
 sky130_as_sc_hs__nand3_2 _48433_ (.A(_19759_),
    .B(_16489_),
    .C(_16490_),
    .Y(_16491_));
 sky130_as_sc_hs__nand3_2 _48437_ (.A(_16492_),
    .B(_16493_),
    .C(_16494_),
    .Y(_16495_));
 sky130_as_sc_hs__and2_2 _48440_ (.A(_16496_),
    .B(_16497_),
    .Y(_16498_));
 sky130_as_sc_hs__nand3_2 _48443_ (.A(_16498_),
    .B(_16499_),
    .C(_16500_),
    .Y(_16501_));
 sky130_as_sc_hs__nor2_2 _48444_ (.A(_16495_),
    .B(_16501_),
    .Y(_16502_));
 sky130_as_sc_hs__and2_2 _48447_ (.A(net137),
    .B(_16504_),
    .Y(_16505_));
 sky130_as_sc_hs__nor2_2 _48448_ (.A(_16445_),
    .B(_16505_),
    .Y(_16506_));
 sky130_as_sc_hs__and2_2 _48451_ (.A(net504),
    .B(_16508_),
    .Y(_16509_));
 sky130_as_sc_hs__and2_2 _48452_ (.A(_16507_),
    .B(_16509_),
    .Y(_01235_));
 sky130_as_sc_hs__or2_2 _48454_ (.A(net15),
    .B(_19751_),
    .Y(_16511_));
 sky130_as_sc_hs__nand3_2 _48455_ (.A(_19759_),
    .B(_16510_),
    .C(_16511_),
    .Y(_16512_));
 sky130_as_sc_hs__nand3_2 _48459_ (.A(_16513_),
    .B(_16514_),
    .C(_16515_),
    .Y(_16516_));
 sky130_as_sc_hs__and2_2 _48462_ (.A(_16517_),
    .B(_16518_),
    .Y(_16519_));
 sky130_as_sc_hs__nand3_2 _48465_ (.A(_16519_),
    .B(_16520_),
    .C(_16521_),
    .Y(_16522_));
 sky130_as_sc_hs__or2_2 _48466_ (.A(_16516_),
    .B(_16522_),
    .Y(_16523_));
 sky130_as_sc_hs__or2_2 _48467_ (.A(_16449_),
    .B(_16523_),
    .Y(_16524_));
 sky130_as_sc_hs__or2_2 _48468_ (.A(\tholin_riscv.intr_vec[17] ),
    .B(_20005_),
    .Y(_16525_));
 sky130_as_sc_hs__nand3_2 _48469_ (.A(net137),
    .B(_16524_),
    .C(_16525_),
    .Y(_16526_));
 sky130_as_sc_hs__and2_2 _48470_ (.A(_16512_),
    .B(_16526_),
    .Y(_16527_));
 sky130_as_sc_hs__or2_2 _48471_ (.A(_16445_),
    .B(_16527_),
    .Y(_16528_));
 sky130_as_sc_hs__and2_2 _48474_ (.A(net527),
    .B(_16530_),
    .Y(_01236_));
 sky130_as_sc_hs__or2_2 _48476_ (.A(net16),
    .B(_19751_),
    .Y(_16532_));
 sky130_as_sc_hs__nand3_2 _48477_ (.A(_19759_),
    .B(_16531_),
    .C(_16532_),
    .Y(_16533_));
 sky130_as_sc_hs__nand3_2 _48481_ (.A(_16534_),
    .B(_16535_),
    .C(_16536_),
    .Y(_16537_));
 sky130_as_sc_hs__and2_2 _48484_ (.A(_16538_),
    .B(_16539_),
    .Y(_16540_));
 sky130_as_sc_hs__nand3_2 _48487_ (.A(_16540_),
    .B(_16541_),
    .C(_16542_),
    .Y(_16543_));
 sky130_as_sc_hs__nor2_2 _48488_ (.A(_16537_),
    .B(_16543_),
    .Y(_16544_));
 sky130_as_sc_hs__and2_2 _48492_ (.A(_16533_),
    .B(_16547_),
    .Y(_16548_));
 sky130_as_sc_hs__or2_2 _48493_ (.A(_16445_),
    .B(_16548_),
    .Y(_16549_));
 sky130_as_sc_hs__and2_2 _48496_ (.A(net504),
    .B(_16551_),
    .Y(_01237_));
 sky130_as_sc_hs__or2_2 _48498_ (.A(net17),
    .B(_19751_),
    .Y(_16553_));
 sky130_as_sc_hs__nand3_2 _48499_ (.A(_19759_),
    .B(_16552_),
    .C(_16553_),
    .Y(_16554_));
 sky130_as_sc_hs__nand3_2 _48503_ (.A(_16555_),
    .B(_16556_),
    .C(_16557_),
    .Y(_16558_));
 sky130_as_sc_hs__and2_2 _48506_ (.A(_16559_),
    .B(_16560_),
    .Y(_16561_));
 sky130_as_sc_hs__nand3_2 _48509_ (.A(_16561_),
    .B(_16562_),
    .C(_16563_),
    .Y(_16564_));
 sky130_as_sc_hs__nor2_2 _48510_ (.A(_16558_),
    .B(_16564_),
    .Y(_16565_));
 sky130_as_sc_hs__and2_2 _48513_ (.A(net137),
    .B(_16567_),
    .Y(_16568_));
 sky130_as_sc_hs__nor2_2 _48514_ (.A(_16445_),
    .B(_16568_),
    .Y(_16569_));
 sky130_as_sc_hs__and2_2 _48517_ (.A(net503),
    .B(_16571_),
    .Y(_16572_));
 sky130_as_sc_hs__and2_2 _48518_ (.A(_16570_),
    .B(_16572_),
    .Y(_01238_));
 sky130_as_sc_hs__or2_2 _48520_ (.A(net18),
    .B(_19751_),
    .Y(_16574_));
 sky130_as_sc_hs__nand3_2 _48521_ (.A(_19759_),
    .B(_16573_),
    .C(_16574_),
    .Y(_16575_));
 sky130_as_sc_hs__nand3_2 _48525_ (.A(_16576_),
    .B(_16577_),
    .C(_16578_),
    .Y(_16579_));
 sky130_as_sc_hs__and2_2 _48528_ (.A(_16580_),
    .B(_16581_),
    .Y(_16582_));
 sky130_as_sc_hs__nand3_2 _48531_ (.A(_16582_),
    .B(_16583_),
    .C(_16584_),
    .Y(_16585_));
 sky130_as_sc_hs__or2_2 _48532_ (.A(_16579_),
    .B(_16585_),
    .Y(_16586_));
 sky130_as_sc_hs__or2_2 _48533_ (.A(_16449_),
    .B(_16586_),
    .Y(_16587_));
 sky130_as_sc_hs__or2_2 _48534_ (.A(\tholin_riscv.intr_vec[20] ),
    .B(_20005_),
    .Y(_16588_));
 sky130_as_sc_hs__nand3_2 _48535_ (.A(net137),
    .B(_16587_),
    .C(_16588_),
    .Y(_16589_));
 sky130_as_sc_hs__and2_2 _48536_ (.A(_16575_),
    .B(_16589_),
    .Y(_16590_));
 sky130_as_sc_hs__or2_2 _48537_ (.A(_16445_),
    .B(_16590_),
    .Y(_16591_));
 sky130_as_sc_hs__and2_2 _48540_ (.A(net520),
    .B(_16593_),
    .Y(_01239_));
 sky130_as_sc_hs__or2_2 _48542_ (.A(net19),
    .B(_19751_),
    .Y(_16595_));
 sky130_as_sc_hs__nand3_2 _48543_ (.A(_19759_),
    .B(_16594_),
    .C(_16595_),
    .Y(_16596_));
 sky130_as_sc_hs__nand3_2 _48547_ (.A(_16597_),
    .B(_16598_),
    .C(_16599_),
    .Y(_16600_));
 sky130_as_sc_hs__and2_2 _48550_ (.A(_16601_),
    .B(_16602_),
    .Y(_16603_));
 sky130_as_sc_hs__nand3_2 _48553_ (.A(_16603_),
    .B(_16604_),
    .C(_16605_),
    .Y(_16606_));
 sky130_as_sc_hs__nor2_2 _48554_ (.A(_16600_),
    .B(_16606_),
    .Y(_16607_));
 sky130_as_sc_hs__and2_2 _48557_ (.A(net137),
    .B(_16609_),
    .Y(_16610_));
 sky130_as_sc_hs__nor2_2 _48558_ (.A(_16445_),
    .B(_16610_),
    .Y(_16611_));
 sky130_as_sc_hs__and2_2 _48561_ (.A(net503),
    .B(_16613_),
    .Y(_16614_));
 sky130_as_sc_hs__and2_2 _48562_ (.A(_16612_),
    .B(_16614_),
    .Y(_01240_));
 sky130_as_sc_hs__or2_2 _48564_ (.A(net20),
    .B(_19751_),
    .Y(_16616_));
 sky130_as_sc_hs__nand3_2 _48565_ (.A(_19759_),
    .B(_16615_),
    .C(_16616_),
    .Y(_16617_));
 sky130_as_sc_hs__nand3_2 _48569_ (.A(_16618_),
    .B(_16619_),
    .C(_16620_),
    .Y(_16621_));
 sky130_as_sc_hs__and2_2 _48572_ (.A(_16622_),
    .B(_16623_),
    .Y(_16624_));
 sky130_as_sc_hs__nand3_2 _48575_ (.A(_16624_),
    .B(_16625_),
    .C(_16626_),
    .Y(_16627_));
 sky130_as_sc_hs__nor2_2 _48576_ (.A(_16621_),
    .B(_16627_),
    .Y(_16628_));
 sky130_as_sc_hs__and2_2 _48579_ (.A(net137),
    .B(_16630_),
    .Y(_16631_));
 sky130_as_sc_hs__nor2_2 _48580_ (.A(_16445_),
    .B(_16631_),
    .Y(_16632_));
 sky130_as_sc_hs__and2_2 _48583_ (.A(net503),
    .B(_16634_),
    .Y(_16635_));
 sky130_as_sc_hs__and2_2 _48584_ (.A(_16633_),
    .B(_16635_),
    .Y(_01241_));
 sky130_as_sc_hs__or2_2 _48586_ (.A(net21),
    .B(_19751_),
    .Y(_16637_));
 sky130_as_sc_hs__nand3_2 _48587_ (.A(_19759_),
    .B(_16636_),
    .C(_16637_),
    .Y(_16638_));
 sky130_as_sc_hs__nand3_2 _48591_ (.A(_16639_),
    .B(_16640_),
    .C(_16641_),
    .Y(_16642_));
 sky130_as_sc_hs__and2_2 _48594_ (.A(_16643_),
    .B(_16644_),
    .Y(_16645_));
 sky130_as_sc_hs__nand3_2 _48597_ (.A(_16645_),
    .B(_16646_),
    .C(_16647_),
    .Y(_16648_));
 sky130_as_sc_hs__or2_2 _48598_ (.A(_16642_),
    .B(_16648_),
    .Y(_16649_));
 sky130_as_sc_hs__or2_2 _48599_ (.A(_16449_),
    .B(_16649_),
    .Y(_16650_));
 sky130_as_sc_hs__or2_2 _48600_ (.A(\tholin_riscv.intr_vec[23] ),
    .B(_20005_),
    .Y(_16651_));
 sky130_as_sc_hs__nand3_2 _48601_ (.A(net137),
    .B(_16650_),
    .C(_16651_),
    .Y(_16652_));
 sky130_as_sc_hs__and2_2 _48602_ (.A(_16638_),
    .B(_16652_),
    .Y(_16653_));
 sky130_as_sc_hs__or2_2 _48603_ (.A(_16445_),
    .B(_16653_),
    .Y(_16654_));
 sky130_as_sc_hs__and2_2 _48606_ (.A(net504),
    .B(_16656_),
    .Y(_01242_));
 sky130_as_sc_hs__or2_2 _48608_ (.A(net4),
    .B(_19751_),
    .Y(_16658_));
 sky130_as_sc_hs__nand3_2 _48609_ (.A(_19759_),
    .B(_16657_),
    .C(_16658_),
    .Y(_16659_));
 sky130_as_sc_hs__nand3_2 _48613_ (.A(_16660_),
    .B(_16661_),
    .C(_16662_),
    .Y(_16663_));
 sky130_as_sc_hs__and2_2 _48616_ (.A(_16664_),
    .B(_16665_),
    .Y(_16666_));
 sky130_as_sc_hs__nand3_2 _48619_ (.A(_16666_),
    .B(_16667_),
    .C(_16668_),
    .Y(_16669_));
 sky130_as_sc_hs__nor2_2 _48620_ (.A(_16663_),
    .B(_16669_),
    .Y(_16670_));
 sky130_as_sc_hs__and2_2 _48624_ (.A(_16659_),
    .B(_16673_),
    .Y(_16674_));
 sky130_as_sc_hs__or2_2 _48625_ (.A(_16445_),
    .B(_16674_),
    .Y(_16675_));
 sky130_as_sc_hs__and2_2 _48628_ (.A(net511),
    .B(_16677_),
    .Y(_01243_));
 sky130_as_sc_hs__or2_2 _48630_ (.A(net5),
    .B(_19751_),
    .Y(_16679_));
 sky130_as_sc_hs__nand3_2 _48631_ (.A(_19759_),
    .B(_16678_),
    .C(_16679_),
    .Y(_16680_));
 sky130_as_sc_hs__nand3_2 _48635_ (.A(_16681_),
    .B(_16682_),
    .C(_16683_),
    .Y(_16684_));
 sky130_as_sc_hs__and2_2 _48638_ (.A(_16685_),
    .B(_16686_),
    .Y(_16687_));
 sky130_as_sc_hs__nand3_2 _48641_ (.A(_16687_),
    .B(_16688_),
    .C(_16689_),
    .Y(_16690_));
 sky130_as_sc_hs__nor2_2 _48642_ (.A(_16684_),
    .B(_16690_),
    .Y(_16691_));
 sky130_as_sc_hs__and2_2 _48645_ (.A(net137),
    .B(_16693_),
    .Y(_16694_));
 sky130_as_sc_hs__nor2_2 _48646_ (.A(_16445_),
    .B(_16694_),
    .Y(_16695_));
 sky130_as_sc_hs__and2_2 _48649_ (.A(net503),
    .B(_16697_),
    .Y(_16698_));
 sky130_as_sc_hs__and2_2 _48650_ (.A(_16696_),
    .B(_16698_),
    .Y(_01244_));
 sky130_as_sc_hs__or2_2 _48652_ (.A(net6),
    .B(_19751_),
    .Y(_16700_));
 sky130_as_sc_hs__nand3_2 _48653_ (.A(_19759_),
    .B(_16699_),
    .C(_16700_),
    .Y(_16701_));
 sky130_as_sc_hs__nand3_2 _48657_ (.A(_16702_),
    .B(_16703_),
    .C(_16704_),
    .Y(_16705_));
 sky130_as_sc_hs__and2_2 _48660_ (.A(_16706_),
    .B(_16707_),
    .Y(_16708_));
 sky130_as_sc_hs__nand3_2 _48663_ (.A(_16708_),
    .B(_16709_),
    .C(_16710_),
    .Y(_16711_));
 sky130_as_sc_hs__or2_2 _48664_ (.A(_16705_),
    .B(_16711_),
    .Y(_16712_));
 sky130_as_sc_hs__or2_2 _48665_ (.A(_16449_),
    .B(_16712_),
    .Y(_16713_));
 sky130_as_sc_hs__or2_2 _48666_ (.A(\tholin_riscv.intr_vec[26] ),
    .B(_20005_),
    .Y(_16714_));
 sky130_as_sc_hs__nand3_2 _48667_ (.A(net137),
    .B(_16713_),
    .C(_16714_),
    .Y(_16715_));
 sky130_as_sc_hs__and2_2 _48668_ (.A(_16701_),
    .B(_16715_),
    .Y(_16716_));
 sky130_as_sc_hs__or2_2 _48669_ (.A(_16445_),
    .B(_16716_),
    .Y(_16717_));
 sky130_as_sc_hs__and2_2 _48672_ (.A(net503),
    .B(_16719_),
    .Y(_01245_));
 sky130_as_sc_hs__or2_2 _48674_ (.A(net7),
    .B(_19751_),
    .Y(_16721_));
 sky130_as_sc_hs__nand3_2 _48675_ (.A(_19759_),
    .B(_16720_),
    .C(_16721_),
    .Y(_16722_));
 sky130_as_sc_hs__nand3_2 _48679_ (.A(_16723_),
    .B(_16724_),
    .C(_16725_),
    .Y(_16726_));
 sky130_as_sc_hs__and2_2 _48682_ (.A(_16727_),
    .B(_16728_),
    .Y(_16729_));
 sky130_as_sc_hs__nand3_2 _48685_ (.A(_16729_),
    .B(_16730_),
    .C(_16731_),
    .Y(_16732_));
 sky130_as_sc_hs__nor2_2 _48686_ (.A(_16726_),
    .B(_16732_),
    .Y(_16733_));
 sky130_as_sc_hs__and2_2 _48690_ (.A(_16722_),
    .B(_16736_),
    .Y(_16737_));
 sky130_as_sc_hs__or2_2 _48691_ (.A(_16445_),
    .B(_16737_),
    .Y(_16738_));
 sky130_as_sc_hs__and2_2 _48694_ (.A(net493),
    .B(_16740_),
    .Y(_01246_));
 sky130_as_sc_hs__or2_2 _48695_ (.A(_19750_),
    .B(_02381_),
    .Y(_16741_));
 sky130_as_sc_hs__or2_2 _48696_ (.A(net8),
    .B(_19751_),
    .Y(_16742_));
 sky130_as_sc_hs__nand3_2 _48697_ (.A(_19759_),
    .B(_16741_),
    .C(_16742_),
    .Y(_16743_));
 sky130_as_sc_hs__nand3_2 _48701_ (.A(_16744_),
    .B(_16745_),
    .C(_16746_),
    .Y(_16747_));
 sky130_as_sc_hs__and2_2 _48704_ (.A(_16748_),
    .B(_16749_),
    .Y(_16750_));
 sky130_as_sc_hs__nand3_2 _48707_ (.A(_16750_),
    .B(_16751_),
    .C(_16752_),
    .Y(_16753_));
 sky130_as_sc_hs__or2_2 _48708_ (.A(_16747_),
    .B(_16753_),
    .Y(_16754_));
 sky130_as_sc_hs__or2_2 _48709_ (.A(_16449_),
    .B(_16754_),
    .Y(_16755_));
 sky130_as_sc_hs__or2_2 _48710_ (.A(\tholin_riscv.intr_vec[28] ),
    .B(_20005_),
    .Y(_16756_));
 sky130_as_sc_hs__nand3_2 _48711_ (.A(net137),
    .B(_16755_),
    .C(_16756_),
    .Y(_16757_));
 sky130_as_sc_hs__and2_2 _48712_ (.A(_16743_),
    .B(_16757_),
    .Y(_16758_));
 sky130_as_sc_hs__or2_2 _48713_ (.A(_16445_),
    .B(_16758_),
    .Y(_16759_));
 sky130_as_sc_hs__and2_2 _48716_ (.A(net493),
    .B(_16761_),
    .Y(_01247_));
 sky130_as_sc_hs__or2_2 _48717_ (.A(_19750_),
    .B(_23598_),
    .Y(_16762_));
 sky130_as_sc_hs__or2_2 _48718_ (.A(net9),
    .B(_19751_),
    .Y(_16763_));
 sky130_as_sc_hs__nand3_2 _48719_ (.A(_19759_),
    .B(_16762_),
    .C(_16763_),
    .Y(_16764_));
 sky130_as_sc_hs__nand3_2 _48723_ (.A(_16765_),
    .B(_16766_),
    .C(_16767_),
    .Y(_16768_));
 sky130_as_sc_hs__and2_2 _48726_ (.A(_16769_),
    .B(_16770_),
    .Y(_16771_));
 sky130_as_sc_hs__nand3_2 _48729_ (.A(_16771_),
    .B(_16772_),
    .C(_16773_),
    .Y(_16774_));
 sky130_as_sc_hs__nor2_2 _48730_ (.A(_16768_),
    .B(_16774_),
    .Y(_16775_));
 sky130_as_sc_hs__and2_2 _48734_ (.A(_16764_),
    .B(_16778_),
    .Y(_16779_));
 sky130_as_sc_hs__or2_2 _48735_ (.A(_16445_),
    .B(_16779_),
    .Y(_16780_));
 sky130_as_sc_hs__and2_2 _48738_ (.A(net517),
    .B(_16782_),
    .Y(_01248_));
 sky130_as_sc_hs__and2_2 _48741_ (.A(net493),
    .B(_16784_),
    .Y(_01249_));
 sky130_as_sc_hs__or2_2 _48742_ (.A(_19936_),
    .B(_06155_),
    .Y(_16785_));
 sky130_as_sc_hs__or2_2 _48743_ (.A(\tholin_riscv.PC[0] ),
    .B(_19937_),
    .Y(_16786_));
 sky130_as_sc_hs__or2_2 _48746_ (.A(net1691),
    .B(_16428_),
    .Y(_16789_));
 sky130_as_sc_hs__and2_2 _48747_ (.A(net500),
    .B(_16789_),
    .Y(_16790_));
 sky130_as_sc_hs__and2_2 _48748_ (.A(_16788_),
    .B(_16790_),
    .Y(_01250_));
 sky130_as_sc_hs__or2_2 _48750_ (.A(\tholin_riscv.PC[1] ),
    .B(_19937_),
    .Y(_16792_));
 sky130_as_sc_hs__or2_2 _48753_ (.A(net1595),
    .B(_16428_),
    .Y(_16795_));
 sky130_as_sc_hs__and2_2 _48754_ (.A(net494),
    .B(net1596),
    .Y(_16796_));
 sky130_as_sc_hs__and2_2 _48755_ (.A(_16794_),
    .B(_16796_),
    .Y(_01251_));
 sky130_as_sc_hs__and2_2 _48761_ (.A(net490),
    .B(_16801_),
    .Y(_16802_));
 sky130_as_sc_hs__and2_2 _48762_ (.A(_16800_),
    .B(_16802_),
    .Y(_01252_));
 sky130_as_sc_hs__or2_2 _48764_ (.A(\tholin_riscv.PC[3] ),
    .B(_19937_),
    .Y(_16804_));
 sky130_as_sc_hs__and2_2 _48768_ (.A(net490),
    .B(_16807_),
    .Y(_16808_));
 sky130_as_sc_hs__and2_2 _48769_ (.A(_16806_),
    .B(_16808_),
    .Y(_01253_));
 sky130_as_sc_hs__or2_2 _48771_ (.A(\tholin_riscv.PC[4] ),
    .B(_19937_),
    .Y(_16810_));
 sky130_as_sc_hs__and2_2 _48775_ (.A(net490),
    .B(_16813_),
    .Y(_16814_));
 sky130_as_sc_hs__and2_2 _48776_ (.A(_16812_),
    .B(_16814_),
    .Y(_01254_));
 sky130_as_sc_hs__or2_2 _48778_ (.A(\tholin_riscv.PC[5] ),
    .B(_19937_),
    .Y(_16816_));
 sky130_as_sc_hs__and2_2 _48782_ (.A(net490),
    .B(_16819_),
    .Y(_16820_));
 sky130_as_sc_hs__and2_2 _48783_ (.A(_16818_),
    .B(_16820_),
    .Y(_01255_));
 sky130_as_sc_hs__or2_2 _48785_ (.A(\tholin_riscv.PC[6] ),
    .B(_19937_),
    .Y(_16822_));
 sky130_as_sc_hs__or2_2 _48788_ (.A(net1703),
    .B(net131),
    .Y(_16825_));
 sky130_as_sc_hs__and2_2 _48789_ (.A(net490),
    .B(_16825_),
    .Y(_16826_));
 sky130_as_sc_hs__and2_2 _48790_ (.A(_16824_),
    .B(_16826_),
    .Y(_01256_));
 sky130_as_sc_hs__or2_2 _48792_ (.A(\tholin_riscv.PC[7] ),
    .B(_19937_),
    .Y(_16828_));
 sky130_as_sc_hs__and2_2 _48796_ (.A(net490),
    .B(_16831_),
    .Y(_16832_));
 sky130_as_sc_hs__and2_2 _48797_ (.A(_16830_),
    .B(_16832_),
    .Y(_01257_));
 sky130_as_sc_hs__or2_2 _48799_ (.A(\tholin_riscv.PC[8] ),
    .B(_19937_),
    .Y(_16834_));
 sky130_as_sc_hs__or2_2 _48802_ (.A(net1638),
    .B(net130),
    .Y(_16837_));
 sky130_as_sc_hs__and2_2 _48803_ (.A(net488),
    .B(net1639),
    .Y(_16838_));
 sky130_as_sc_hs__and2_2 _48804_ (.A(_16836_),
    .B(_16838_),
    .Y(_01258_));
 sky130_as_sc_hs__or2_2 _48806_ (.A(\tholin_riscv.PC[9] ),
    .B(_19937_),
    .Y(_16840_));
 sky130_as_sc_hs__or2_2 _48809_ (.A(net1612),
    .B(net130),
    .Y(_16843_));
 sky130_as_sc_hs__and2_2 _48810_ (.A(net488),
    .B(net1613),
    .Y(_16844_));
 sky130_as_sc_hs__and2_2 _48811_ (.A(_16842_),
    .B(_16844_),
    .Y(_01259_));
 sky130_as_sc_hs__or2_2 _48813_ (.A(\tholin_riscv.PC[10] ),
    .B(_19937_),
    .Y(_16846_));
 sky130_as_sc_hs__or2_2 _48816_ (.A(net1565),
    .B(net130),
    .Y(_16849_));
 sky130_as_sc_hs__and2_2 _48817_ (.A(net488),
    .B(net1566),
    .Y(_16850_));
 sky130_as_sc_hs__and2_2 _48818_ (.A(_16848_),
    .B(net1567),
    .Y(_01260_));
 sky130_as_sc_hs__or2_2 _48820_ (.A(\tholin_riscv.PC[11] ),
    .B(_19937_),
    .Y(_16852_));
 sky130_as_sc_hs__or2_2 _48823_ (.A(net1398),
    .B(net130),
    .Y(_16855_));
 sky130_as_sc_hs__and2_2 _48824_ (.A(net488),
    .B(net1399),
    .Y(_16856_));
 sky130_as_sc_hs__and2_2 _48825_ (.A(_16854_),
    .B(net1400),
    .Y(_01261_));
 sky130_as_sc_hs__or2_2 _48827_ (.A(\tholin_riscv.PC[12] ),
    .B(_19937_),
    .Y(_16858_));
 sky130_as_sc_hs__or2_2 _48830_ (.A(net1610),
    .B(net130),
    .Y(_16861_));
 sky130_as_sc_hs__and2_2 _48831_ (.A(net490),
    .B(net1611),
    .Y(_16862_));
 sky130_as_sc_hs__and2_2 _48832_ (.A(_16860_),
    .B(_16862_),
    .Y(_01262_));
 sky130_as_sc_hs__or2_2 _48834_ (.A(\tholin_riscv.PC[13] ),
    .B(_19937_),
    .Y(_16864_));
 sky130_as_sc_hs__or2_2 _48837_ (.A(net1618),
    .B(net130),
    .Y(_16867_));
 sky130_as_sc_hs__and2_2 _48838_ (.A(net488),
    .B(net1619),
    .Y(_16868_));
 sky130_as_sc_hs__and2_2 _48839_ (.A(_16866_),
    .B(_16868_),
    .Y(_01263_));
 sky130_as_sc_hs__or2_2 _48841_ (.A(\tholin_riscv.PC[14] ),
    .B(_19937_),
    .Y(_16870_));
 sky130_as_sc_hs__or2_2 _48844_ (.A(net1483),
    .B(net131),
    .Y(_16873_));
 sky130_as_sc_hs__and2_2 _48845_ (.A(net490),
    .B(net1484),
    .Y(_16874_));
 sky130_as_sc_hs__and2_2 _48846_ (.A(_16872_),
    .B(net1485),
    .Y(_01264_));
 sky130_as_sc_hs__or2_2 _48848_ (.A(\tholin_riscv.PC[15] ),
    .B(_19937_),
    .Y(_16876_));
 sky130_as_sc_hs__or2_2 _48851_ (.A(net1590),
    .B(net131),
    .Y(_16879_));
 sky130_as_sc_hs__and2_2 _48852_ (.A(net490),
    .B(net1591),
    .Y(_16880_));
 sky130_as_sc_hs__and2_2 _48853_ (.A(_16878_),
    .B(net1592),
    .Y(_01265_));
 sky130_as_sc_hs__or2_2 _48855_ (.A(\tholin_riscv.PC[16] ),
    .B(_19937_),
    .Y(_16882_));
 sky130_as_sc_hs__or2_2 _48858_ (.A(net1598),
    .B(net131),
    .Y(_16885_));
 sky130_as_sc_hs__and2_2 _48859_ (.A(net490),
    .B(net1599),
    .Y(_16886_));
 sky130_as_sc_hs__and2_2 _48860_ (.A(_16884_),
    .B(_16886_),
    .Y(_01266_));
 sky130_as_sc_hs__or2_2 _48862_ (.A(\tholin_riscv.PC[17] ),
    .B(_19937_),
    .Y(_16888_));
 sky130_as_sc_hs__or2_2 _48865_ (.A(net1632),
    .B(net131),
    .Y(_16891_));
 sky130_as_sc_hs__and2_2 _48866_ (.A(net491),
    .B(net1633),
    .Y(_16892_));
 sky130_as_sc_hs__and2_2 _48867_ (.A(_16890_),
    .B(_16892_),
    .Y(_01267_));
 sky130_as_sc_hs__or2_2 _48869_ (.A(\tholin_riscv.PC[18] ),
    .B(_19937_),
    .Y(_16894_));
 sky130_as_sc_hs__or2_2 _48872_ (.A(net1401),
    .B(net131),
    .Y(_16897_));
 sky130_as_sc_hs__and2_2 _48873_ (.A(net491),
    .B(net1402),
    .Y(_16898_));
 sky130_as_sc_hs__and2_2 _48874_ (.A(_16896_),
    .B(net1403),
    .Y(_01268_));
 sky130_as_sc_hs__or2_2 _48876_ (.A(\tholin_riscv.PC[19] ),
    .B(_19937_),
    .Y(_16900_));
 sky130_as_sc_hs__or2_2 _48879_ (.A(net1574),
    .B(net131),
    .Y(_16903_));
 sky130_as_sc_hs__and2_2 _48880_ (.A(net491),
    .B(net1575),
    .Y(_16904_));
 sky130_as_sc_hs__and2_2 _48881_ (.A(_16902_),
    .B(net1576),
    .Y(_01269_));
 sky130_as_sc_hs__or2_2 _48883_ (.A(\tholin_riscv.PC[20] ),
    .B(_19937_),
    .Y(_16906_));
 sky130_as_sc_hs__or2_2 _48886_ (.A(net1616),
    .B(net130),
    .Y(_16909_));
 sky130_as_sc_hs__and2_2 _48887_ (.A(net488),
    .B(net1617),
    .Y(_16910_));
 sky130_as_sc_hs__and2_2 _48888_ (.A(_16908_),
    .B(_16910_),
    .Y(_01270_));
 sky130_as_sc_hs__or2_2 _48890_ (.A(\tholin_riscv.PC[21] ),
    .B(_19937_),
    .Y(_16912_));
 sky130_as_sc_hs__or2_2 _48893_ (.A(net1603),
    .B(net130),
    .Y(_16915_));
 sky130_as_sc_hs__and2_2 _48894_ (.A(net489),
    .B(net1604),
    .Y(_16916_));
 sky130_as_sc_hs__and2_2 _48895_ (.A(_16914_),
    .B(_16916_),
    .Y(_01271_));
 sky130_as_sc_hs__or2_2 _48897_ (.A(\tholin_riscv.PC[22] ),
    .B(_19937_),
    .Y(_16918_));
 sky130_as_sc_hs__or2_2 _48900_ (.A(net1518),
    .B(net131),
    .Y(_16921_));
 sky130_as_sc_hs__and2_2 _48901_ (.A(net489),
    .B(net1519),
    .Y(_16922_));
 sky130_as_sc_hs__and2_2 _48902_ (.A(_16920_),
    .B(net1520),
    .Y(_01272_));
 sky130_as_sc_hs__or2_2 _48904_ (.A(\tholin_riscv.PC[23] ),
    .B(_19937_),
    .Y(_16924_));
 sky130_as_sc_hs__or2_2 _48907_ (.A(net1512),
    .B(net131),
    .Y(_16927_));
 sky130_as_sc_hs__and2_2 _48908_ (.A(net489),
    .B(net1513),
    .Y(_16928_));
 sky130_as_sc_hs__and2_2 _48909_ (.A(_16926_),
    .B(net1514),
    .Y(_01273_));
 sky130_as_sc_hs__or2_2 _48911_ (.A(\tholin_riscv.PC[24] ),
    .B(_19937_),
    .Y(_16930_));
 sky130_as_sc_hs__or2_2 _48914_ (.A(net1605),
    .B(net130),
    .Y(_16933_));
 sky130_as_sc_hs__and2_2 _48915_ (.A(net488),
    .B(net1606),
    .Y(_16934_));
 sky130_as_sc_hs__and2_2 _48916_ (.A(_16932_),
    .B(_16934_),
    .Y(_01274_));
 sky130_as_sc_hs__or2_2 _48918_ (.A(\tholin_riscv.PC[25] ),
    .B(_19937_),
    .Y(_16936_));
 sky130_as_sc_hs__or2_2 _48921_ (.A(net1600),
    .B(net130),
    .Y(_16939_));
 sky130_as_sc_hs__and2_2 _48922_ (.A(net488),
    .B(net1601),
    .Y(_16940_));
 sky130_as_sc_hs__and2_2 _48923_ (.A(_16938_),
    .B(_16940_),
    .Y(_01275_));
 sky130_as_sc_hs__or2_2 _48925_ (.A(\tholin_riscv.PC[26] ),
    .B(_19937_),
    .Y(_16942_));
 sky130_as_sc_hs__or2_2 _48928_ (.A(net1562),
    .B(net130),
    .Y(_16945_));
 sky130_as_sc_hs__and2_2 _48929_ (.A(net488),
    .B(net1563),
    .Y(_16946_));
 sky130_as_sc_hs__and2_2 _48930_ (.A(_16944_),
    .B(net1564),
    .Y(_01276_));
 sky130_as_sc_hs__or2_2 _48932_ (.A(\tholin_riscv.PC[27] ),
    .B(_19937_),
    .Y(_16948_));
 sky130_as_sc_hs__or2_2 _48935_ (.A(net1386),
    .B(net130),
    .Y(_16951_));
 sky130_as_sc_hs__and2_2 _48936_ (.A(net488),
    .B(net1387),
    .Y(_16952_));
 sky130_as_sc_hs__and2_2 _48937_ (.A(_16950_),
    .B(net1388),
    .Y(_01277_));
 sky130_as_sc_hs__or2_2 _48939_ (.A(\tholin_riscv.PC[28] ),
    .B(_19937_),
    .Y(_16954_));
 sky130_as_sc_hs__or2_2 _48942_ (.A(net1622),
    .B(net130),
    .Y(_16957_));
 sky130_as_sc_hs__and2_2 _48943_ (.A(net489),
    .B(net1623),
    .Y(_16958_));
 sky130_as_sc_hs__and2_2 _48944_ (.A(_16956_),
    .B(_16958_),
    .Y(_01278_));
 sky130_as_sc_hs__or2_2 _48946_ (.A(\tholin_riscv.PC[29] ),
    .B(_19937_),
    .Y(_16960_));
 sky130_as_sc_hs__or2_2 _48949_ (.A(net1614),
    .B(net130),
    .Y(_16963_));
 sky130_as_sc_hs__and2_2 _48950_ (.A(net488),
    .B(net1615),
    .Y(_16964_));
 sky130_as_sc_hs__and2_2 _48951_ (.A(_16962_),
    .B(_16964_),
    .Y(_01279_));
 sky130_as_sc_hs__or2_2 _48952_ (.A(_19936_),
    .B(_12575_),
    .Y(_16965_));
 sky130_as_sc_hs__or2_2 _48953_ (.A(\tholin_riscv.PC[30] ),
    .B(_19937_),
    .Y(_16966_));
 sky130_as_sc_hs__or2_2 _48956_ (.A(net1571),
    .B(net130),
    .Y(_16969_));
 sky130_as_sc_hs__and2_2 _48957_ (.A(net489),
    .B(net1572),
    .Y(_16970_));
 sky130_as_sc_hs__and2_2 _48958_ (.A(_16968_),
    .B(net1573),
    .Y(_01280_));
 sky130_as_sc_hs__or2_2 _48960_ (.A(\tholin_riscv.PC[31] ),
    .B(_19937_),
    .Y(_16972_));
 sky130_as_sc_hs__or2_2 _48963_ (.A(net1358),
    .B(net130),
    .Y(_16975_));
 sky130_as_sc_hs__and2_2 _48964_ (.A(net488),
    .B(net1359),
    .Y(_16976_));
 sky130_as_sc_hs__and2_2 _48965_ (.A(_16974_),
    .B(net1360),
    .Y(_01281_));
 sky130_as_sc_hs__or2_2 _48966_ (.A(net1316),
    .B(net105),
    .Y(_16977_));
 sky130_as_sc_hs__and2_2 _48968_ (.A(net484),
    .B(net1317),
    .Y(_16979_));
 sky130_as_sc_hs__and2_2 _48969_ (.A(_16978_),
    .B(net1318),
    .Y(_01282_));
 sky130_as_sc_hs__or2_2 _48970_ (.A(net1220),
    .B(net105),
    .Y(_16980_));
 sky130_as_sc_hs__and2_2 _48972_ (.A(net484),
    .B(net1221),
    .Y(_16982_));
 sky130_as_sc_hs__and2_2 _48973_ (.A(_16981_),
    .B(net1222),
    .Y(_01283_));
 sky130_as_sc_hs__or2_2 _48974_ (.A(net1217),
    .B(net105),
    .Y(_16983_));
 sky130_as_sc_hs__and2_2 _48976_ (.A(net485),
    .B(net1218),
    .Y(_16985_));
 sky130_as_sc_hs__and2_2 _48977_ (.A(_16984_),
    .B(net1219),
    .Y(_01284_));
 sky130_as_sc_hs__or2_2 _48978_ (.A(net1141),
    .B(net105),
    .Y(_16986_));
 sky130_as_sc_hs__and2_2 _48980_ (.A(net484),
    .B(net1142),
    .Y(_16988_));
 sky130_as_sc_hs__and2_2 _48981_ (.A(_16987_),
    .B(net1143),
    .Y(_01285_));
 sky130_as_sc_hs__or2_2 _48982_ (.A(net1295),
    .B(net105),
    .Y(_16989_));
 sky130_as_sc_hs__and2_2 _48984_ (.A(net484),
    .B(net1296),
    .Y(_16991_));
 sky130_as_sc_hs__and2_2 _48985_ (.A(_16990_),
    .B(net1297),
    .Y(_01286_));
 sky130_as_sc_hs__or2_2 _48986_ (.A(net1266),
    .B(net106),
    .Y(_16992_));
 sky130_as_sc_hs__or2_2 _48987_ (.A(\tholin_riscv.Bimm[11] ),
    .B(_19931_),
    .Y(_16993_));
 sky130_as_sc_hs__and2_2 _48988_ (.A(net491),
    .B(net1267),
    .Y(_16994_));
 sky130_as_sc_hs__and2_2 _48989_ (.A(_16993_),
    .B(net1268),
    .Y(_01287_));
 sky130_as_sc_hs__or2_2 _48990_ (.A(net1277),
    .B(net106),
    .Y(_16995_));
 sky130_as_sc_hs__or2_2 _48991_ (.A(net1260),
    .B(_19931_),
    .Y(_16996_));
 sky130_as_sc_hs__and2_2 _48992_ (.A(net493),
    .B(net1278),
    .Y(_16997_));
 sky130_as_sc_hs__and2_2 _48993_ (.A(_16996_),
    .B(net1279),
    .Y(_01288_));
 sky130_as_sc_hs__or2_2 _48994_ (.A(net1147),
    .B(net106),
    .Y(_16998_));
 sky130_as_sc_hs__or2_2 _48995_ (.A(net1780),
    .B(_19931_),
    .Y(_16999_));
 sky130_as_sc_hs__and2_2 _48996_ (.A(net493),
    .B(net1148),
    .Y(_17000_));
 sky130_as_sc_hs__and2_2 _48997_ (.A(_16999_),
    .B(net1149),
    .Y(_01289_));
 sky130_as_sc_hs__or2_2 _48998_ (.A(net1241),
    .B(net106),
    .Y(_17001_));
 sky130_as_sc_hs__or2_2 _48999_ (.A(net1791),
    .B(_19931_),
    .Y(_17002_));
 sky130_as_sc_hs__and2_2 _49000_ (.A(net493),
    .B(net1242),
    .Y(_17003_));
 sky130_as_sc_hs__and2_2 _49001_ (.A(_17002_),
    .B(net1243),
    .Y(_01290_));
 sky130_as_sc_hs__or2_2 _49002_ (.A(net1270),
    .B(net106),
    .Y(_17004_));
 sky130_as_sc_hs__or2_2 _49003_ (.A(net1792),
    .B(_19931_),
    .Y(_17005_));
 sky130_as_sc_hs__and2_2 _49004_ (.A(net493),
    .B(net1271),
    .Y(_17006_));
 sky130_as_sc_hs__and2_2 _49005_ (.A(_17005_),
    .B(net1272),
    .Y(_01291_));
 sky130_as_sc_hs__or2_2 _49006_ (.A(net1263),
    .B(net105),
    .Y(_17007_));
 sky130_as_sc_hs__and2_2 _49008_ (.A(net484),
    .B(net1264),
    .Y(_17009_));
 sky130_as_sc_hs__and2_2 _49009_ (.A(_17008_),
    .B(net1265),
    .Y(_01292_));
 sky130_as_sc_hs__or2_2 _49010_ (.A(net1245),
    .B(net105),
    .Y(_17010_));
 sky130_as_sc_hs__and2_2 _49012_ (.A(net485),
    .B(net1246),
    .Y(_17012_));
 sky130_as_sc_hs__and2_2 _49013_ (.A(_17011_),
    .B(net1247),
    .Y(_01293_));
 sky130_as_sc_hs__or2_2 _49014_ (.A(net1120),
    .B(net106),
    .Y(_17013_));
 sky130_as_sc_hs__or2_2 _49015_ (.A(net411),
    .B(_19931_),
    .Y(_17014_));
 sky130_as_sc_hs__and2_2 _49016_ (.A(net493),
    .B(net1121),
    .Y(_17015_));
 sky130_as_sc_hs__and2_2 _49017_ (.A(_17014_),
    .B(net1122),
    .Y(_01294_));
 sky130_as_sc_hs__or2_2 _49018_ (.A(net1106),
    .B(net105),
    .Y(_17016_));
 sky130_as_sc_hs__and2_2 _49020_ (.A(net485),
    .B(net1107),
    .Y(_17018_));
 sky130_as_sc_hs__and2_2 _49021_ (.A(_17017_),
    .B(net1108),
    .Y(_01295_));
 sky130_as_sc_hs__or2_2 _49022_ (.A(net1539),
    .B(net105),
    .Y(_17019_));
 sky130_as_sc_hs__and2_2 _49024_ (.A(net499),
    .B(net1540),
    .Y(_17021_));
 sky130_as_sc_hs__and2_2 _49025_ (.A(_17020_),
    .B(net1541),
    .Y(_01296_));
 sky130_as_sc_hs__or2_2 _49026_ (.A(net1337),
    .B(net105),
    .Y(_17022_));
 sky130_as_sc_hs__and2_2 _49028_ (.A(net484),
    .B(net1338),
    .Y(_17024_));
 sky130_as_sc_hs__and2_2 _49029_ (.A(_17023_),
    .B(net1339),
    .Y(_01297_));
 sky130_as_sc_hs__or2_2 _49030_ (.A(net1076),
    .B(net105),
    .Y(_17025_));
 sky130_as_sc_hs__and2_2 _49032_ (.A(net485),
    .B(net1077),
    .Y(_17027_));
 sky130_as_sc_hs__and2_2 _49033_ (.A(_17026_),
    .B(net1078),
    .Y(_01298_));
 sky130_as_sc_hs__or2_2 _49034_ (.A(net1548),
    .B(net106),
    .Y(_17028_));
 sky130_as_sc_hs__and2_2 _49036_ (.A(net499),
    .B(net1549),
    .Y(_17030_));
 sky130_as_sc_hs__and2_2 _49037_ (.A(_17029_),
    .B(net1550),
    .Y(_01299_));
 sky130_as_sc_hs__or2_2 _49038_ (.A(net1086),
    .B(net106),
    .Y(_17031_));
 sky130_as_sc_hs__or2_2 _49039_ (.A(\tholin_riscv.Iimm[0] ),
    .B(_19931_),
    .Y(_17032_));
 sky130_as_sc_hs__and2_2 _49040_ (.A(net491),
    .B(net1087),
    .Y(_17033_));
 sky130_as_sc_hs__and2_2 _49041_ (.A(_17032_),
    .B(net1088),
    .Y(_01300_));
 sky130_as_sc_hs__or2_2 _49042_ (.A(net1144),
    .B(net105),
    .Y(_17034_));
 sky130_as_sc_hs__and2_2 _49044_ (.A(net484),
    .B(net1145),
    .Y(_17036_));
 sky130_as_sc_hs__and2_2 _49045_ (.A(_17035_),
    .B(net1146),
    .Y(_01301_));
 sky130_as_sc_hs__or2_2 _49046_ (.A(net1524),
    .B(net105),
    .Y(_17037_));
 sky130_as_sc_hs__or2_2 _49047_ (.A(\tholin_riscv.Iimm[2] ),
    .B(_19931_),
    .Y(_17038_));
 sky130_as_sc_hs__and2_2 _49048_ (.A(net497),
    .B(net1525),
    .Y(_17039_));
 sky130_as_sc_hs__and2_2 _49049_ (.A(_17038_),
    .B(_17039_),
    .Y(_01302_));
 sky130_as_sc_hs__or2_2 _49050_ (.A(net1113),
    .B(net105),
    .Y(_17040_));
 sky130_as_sc_hs__and2_2 _49052_ (.A(net485),
    .B(net1114),
    .Y(_17042_));
 sky130_as_sc_hs__and2_2 _49053_ (.A(_17041_),
    .B(net1115),
    .Y(_01303_));
 sky130_as_sc_hs__or2_2 _49054_ (.A(net1195),
    .B(net105),
    .Y(_17043_));
 sky130_as_sc_hs__and2_2 _49056_ (.A(net484),
    .B(net1196),
    .Y(_17045_));
 sky130_as_sc_hs__and2_2 _49057_ (.A(_17044_),
    .B(net1197),
    .Y(_01304_));
 sky130_as_sc_hs__or2_2 _49058_ (.A(net1408),
    .B(net106),
    .Y(_17046_));
 sky130_as_sc_hs__or2_2 _49059_ (.A(\tholin_riscv.Bimm[5] ),
    .B(_19931_),
    .Y(_17047_));
 sky130_as_sc_hs__and2_2 _49060_ (.A(net497),
    .B(net1409),
    .Y(_17048_));
 sky130_as_sc_hs__and2_2 _49061_ (.A(_17047_),
    .B(net1410),
    .Y(_01305_));
 sky130_as_sc_hs__or2_2 _49062_ (.A(net1151),
    .B(net106),
    .Y(_17049_));
 sky130_as_sc_hs__or2_2 _49063_ (.A(\tholin_riscv.Bimm[6] ),
    .B(_19931_),
    .Y(_17050_));
 sky130_as_sc_hs__and2_2 _49064_ (.A(net493),
    .B(net1152),
    .Y(_17051_));
 sky130_as_sc_hs__and2_2 _49065_ (.A(_17050_),
    .B(net1153),
    .Y(_01306_));
 sky130_as_sc_hs__or2_2 _49066_ (.A(net1182),
    .B(net105),
    .Y(_17052_));
 sky130_as_sc_hs__and2_2 _49068_ (.A(net484),
    .B(net1183),
    .Y(_17054_));
 sky130_as_sc_hs__and2_2 _49069_ (.A(_17053_),
    .B(net1184),
    .Y(_01307_));
 sky130_as_sc_hs__or2_2 _49070_ (.A(net1593),
    .B(net106),
    .Y(_17055_));
 sky130_as_sc_hs__and2_2 _49072_ (.A(net499),
    .B(net1594),
    .Y(_17057_));
 sky130_as_sc_hs__and2_2 _49073_ (.A(_17056_),
    .B(_17057_),
    .Y(_01308_));
 sky130_as_sc_hs__or2_2 _49074_ (.A(net1229),
    .B(net106),
    .Y(_17058_));
 sky130_as_sc_hs__or2_2 _49075_ (.A(net1832),
    .B(_19931_),
    .Y(_17059_));
 sky130_as_sc_hs__and2_2 _49076_ (.A(net495),
    .B(net1230),
    .Y(_17060_));
 sky130_as_sc_hs__and2_2 _49077_ (.A(_17059_),
    .B(net1231),
    .Y(_01309_));
 sky130_as_sc_hs__or2_2 _49078_ (.A(net1425),
    .B(net106),
    .Y(_17061_));
 sky130_as_sc_hs__or2_2 _49079_ (.A(\tholin_riscv.Bimm[10] ),
    .B(_19931_),
    .Y(_17062_));
 sky130_as_sc_hs__and2_2 _49080_ (.A(net497),
    .B(net1426),
    .Y(_17063_));
 sky130_as_sc_hs__and2_2 _49081_ (.A(_17062_),
    .B(net1427),
    .Y(_01310_));
 sky130_as_sc_hs__or2_2 _49082_ (.A(net1116),
    .B(net106),
    .Y(_17064_));
 sky130_as_sc_hs__or2_2 _49083_ (.A(\tholin_riscv.Bimm[12] ),
    .B(_19931_),
    .Y(_17065_));
 sky130_as_sc_hs__and2_2 _49084_ (.A(net493),
    .B(net1117),
    .Y(_17066_));
 sky130_as_sc_hs__and2_2 _49085_ (.A(_17065_),
    .B(net1118),
    .Y(_01311_));
 sky130_as_sc_hs__and2_2 _49086_ (.A(net544),
    .B(net747),
    .Y(_17067_));
 sky130_as_sc_hs__and2_2 _49087_ (.A(net884),
    .B(_17067_),
    .Y(_17068_));
 sky130_as_sc_hs__and2_2 _49088_ (.A(net963),
    .B(_17068_),
    .Y(_17069_));
 sky130_as_sc_hs__and2_2 _49089_ (.A(net984),
    .B(_17069_),
    .Y(_17070_));
 sky130_as_sc_hs__and2_2 _49090_ (.A(_17070_),
    .B(net880),
    .Y(_17071_));
 sky130_as_sc_hs__and2_2 _49091_ (.A(_17071_),
    .B(net1109),
    .Y(_17072_));
 sky130_as_sc_hs__and2_2 _49092_ (.A(net927),
    .B(_17072_),
    .Y(_17073_));
 sky130_as_sc_hs__and2_2 _49093_ (.A(net1004),
    .B(_17073_),
    .Y(_17074_));
 sky130_as_sc_hs__and2_2 _49094_ (.A(net1008),
    .B(_17074_),
    .Y(_17075_));
 sky130_as_sc_hs__and2_2 _49095_ (.A(net980),
    .B(_17075_),
    .Y(_17076_));
 sky130_as_sc_hs__and2_2 _49096_ (.A(net976),
    .B(_17076_),
    .Y(_17077_));
 sky130_as_sc_hs__and2_2 _49097_ (.A(net1028),
    .B(_17077_),
    .Y(_17078_));
 sky130_as_sc_hs__and2_2 _49098_ (.A(net919),
    .B(_17078_),
    .Y(_17079_));
 sky130_as_sc_hs__and2_2 _49099_ (.A(net996),
    .B(_17079_),
    .Y(_17080_));
 sky130_as_sc_hs__and2_2 _49100_ (.A(net1065),
    .B(_17080_),
    .Y(_17081_));
 sky130_as_sc_hs__and2_2 _49101_ (.A(net1053),
    .B(_17081_),
    .Y(_17082_));
 sky130_as_sc_hs__and2_2 _49102_ (.A(net935),
    .B(_17082_),
    .Y(_17083_));
 sky130_as_sc_hs__and2_2 _49103_ (.A(net899),
    .B(_17083_),
    .Y(_17084_));
 sky130_as_sc_hs__and2_2 _49104_ (.A(_17084_),
    .B(net1038),
    .Y(_17085_));
 sky130_as_sc_hs__and2_2 _49105_ (.A(net911),
    .B(_17085_),
    .Y(_17086_));
 sky130_as_sc_hs__and2_2 _49106_ (.A(net891),
    .B(_17086_),
    .Y(_17087_));
 sky130_as_sc_hs__and2_2 _49107_ (.A(net931),
    .B(_17087_),
    .Y(_17088_));
 sky130_as_sc_hs__and2_2 _49108_ (.A(_17088_),
    .B(net1034),
    .Y(_17089_));
 sky130_as_sc_hs__and2_2 _49109_ (.A(net992),
    .B(_17089_),
    .Y(_17090_));
 sky130_as_sc_hs__and2_2 _49110_ (.A(_17090_),
    .B(net760),
    .Y(_17091_));
 sky130_as_sc_hs__and2_2 _49111_ (.A(net959),
    .B(_17091_),
    .Y(_17092_));
 sky130_as_sc_hs__and2_2 _49112_ (.A(net1057),
    .B(_17092_),
    .Y(_17093_));
 sky130_as_sc_hs__and2_2 _49113_ (.A(net1096),
    .B(_17093_),
    .Y(_17094_));
 sky130_as_sc_hs__and2_2 _49114_ (.A(_17094_),
    .B(net955),
    .Y(_17095_));
 sky130_as_sc_hs__and2_2 _49115_ (.A(net775),
    .B(_17095_),
    .Y(_17096_));
 sky130_as_sc_hs__or2_2 _49116_ (.A(\tholin_riscv.tmr0_pre_ctr[31] ),
    .B(_17096_),
    .Y(_17097_));
 sky130_as_sc_hs__nor2_2 _49120_ (.A(net911),
    .B(_17085_),
    .Y(_17101_));
 sky130_as_sc_hs__or2_2 _49121_ (.A(_17086_),
    .B(net912),
    .Y(_17102_));
 sky130_as_sc_hs__nor2_2 _49123_ (.A(net1038),
    .B(_17084_),
    .Y(_17104_));
 sky130_as_sc_hs__or2_2 _49124_ (.A(_17085_),
    .B(net1039),
    .Y(_17105_));
 sky130_as_sc_hs__or2_2 _49125_ (.A(\tholin_riscv.tmr0_pre[19] ),
    .B(_17105_),
    .Y(_17106_));
 sky130_as_sc_hs__nor2_2 _49126_ (.A(net996),
    .B(_17079_),
    .Y(_17107_));
 sky130_as_sc_hs__or2_2 _49127_ (.A(_17080_),
    .B(net997),
    .Y(_17108_));
 sky130_as_sc_hs__or2_2 _49128_ (.A(\tholin_riscv.tmr0_pre[14] ),
    .B(_17108_),
    .Y(_17109_));
 sky130_as_sc_hs__nor2_2 _49129_ (.A(net919),
    .B(_17078_),
    .Y(_17110_));
 sky130_as_sc_hs__or2_2 _49130_ (.A(_17079_),
    .B(net920),
    .Y(_17111_));
 sky130_as_sc_hs__nor2_2 _49132_ (.A(net1028),
    .B(_17077_),
    .Y(_17113_));
 sky130_as_sc_hs__or2_2 _49133_ (.A(_17078_),
    .B(net1029),
    .Y(_17114_));
 sky130_as_sc_hs__nor2_2 _49135_ (.A(net984),
    .B(_17069_),
    .Y(_17116_));
 sky130_as_sc_hs__or2_2 _49136_ (.A(_17070_),
    .B(net985),
    .Y(_17117_));
 sky130_as_sc_hs__or2_2 _49137_ (.A(\tholin_riscv.tmr0_pre[4] ),
    .B(_17117_),
    .Y(_17118_));
 sky130_as_sc_hs__nor2_2 _49138_ (.A(net963),
    .B(_17068_),
    .Y(_17119_));
 sky130_as_sc_hs__or2_2 _49139_ (.A(_17069_),
    .B(net964),
    .Y(_17120_));
 sky130_as_sc_hs__or2_2 _49140_ (.A(\tholin_riscv.tmr0_pre[3] ),
    .B(_17120_),
    .Y(_17121_));
 sky130_as_sc_hs__nor2_2 _49142_ (.A(net884),
    .B(_17067_),
    .Y(_17123_));
 sky130_as_sc_hs__or2_2 _49143_ (.A(_17068_),
    .B(net885),
    .Y(_17124_));
 sky130_as_sc_hs__or2_2 _49144_ (.A(\tholin_riscv.tmr0_pre[2] ),
    .B(_17124_),
    .Y(_17125_));
 sky130_as_sc_hs__nor2_2 _49146_ (.A(net544),
    .B(net747),
    .Y(_17127_));
 sky130_as_sc_hs__or2_2 _49147_ (.A(_17067_),
    .B(net748),
    .Y(_17128_));
 sky130_as_sc_hs__or2_2 _49148_ (.A(\tholin_riscv.tmr0_pre[1] ),
    .B(_17128_),
    .Y(_17129_));
 sky130_as_sc_hs__nand3_2 _49152_ (.A(_17125_),
    .B(_17129_),
    .C(_17132_),
    .Y(_17133_));
 sky130_as_sc_hs__nand3_2 _49153_ (.A(_17122_),
    .B(_17126_),
    .C(_17133_),
    .Y(_17134_));
 sky130_as_sc_hs__nand3_2 _49154_ (.A(_17118_),
    .B(_17121_),
    .C(_17134_),
    .Y(_17135_));
 sky130_as_sc_hs__nor2_2 _49155_ (.A(net880),
    .B(_17070_),
    .Y(_17136_));
 sky130_as_sc_hs__or2_2 _49156_ (.A(_17071_),
    .B(net881),
    .Y(_17137_));
 sky130_as_sc_hs__nand3_2 _49159_ (.A(_17135_),
    .B(_17138_),
    .C(_17139_),
    .Y(_17140_));
 sky130_as_sc_hs__or2_2 _49160_ (.A(\tholin_riscv.tmr0_pre[5] ),
    .B(_17137_),
    .Y(_17141_));
 sky130_as_sc_hs__nor2_2 _49161_ (.A(net1109),
    .B(_17071_),
    .Y(_17142_));
 sky130_as_sc_hs__or2_2 _49162_ (.A(_17072_),
    .B(net1110),
    .Y(_17143_));
 sky130_as_sc_hs__or2_2 _49163_ (.A(\tholin_riscv.tmr0_pre[6] ),
    .B(_17143_),
    .Y(_17144_));
 sky130_as_sc_hs__nand3_2 _49164_ (.A(_17140_),
    .B(_17141_),
    .C(_17144_),
    .Y(_17145_));
 sky130_as_sc_hs__nor2_2 _49166_ (.A(net927),
    .B(_17072_),
    .Y(_17147_));
 sky130_as_sc_hs__or2_2 _49167_ (.A(_17073_),
    .B(net928),
    .Y(_17148_));
 sky130_as_sc_hs__nand3_2 _49169_ (.A(_17145_),
    .B(_17146_),
    .C(_17149_),
    .Y(_17150_));
 sky130_as_sc_hs__or2_2 _49170_ (.A(\tholin_riscv.tmr0_pre[7] ),
    .B(_17148_),
    .Y(_17151_));
 sky130_as_sc_hs__nor2_2 _49171_ (.A(net1004),
    .B(_17073_),
    .Y(_17152_));
 sky130_as_sc_hs__or2_2 _49172_ (.A(_17074_),
    .B(net1005),
    .Y(_17153_));
 sky130_as_sc_hs__or2_2 _49173_ (.A(\tholin_riscv.tmr0_pre[8] ),
    .B(_17153_),
    .Y(_17154_));
 sky130_as_sc_hs__nand3_2 _49174_ (.A(_17150_),
    .B(_17151_),
    .C(_17154_),
    .Y(_17155_));
 sky130_as_sc_hs__nor2_2 _49176_ (.A(net1008),
    .B(_17074_),
    .Y(_17157_));
 sky130_as_sc_hs__or2_2 _49177_ (.A(_17075_),
    .B(net1009),
    .Y(_17158_));
 sky130_as_sc_hs__nand3_2 _49179_ (.A(_17155_),
    .B(_17156_),
    .C(_17159_),
    .Y(_17160_));
 sky130_as_sc_hs__or2_2 _49180_ (.A(\tholin_riscv.tmr0_pre[9] ),
    .B(_17158_),
    .Y(_17161_));
 sky130_as_sc_hs__nor2_2 _49181_ (.A(net980),
    .B(_17075_),
    .Y(_17162_));
 sky130_as_sc_hs__or2_2 _49182_ (.A(_17076_),
    .B(net981),
    .Y(_17163_));
 sky130_as_sc_hs__or2_2 _49183_ (.A(\tholin_riscv.tmr0_pre[10] ),
    .B(_17163_),
    .Y(_17164_));
 sky130_as_sc_hs__nand3_2 _49184_ (.A(_17160_),
    .B(_17161_),
    .C(_17164_),
    .Y(_17165_));
 sky130_as_sc_hs__nor2_2 _49186_ (.A(net976),
    .B(_17076_),
    .Y(_17167_));
 sky130_as_sc_hs__or2_2 _49187_ (.A(_17077_),
    .B(net977),
    .Y(_17168_));
 sky130_as_sc_hs__nand3_2 _49189_ (.A(_17165_),
    .B(_17166_),
    .C(_17169_),
    .Y(_17170_));
 sky130_as_sc_hs__or2_2 _49190_ (.A(\tholin_riscv.tmr0_pre[12] ),
    .B(_17114_),
    .Y(_17171_));
 sky130_as_sc_hs__or2_2 _49191_ (.A(\tholin_riscv.tmr0_pre[11] ),
    .B(_17168_),
    .Y(_17172_));
 sky130_as_sc_hs__nand3_2 _49192_ (.A(_17170_),
    .B(_17171_),
    .C(_17172_),
    .Y(_17173_));
 sky130_as_sc_hs__or2_2 _49194_ (.A(\tholin_riscv.tmr0_pre[13] ),
    .B(_17111_),
    .Y(_17175_));
 sky130_as_sc_hs__nor2_2 _49198_ (.A(net1065),
    .B(_17080_),
    .Y(_17179_));
 sky130_as_sc_hs__or2_2 _49199_ (.A(_17081_),
    .B(net1066),
    .Y(_17180_));
 sky130_as_sc_hs__nand3_2 _49202_ (.A(_17178_),
    .B(_17181_),
    .C(_17182_),
    .Y(_17183_));
 sky130_as_sc_hs__or2_2 _49203_ (.A(\tholin_riscv.tmr0_pre[15] ),
    .B(_17180_),
    .Y(_17184_));
 sky130_as_sc_hs__nor2_2 _49204_ (.A(net1053),
    .B(_17081_),
    .Y(_17185_));
 sky130_as_sc_hs__or2_2 _49205_ (.A(_17082_),
    .B(net1054),
    .Y(_17186_));
 sky130_as_sc_hs__or2_2 _49206_ (.A(\tholin_riscv.tmr0_pre[16] ),
    .B(_17186_),
    .Y(_17187_));
 sky130_as_sc_hs__nand3_2 _49207_ (.A(_17183_),
    .B(_17184_),
    .C(_17187_),
    .Y(_17188_));
 sky130_as_sc_hs__nor2_2 _49209_ (.A(net935),
    .B(_17082_),
    .Y(_17190_));
 sky130_as_sc_hs__or2_2 _49210_ (.A(_17083_),
    .B(net936),
    .Y(_17191_));
 sky130_as_sc_hs__nand3_2 _49212_ (.A(_17188_),
    .B(_17189_),
    .C(_17192_),
    .Y(_17193_));
 sky130_as_sc_hs__nor2_2 _49213_ (.A(net899),
    .B(_17083_),
    .Y(_17194_));
 sky130_as_sc_hs__or2_2 _49214_ (.A(_17084_),
    .B(net900),
    .Y(_17195_));
 sky130_as_sc_hs__or2_2 _49215_ (.A(\tholin_riscv.tmr0_pre[18] ),
    .B(_17195_),
    .Y(_17196_));
 sky130_as_sc_hs__or2_2 _49216_ (.A(\tholin_riscv.tmr0_pre[17] ),
    .B(_17191_),
    .Y(_17197_));
 sky130_as_sc_hs__nand3_2 _49217_ (.A(_17193_),
    .B(_17196_),
    .C(_17197_),
    .Y(_17198_));
 sky130_as_sc_hs__nand3_2 _49220_ (.A(_17198_),
    .B(_17199_),
    .C(_17200_),
    .Y(_17201_));
 sky130_as_sc_hs__nor2_2 _49223_ (.A(net891),
    .B(_17086_),
    .Y(_17204_));
 sky130_as_sc_hs__or2_2 _49224_ (.A(_17087_),
    .B(net892),
    .Y(_17205_));
 sky130_as_sc_hs__or2_2 _49225_ (.A(\tholin_riscv.tmr0_pre[21] ),
    .B(_17205_),
    .Y(_17206_));
 sky130_as_sc_hs__or2_2 _49226_ (.A(\tholin_riscv.tmr0_pre[20] ),
    .B(_17102_),
    .Y(_17207_));
 sky130_as_sc_hs__nand3_2 _49227_ (.A(_17203_),
    .B(_17206_),
    .C(_17207_),
    .Y(_17208_));
 sky130_as_sc_hs__nor2_2 _49228_ (.A(net931),
    .B(_17087_),
    .Y(_17209_));
 sky130_as_sc_hs__or2_2 _49229_ (.A(_17088_),
    .B(net932),
    .Y(_17210_));
 sky130_as_sc_hs__nand3_2 _49232_ (.A(_17208_),
    .B(_17211_),
    .C(_17212_),
    .Y(_17213_));
 sky130_as_sc_hs__nor2_2 _49233_ (.A(net1034),
    .B(_17088_),
    .Y(_17214_));
 sky130_as_sc_hs__or2_2 _49234_ (.A(_17089_),
    .B(net1035),
    .Y(_17215_));
 sky130_as_sc_hs__or2_2 _49235_ (.A(\tholin_riscv.tmr0_pre[23] ),
    .B(_17215_),
    .Y(_17216_));
 sky130_as_sc_hs__or2_2 _49236_ (.A(\tholin_riscv.tmr0_pre[22] ),
    .B(_17210_),
    .Y(_17217_));
 sky130_as_sc_hs__nand3_2 _49237_ (.A(_17213_),
    .B(_17216_),
    .C(_17217_),
    .Y(_17218_));
 sky130_as_sc_hs__nor2_2 _49238_ (.A(net992),
    .B(_17089_),
    .Y(_17219_));
 sky130_as_sc_hs__or2_2 _49239_ (.A(_17090_),
    .B(net993),
    .Y(_17220_));
 sky130_as_sc_hs__or2_2 _49242_ (.A(\tholin_riscv.tmr0_pre[24] ),
    .B(_17220_),
    .Y(_17223_));
 sky130_as_sc_hs__nor2_2 _49243_ (.A(net760),
    .B(_17090_),
    .Y(_17224_));
 sky130_as_sc_hs__nor2_2 _49244_ (.A(_17091_),
    .B(net761),
    .Y(_17225_));
 sky130_as_sc_hs__nor2_2 _49245_ (.A(net959),
    .B(_17091_),
    .Y(_17226_));
 sky130_as_sc_hs__or2_2 _49246_ (.A(_17092_),
    .B(net960),
    .Y(_17227_));
 sky130_as_sc_hs__nor2_2 _49248_ (.A(net1057),
    .B(_17092_),
    .Y(_17229_));
 sky130_as_sc_hs__or2_2 _49249_ (.A(_17093_),
    .B(net1058),
    .Y(_17230_));
 sky130_as_sc_hs__or2_2 _49250_ (.A(\tholin_riscv.tmr0_pre[27] ),
    .B(_17230_),
    .Y(_17231_));
 sky130_as_sc_hs__or2_2 _49251_ (.A(\tholin_riscv.tmr0_pre[26] ),
    .B(_17227_),
    .Y(_17232_));
 sky130_as_sc_hs__or2_2 _49257_ (.A(\tholin_riscv.tmr0_pre[25] ),
    .B(_17235_),
    .Y(_17238_));
 sky130_as_sc_hs__nand3_2 _49258_ (.A(_17232_),
    .B(_17237_),
    .C(_17238_),
    .Y(_17239_));
 sky130_as_sc_hs__nor2_2 _49261_ (.A(net1096),
    .B(_17093_),
    .Y(_17242_));
 sky130_as_sc_hs__or2_2 _49262_ (.A(_17094_),
    .B(net1097),
    .Y(_17243_));
 sky130_as_sc_hs__nand3_2 _49265_ (.A(_17241_),
    .B(_17244_),
    .C(_17245_),
    .Y(_17246_));
 sky130_as_sc_hs__nor2_2 _49266_ (.A(net955),
    .B(_17094_),
    .Y(_17247_));
 sky130_as_sc_hs__or2_2 _49267_ (.A(_17095_),
    .B(net956),
    .Y(_17248_));
 sky130_as_sc_hs__or2_2 _49268_ (.A(\tholin_riscv.tmr0_pre[29] ),
    .B(_17248_),
    .Y(_17249_));
 sky130_as_sc_hs__or2_2 _49269_ (.A(\tholin_riscv.tmr0_pre[28] ),
    .B(_17243_),
    .Y(_17250_));
 sky130_as_sc_hs__nand3_2 _49270_ (.A(_17246_),
    .B(_17249_),
    .C(_17250_),
    .Y(_17251_));
 sky130_as_sc_hs__nor2_2 _49271_ (.A(net775),
    .B(_17095_),
    .Y(_17252_));
 sky130_as_sc_hs__or2_2 _49272_ (.A(net776),
    .B(_17252_),
    .Y(_17253_));
 sky130_as_sc_hs__nand3_2 _49275_ (.A(_17251_),
    .B(_17254_),
    .C(_17255_),
    .Y(_17256_));
 sky130_as_sc_hs__or2_2 _49276_ (.A(\tholin_riscv.tmr0_pre[31] ),
    .B(_17099_),
    .Y(_17257_));
 sky130_as_sc_hs__or2_2 _49277_ (.A(\tholin_riscv.tmr0_pre[30] ),
    .B(_17253_),
    .Y(_17258_));
 sky130_as_sc_hs__nand3_2 _49278_ (.A(_17256_),
    .B(_17257_),
    .C(_17258_),
    .Y(_17259_));
 sky130_as_sc_hs__inv_2 _49281_ (.Y(_17262_),
    .A(_17261_));
 sky130_as_sc_hs__nor2_2 _49282_ (.A(net1714),
    .B(_17261_),
    .Y(_01312_));
 sky130_as_sc_hs__nor2_2 _49283_ (.A(net749),
    .B(_17261_),
    .Y(_01313_));
 sky130_as_sc_hs__nor2_2 _49284_ (.A(net886),
    .B(_17261_),
    .Y(_01314_));
 sky130_as_sc_hs__nor2_2 _49285_ (.A(net965),
    .B(_17261_),
    .Y(_01315_));
 sky130_as_sc_hs__nor2_2 _49286_ (.A(net986),
    .B(_17261_),
    .Y(_01316_));
 sky130_as_sc_hs__nor2_2 _49287_ (.A(net882),
    .B(_17261_),
    .Y(_01317_));
 sky130_as_sc_hs__nor2_2 _49288_ (.A(net1111),
    .B(_17261_),
    .Y(_01318_));
 sky130_as_sc_hs__nor2_2 _49289_ (.A(net929),
    .B(_17261_),
    .Y(_01319_));
 sky130_as_sc_hs__nor2_2 _49290_ (.A(net1006),
    .B(_17261_),
    .Y(_01320_));
 sky130_as_sc_hs__nor2_2 _49291_ (.A(net1010),
    .B(_17261_),
    .Y(_01321_));
 sky130_as_sc_hs__nor2_2 _49292_ (.A(net982),
    .B(_17261_),
    .Y(_01322_));
 sky130_as_sc_hs__nor2_2 _49293_ (.A(net978),
    .B(_17261_),
    .Y(_01323_));
 sky130_as_sc_hs__nor2_2 _49294_ (.A(net1030),
    .B(_17261_),
    .Y(_01324_));
 sky130_as_sc_hs__nor2_2 _49295_ (.A(net921),
    .B(_17261_),
    .Y(_01325_));
 sky130_as_sc_hs__nor2_2 _49296_ (.A(net998),
    .B(_17261_),
    .Y(_01326_));
 sky130_as_sc_hs__nor2_2 _49297_ (.A(net1067),
    .B(_17261_),
    .Y(_01327_));
 sky130_as_sc_hs__nor2_2 _49298_ (.A(net1055),
    .B(_17261_),
    .Y(_01328_));
 sky130_as_sc_hs__nor2_2 _49299_ (.A(net937),
    .B(_17261_),
    .Y(_01329_));
 sky130_as_sc_hs__nor2_2 _49300_ (.A(net901),
    .B(_17261_),
    .Y(_01330_));
 sky130_as_sc_hs__nor2_2 _49301_ (.A(net1040),
    .B(_17261_),
    .Y(_01331_));
 sky130_as_sc_hs__nor2_2 _49302_ (.A(net913),
    .B(_17261_),
    .Y(_01332_));
 sky130_as_sc_hs__nor2_2 _49303_ (.A(net893),
    .B(_17261_),
    .Y(_01333_));
 sky130_as_sc_hs__nor2_2 _49304_ (.A(net933),
    .B(_17261_),
    .Y(_01334_));
 sky130_as_sc_hs__nor2_2 _49305_ (.A(net1036),
    .B(_17261_),
    .Y(_01335_));
 sky130_as_sc_hs__nor2_2 _49306_ (.A(net994),
    .B(_17261_),
    .Y(_01336_));
 sky130_as_sc_hs__and2_2 _49307_ (.A(net762),
    .B(_17262_),
    .Y(_01337_));
 sky130_as_sc_hs__nor2_2 _49308_ (.A(net961),
    .B(_17261_),
    .Y(_01338_));
 sky130_as_sc_hs__nor2_2 _49309_ (.A(net1059),
    .B(_17261_),
    .Y(_01339_));
 sky130_as_sc_hs__nor2_2 _49310_ (.A(net1098),
    .B(_17261_),
    .Y(_01340_));
 sky130_as_sc_hs__nor2_2 _49311_ (.A(net957),
    .B(_17261_),
    .Y(_01341_));
 sky130_as_sc_hs__nor2_2 _49312_ (.A(net777),
    .B(_17261_),
    .Y(_01342_));
 sky130_as_sc_hs__nor2_2 _49313_ (.A(_17099_),
    .B(_17261_),
    .Y(_01343_));
 sky130_as_sc_hs__and2_2 _49314_ (.A(_19901_),
    .B(_20032_),
    .Y(_17263_));
 sky130_as_sc_hs__nor2_2 _49319_ (.A(\tholin_riscv.tmr1_top[30] ),
    .B(_19722_),
    .Y(_17268_));
 sky130_as_sc_hs__nor2_2 _49320_ (.A(\tholin_riscv.tmr1_top[31] ),
    .B(_19721_),
    .Y(_17269_));
 sky130_as_sc_hs__nor2_2 _49321_ (.A(_17268_),
    .B(_17269_),
    .Y(_17270_));
 sky130_as_sc_hs__nor2_2 _49322_ (.A(\tholin_riscv.tmr1_top[29] ),
    .B(_19723_),
    .Y(_17271_));
 sky130_as_sc_hs__nor2_2 _49323_ (.A(\tholin_riscv.tmr1_top[28] ),
    .B(_19724_),
    .Y(_17272_));
 sky130_as_sc_hs__nor2_2 _49324_ (.A(_17271_),
    .B(_17272_),
    .Y(_17273_));
 sky130_as_sc_hs__nor2_2 _49325_ (.A(\tholin_riscv.tmr1_top[27] ),
    .B(_19725_),
    .Y(_17274_));
 sky130_as_sc_hs__nor2_2 _49326_ (.A(\tholin_riscv.tmr1_top[26] ),
    .B(_19726_),
    .Y(_17275_));
 sky130_as_sc_hs__nor2_2 _49327_ (.A(_17274_),
    .B(_17275_),
    .Y(_17276_));
 sky130_as_sc_hs__nor2_2 _49328_ (.A(\tholin_riscv.tmr1_top[24] ),
    .B(_19691_),
    .Y(_17277_));
 sky130_as_sc_hs__nor2_2 _49329_ (.A(\tholin_riscv.tmr1_top[25] ),
    .B(_19727_),
    .Y(_17278_));
 sky130_as_sc_hs__or2_2 _49330_ (.A(_17277_),
    .B(_17278_),
    .Y(_17279_));
 sky130_as_sc_hs__and2_2 _49333_ (.A(_17280_),
    .B(_17281_),
    .Y(_17282_));
 sky130_as_sc_hs__and2_2 _49338_ (.A(_17285_),
    .B(_17286_),
    .Y(_17287_));
 sky130_as_sc_hs__and2_2 _49343_ (.A(_17290_),
    .B(_17291_),
    .Y(_17292_));
 sky130_as_sc_hs__nor2_2 _49348_ (.A(\tholin_riscv.tmr1_top[22] ),
    .B(_19687_),
    .Y(_17297_));
 sky130_as_sc_hs__nor2_2 _49349_ (.A(\tholin_riscv.tmr1_top[23] ),
    .B(_19689_),
    .Y(_17298_));
 sky130_as_sc_hs__nor2_2 _49350_ (.A(_17297_),
    .B(_17298_),
    .Y(_17299_));
 sky130_as_sc_hs__nor2_2 _49351_ (.A(\tholin_riscv.tmr1_top[21] ),
    .B(_19685_),
    .Y(_17300_));
 sky130_as_sc_hs__nor2_2 _49352_ (.A(\tholin_riscv.tmr1_top[20] ),
    .B(_19683_),
    .Y(_17301_));
 sky130_as_sc_hs__nor2_2 _49353_ (.A(_17300_),
    .B(_17301_),
    .Y(_17302_));
 sky130_as_sc_hs__nor2_2 _49354_ (.A(\tholin_riscv.tmr1_top[19] ),
    .B(_19728_),
    .Y(_17303_));
 sky130_as_sc_hs__nor2_2 _49355_ (.A(\tholin_riscv.tmr1_top[18] ),
    .B(_19729_),
    .Y(_17304_));
 sky130_as_sc_hs__nor2_2 _49356_ (.A(_17303_),
    .B(_17304_),
    .Y(_17305_));
 sky130_as_sc_hs__nor2_2 _49357_ (.A(\tholin_riscv.tmr1_top[16] ),
    .B(_19731_),
    .Y(_17306_));
 sky130_as_sc_hs__nor2_2 _49358_ (.A(\tholin_riscv.tmr1_top[17] ),
    .B(_19730_),
    .Y(_17307_));
 sky130_as_sc_hs__or2_2 _49359_ (.A(_17306_),
    .B(_17307_),
    .Y(_17308_));
 sky130_as_sc_hs__and2_2 _49362_ (.A(_17309_),
    .B(_17310_),
    .Y(_17311_));
 sky130_as_sc_hs__and2_2 _49367_ (.A(_17314_),
    .B(_17315_),
    .Y(_17316_));
 sky130_as_sc_hs__and2_2 _49372_ (.A(_17319_),
    .B(_17320_),
    .Y(_17321_));
 sky130_as_sc_hs__nor2_2 _49376_ (.A(\tholin_riscv.tmr1_top[14] ),
    .B(_19733_),
    .Y(_17325_));
 sky130_as_sc_hs__nor2_2 _49377_ (.A(\tholin_riscv.tmr1_top[15] ),
    .B(_19732_),
    .Y(_17326_));
 sky130_as_sc_hs__or2_2 _49378_ (.A(_17325_),
    .B(_17326_),
    .Y(_17327_));
 sky130_as_sc_hs__or2_2 _49381_ (.A(\tholin_riscv.tmr1_top[13] ),
    .B(_19734_),
    .Y(_17330_));
 sky130_as_sc_hs__or2_2 _49382_ (.A(\tholin_riscv.tmr1_top[12] ),
    .B(_19735_),
    .Y(_17331_));
 sky130_as_sc_hs__nor2_2 _49384_ (.A(\tholin_riscv.tmr1_top[11] ),
    .B(_19736_),
    .Y(_17333_));
 sky130_as_sc_hs__nor2_2 _49385_ (.A(\tholin_riscv.tmr1_top[10] ),
    .B(_19737_),
    .Y(_17334_));
 sky130_as_sc_hs__or2_2 _49386_ (.A(_17333_),
    .B(_17334_),
    .Y(_17335_));
 sky130_as_sc_hs__or2_2 _49389_ (.A(\tholin_riscv.tmr1_top[8] ),
    .B(_19739_),
    .Y(_17338_));
 sky130_as_sc_hs__or2_2 _49390_ (.A(\tholin_riscv.tmr1_top[9] ),
    .B(_19738_),
    .Y(_17339_));
 sky130_as_sc_hs__or2_2 _49392_ (.A(\tholin_riscv.tmr1_top[1] ),
    .B(_19746_),
    .Y(_17341_));
 sky130_as_sc_hs__nand3_2 _49394_ (.A(\tholin_riscv.tmr1_top[0] ),
    .B(_19747_),
    .C(_17341_),
    .Y(_17343_));
 sky130_as_sc_hs__nand3_2 _49395_ (.A(_17340_),
    .B(_17342_),
    .C(_17343_),
    .Y(_17344_));
 sky130_as_sc_hs__or2_2 _49396_ (.A(\tholin_riscv.tmr1_top[3] ),
    .B(_19744_),
    .Y(_17345_));
 sky130_as_sc_hs__or2_2 _49397_ (.A(\tholin_riscv.tmr1_top[2] ),
    .B(_19745_),
    .Y(_17346_));
 sky130_as_sc_hs__nand3_2 _49398_ (.A(_17344_),
    .B(_17345_),
    .C(_17346_),
    .Y(_17347_));
 sky130_as_sc_hs__nand3_2 _49401_ (.A(_17347_),
    .B(_17348_),
    .C(_17349_),
    .Y(_17350_));
 sky130_as_sc_hs__or2_2 _49402_ (.A(\tholin_riscv.tmr1_top[5] ),
    .B(_19742_),
    .Y(_17351_));
 sky130_as_sc_hs__or2_2 _49403_ (.A(\tholin_riscv.tmr1_top[4] ),
    .B(_19743_),
    .Y(_17352_));
 sky130_as_sc_hs__nand3_2 _49404_ (.A(_17350_),
    .B(_17351_),
    .C(_17352_),
    .Y(_17353_));
 sky130_as_sc_hs__or2_2 _49405_ (.A(\tholin_riscv.tmr1_top[6] ),
    .B(_19741_),
    .Y(_17354_));
 sky130_as_sc_hs__and2_2 _49407_ (.A(_17354_),
    .B(_17355_),
    .Y(_17356_));
 sky130_as_sc_hs__and2_2 _49410_ (.A(_17357_),
    .B(_17358_),
    .Y(_17359_));
 sky130_as_sc_hs__nand3_2 _49411_ (.A(_17353_),
    .B(_17356_),
    .C(_17359_),
    .Y(_17360_));
 sky130_as_sc_hs__nand2b_2 _49412_ (.B(_17355_),
    .Y(_17361_),
    .A(_17354_));
 sky130_as_sc_hs__or2_2 _49413_ (.A(\tholin_riscv.tmr1_top[7] ),
    .B(_19740_),
    .Y(_17362_));
 sky130_as_sc_hs__nand3_2 _49414_ (.A(_17360_),
    .B(_17361_),
    .C(_17362_),
    .Y(_17363_));
 sky130_as_sc_hs__nand3_2 _49417_ (.A(_17338_),
    .B(_17339_),
    .C(_17365_),
    .Y(_17366_));
 sky130_as_sc_hs__nand3_2 _49420_ (.A(_17336_),
    .B(_17367_),
    .C(_17368_),
    .Y(_17369_));
 sky130_as_sc_hs__nor2_2 _49421_ (.A(_17335_),
    .B(_17369_),
    .Y(_17370_));
 sky130_as_sc_hs__nand3_2 _49425_ (.A(_17330_),
    .B(_17331_),
    .C(_17373_),
    .Y(_17374_));
 sky130_as_sc_hs__nand3_2 _49428_ (.A(_17328_),
    .B(_17375_),
    .C(_17376_),
    .Y(_17377_));
 sky130_as_sc_hs__nor2_2 _49429_ (.A(_17327_),
    .B(_17377_),
    .Y(_17378_));
 sky130_as_sc_hs__nand2b_2 _49432_ (.B(_17311_),
    .Y(_17381_),
    .A(_17308_));
 sky130_as_sc_hs__nor2_2 _49434_ (.A(_17381_),
    .B(_17382_),
    .Y(_17383_));
 sky130_as_sc_hs__nand3_2 _49436_ (.A(_17296_),
    .B(_17299_),
    .C(_17384_),
    .Y(_17385_));
 sky130_as_sc_hs__nor2_2 _49438_ (.A(_17385_),
    .B(_17386_),
    .Y(_17387_));
 sky130_as_sc_hs__nand3_2 _49439_ (.A(_17380_),
    .B(_17383_),
    .C(_17387_),
    .Y(_17388_));
 sky130_as_sc_hs__nand2b_2 _49441_ (.B(_17282_),
    .Y(_17390_),
    .A(_17279_));
 sky130_as_sc_hs__nor2_2 _49443_ (.A(_17390_),
    .B(_17391_),
    .Y(_17392_));
 sky130_as_sc_hs__nand3_2 _49445_ (.A(_17267_),
    .B(_17270_),
    .C(_17393_),
    .Y(_17394_));
 sky130_as_sc_hs__nor2_2 _49447_ (.A(_17394_),
    .B(_17395_),
    .Y(_17396_));
 sky130_as_sc_hs__nand3_2 _49448_ (.A(_17389_),
    .B(_17392_),
    .C(_17396_),
    .Y(_17397_));
 sky130_as_sc_hs__and2_2 _49449_ (.A(_17295_),
    .B(_17397_),
    .Y(_17398_));
 sky130_as_sc_hs__and2_2 _49450_ (.A(_19747_),
    .B(net97),
    .Y(_17399_));
 sky130_as_sc_hs__nor2_2 _49451_ (.A(_16370_),
    .B(_17399_),
    .Y(_17400_));
 sky130_as_sc_hs__nor2_2 _49452_ (.A(_17263_),
    .B(_17400_),
    .Y(_17401_));
 sky130_as_sc_hs__and2_2 _49455_ (.A(net506),
    .B(_17403_),
    .Y(_01344_));
 sky130_as_sc_hs__nor2b_2 _49456_ (.A(_16370_),
    .Y(_17404_),
    .B(net96));
 sky130_as_sc_hs__nand3_2 _49457_ (.A(_19746_),
    .B(net783),
    .C(net81),
    .Y(_17405_));
 sky130_as_sc_hs__or2_2 _49458_ (.A(_19746_),
    .B(_17400_),
    .Y(_17406_));
 sky130_as_sc_hs__nand3_2 _49459_ (.A(_17264_),
    .B(net784),
    .C(_17406_),
    .Y(_17407_));
 sky130_as_sc_hs__or2_2 _49460_ (.A(\tholin_riscv.instr[1] ),
    .B(_17264_),
    .Y(_17408_));
 sky130_as_sc_hs__and2_2 _49461_ (.A(net506),
    .B(_17408_),
    .Y(_17409_));
 sky130_as_sc_hs__and2_2 _49462_ (.A(net785),
    .B(_17409_),
    .Y(_01345_));
 sky130_as_sc_hs__nor2_2 _49464_ (.A(\tholin_riscv.tmr1[2] ),
    .B(_17410_),
    .Y(_17411_));
 sky130_as_sc_hs__and2_2 _49466_ (.A(net97),
    .B(_17410_),
    .Y(_17413_));
 sky130_as_sc_hs__or2_2 _49467_ (.A(_16370_),
    .B(_17413_),
    .Y(_17414_));
 sky130_as_sc_hs__nand3_2 _49469_ (.A(_17264_),
    .B(_17412_),
    .C(_17415_),
    .Y(_17416_));
 sky130_as_sc_hs__and2_2 _49471_ (.A(net506),
    .B(_17417_),
    .Y(_17418_));
 sky130_as_sc_hs__and2_2 _49472_ (.A(_17416_),
    .B(_17418_),
    .Y(_01346_));
 sky130_as_sc_hs__nor2_2 _49473_ (.A(_19745_),
    .B(_17410_),
    .Y(_17419_));
 sky130_as_sc_hs__inv_2 _49474_ (.Y(_17420_),
    .A(_17419_));
 sky130_as_sc_hs__nand3_2 _49475_ (.A(net1128),
    .B(net81),
    .C(_17419_),
    .Y(_17421_));
 sky130_as_sc_hs__and2_2 _49476_ (.A(net97),
    .B(_17420_),
    .Y(_17422_));
 sky130_as_sc_hs__or2_2 _49477_ (.A(_16370_),
    .B(_17422_),
    .Y(_17423_));
 sky130_as_sc_hs__nand3_2 _49479_ (.A(_17264_),
    .B(net1129),
    .C(_17424_),
    .Y(_17425_));
 sky130_as_sc_hs__and2_2 _49481_ (.A(net505),
    .B(_17426_),
    .Y(_17427_));
 sky130_as_sc_hs__and2_2 _49482_ (.A(net1130),
    .B(_17427_),
    .Y(_01347_));
 sky130_as_sc_hs__and2_2 _49483_ (.A(\tholin_riscv.tmr1[3] ),
    .B(_17419_),
    .Y(_17428_));
 sky130_as_sc_hs__inv_2 _49484_ (.Y(_17429_),
    .A(_17428_));
 sky130_as_sc_hs__nand3_2 _49485_ (.A(net803),
    .B(net81),
    .C(_17428_),
    .Y(_17430_));
 sky130_as_sc_hs__and2_2 _49486_ (.A(net97),
    .B(_17429_),
    .Y(_17431_));
 sky130_as_sc_hs__or2_2 _49487_ (.A(_16370_),
    .B(_17431_),
    .Y(_17432_));
 sky130_as_sc_hs__nand3_2 _49489_ (.A(_17264_),
    .B(net804),
    .C(_17433_),
    .Y(_17434_));
 sky130_as_sc_hs__and2_2 _49491_ (.A(net505),
    .B(_17435_),
    .Y(_17436_));
 sky130_as_sc_hs__and2_2 _49492_ (.A(net805),
    .B(_17436_),
    .Y(_01348_));
 sky130_as_sc_hs__nor2_2 _49494_ (.A(\tholin_riscv.tmr1[5] ),
    .B(_17437_),
    .Y(_17438_));
 sky130_as_sc_hs__and2_2 _49496_ (.A(net96),
    .B(_17437_),
    .Y(_17440_));
 sky130_as_sc_hs__or2_2 _49497_ (.A(_16370_),
    .B(_17440_),
    .Y(_17441_));
 sky130_as_sc_hs__nand3_2 _49499_ (.A(_17264_),
    .B(_17439_),
    .C(_17442_),
    .Y(_17443_));
 sky130_as_sc_hs__and2_2 _49501_ (.A(net505),
    .B(_17444_),
    .Y(_17445_));
 sky130_as_sc_hs__and2_2 _49502_ (.A(_17443_),
    .B(_17445_),
    .Y(_01349_));
 sky130_as_sc_hs__nor2_2 _49503_ (.A(_19742_),
    .B(_17437_),
    .Y(_17446_));
 sky130_as_sc_hs__inv_2 _49504_ (.Y(_17447_),
    .A(_17446_));
 sky130_as_sc_hs__nand3_2 _49505_ (.A(net1159),
    .B(net81),
    .C(_17446_),
    .Y(_17448_));
 sky130_as_sc_hs__and2_2 _49506_ (.A(net96),
    .B(_17447_),
    .Y(_17449_));
 sky130_as_sc_hs__or2_2 _49507_ (.A(_16370_),
    .B(_17449_),
    .Y(_17450_));
 sky130_as_sc_hs__nand3_2 _49509_ (.A(_17264_),
    .B(net1160),
    .C(_17451_),
    .Y(_17452_));
 sky130_as_sc_hs__and2_2 _49511_ (.A(net507),
    .B(_17453_),
    .Y(_17454_));
 sky130_as_sc_hs__and2_2 _49512_ (.A(net1161),
    .B(_17454_),
    .Y(_01350_));
 sky130_as_sc_hs__and2_2 _49513_ (.A(\tholin_riscv.tmr1[6] ),
    .B(_17446_),
    .Y(_17455_));
 sky130_as_sc_hs__inv_2 _49514_ (.Y(_17456_),
    .A(_17455_));
 sky130_as_sc_hs__nand3_2 _49515_ (.A(net856),
    .B(net81),
    .C(_17455_),
    .Y(_17457_));
 sky130_as_sc_hs__and2_2 _49516_ (.A(net96),
    .B(_17456_),
    .Y(_17458_));
 sky130_as_sc_hs__or2_2 _49517_ (.A(_16370_),
    .B(_17458_),
    .Y(_17459_));
 sky130_as_sc_hs__nand3_2 _49519_ (.A(_17264_),
    .B(net857),
    .C(_17460_),
    .Y(_17461_));
 sky130_as_sc_hs__or2_2 _49520_ (.A(\tholin_riscv.Bimm[11] ),
    .B(_17264_),
    .Y(_17462_));
 sky130_as_sc_hs__and2_2 _49521_ (.A(net507),
    .B(_17462_),
    .Y(_17463_));
 sky130_as_sc_hs__and2_2 _49522_ (.A(net858),
    .B(_17463_),
    .Y(_01351_));
 sky130_as_sc_hs__nor2_2 _49524_ (.A(\tholin_riscv.tmr1[8] ),
    .B(_17464_),
    .Y(_17465_));
 sky130_as_sc_hs__and2_2 _49526_ (.A(net98),
    .B(_17464_),
    .Y(_17467_));
 sky130_as_sc_hs__or2_2 _49527_ (.A(_16370_),
    .B(_17467_),
    .Y(_17468_));
 sky130_as_sc_hs__nand3_2 _49529_ (.A(_17264_),
    .B(_17466_),
    .C(_17469_),
    .Y(_17470_));
 sky130_as_sc_hs__or2_2 _49530_ (.A(net1260),
    .B(_17264_),
    .Y(_17471_));
 sky130_as_sc_hs__and2_2 _49531_ (.A(net512),
    .B(_17471_),
    .Y(_17472_));
 sky130_as_sc_hs__and2_2 _49532_ (.A(_17470_),
    .B(_17472_),
    .Y(_01352_));
 sky130_as_sc_hs__nor2_2 _49533_ (.A(_19739_),
    .B(_17464_),
    .Y(_17473_));
 sky130_as_sc_hs__inv_2 _49534_ (.Y(_17474_),
    .A(_17473_));
 sky130_as_sc_hs__nand3_2 _49535_ (.A(net1070),
    .B(net81),
    .C(_17473_),
    .Y(_17475_));
 sky130_as_sc_hs__and2_2 _49536_ (.A(net98),
    .B(_17474_),
    .Y(_17476_));
 sky130_as_sc_hs__or2_2 _49537_ (.A(_16370_),
    .B(_17476_),
    .Y(_17477_));
 sky130_as_sc_hs__nand3_2 _49539_ (.A(_17264_),
    .B(net1071),
    .C(_17478_),
    .Y(_17479_));
 sky130_as_sc_hs__or2_2 _49540_ (.A(\tholin_riscv.Bimm[2] ),
    .B(_17264_),
    .Y(_17480_));
 sky130_as_sc_hs__and2_2 _49541_ (.A(net512),
    .B(_17480_),
    .Y(_17481_));
 sky130_as_sc_hs__and2_2 _49542_ (.A(_17479_),
    .B(_17481_),
    .Y(_01353_));
 sky130_as_sc_hs__and2_2 _49543_ (.A(\tholin_riscv.tmr1[9] ),
    .B(_17473_),
    .Y(_17482_));
 sky130_as_sc_hs__inv_2 _49544_ (.Y(_17483_),
    .A(_17482_));
 sky130_as_sc_hs__nand3_2 _49545_ (.A(net815),
    .B(net81),
    .C(_17482_),
    .Y(_17484_));
 sky130_as_sc_hs__and2_2 _49546_ (.A(net98),
    .B(_17483_),
    .Y(_17485_));
 sky130_as_sc_hs__or2_2 _49547_ (.A(_16370_),
    .B(_17485_),
    .Y(_17486_));
 sky130_as_sc_hs__nand3_2 _49549_ (.A(_17264_),
    .B(net816),
    .C(_17487_),
    .Y(_17488_));
 sky130_as_sc_hs__or2_2 _49550_ (.A(net1791),
    .B(_17264_),
    .Y(_17489_));
 sky130_as_sc_hs__and2_2 _49551_ (.A(net512),
    .B(_17489_),
    .Y(_17490_));
 sky130_as_sc_hs__and2_2 _49552_ (.A(net817),
    .B(_17490_),
    .Y(_01354_));
 sky130_as_sc_hs__nor2_2 _49554_ (.A(\tholin_riscv.tmr1[11] ),
    .B(_17491_),
    .Y(_17492_));
 sky130_as_sc_hs__and2_2 _49556_ (.A(net97),
    .B(_17491_),
    .Y(_17494_));
 sky130_as_sc_hs__or2_2 _49557_ (.A(_16370_),
    .B(_17494_),
    .Y(_17495_));
 sky130_as_sc_hs__nand3_2 _49559_ (.A(_17264_),
    .B(_17493_),
    .C(_17496_),
    .Y(_17497_));
 sky130_as_sc_hs__or2_2 _49560_ (.A(net1792),
    .B(_17264_),
    .Y(_17498_));
 sky130_as_sc_hs__and2_2 _49561_ (.A(net507),
    .B(_17498_),
    .Y(_17499_));
 sky130_as_sc_hs__and2_2 _49562_ (.A(_17497_),
    .B(_17499_),
    .Y(_01355_));
 sky130_as_sc_hs__nor2_2 _49563_ (.A(_19736_),
    .B(_17491_),
    .Y(_17500_));
 sky130_as_sc_hs__inv_2 _49564_ (.Y(_17501_),
    .A(_17500_));
 sky130_as_sc_hs__nand3_2 _49565_ (.A(net1311),
    .B(_17404_),
    .C(_17500_),
    .Y(_17502_));
 sky130_as_sc_hs__and2_2 _49566_ (.A(net97),
    .B(_17501_),
    .Y(_17503_));
 sky130_as_sc_hs__or2_2 _49567_ (.A(_16370_),
    .B(_17503_),
    .Y(_17504_));
 sky130_as_sc_hs__nand3_2 _49569_ (.A(_17264_),
    .B(net1312),
    .C(_17505_),
    .Y(_17506_));
 sky130_as_sc_hs__and2_2 _49571_ (.A(net507),
    .B(_17507_),
    .Y(_17508_));
 sky130_as_sc_hs__and2_2 _49572_ (.A(_17506_),
    .B(_17508_),
    .Y(_01356_));
 sky130_as_sc_hs__and2_2 _49573_ (.A(\tholin_riscv.tmr1[12] ),
    .B(_17500_),
    .Y(_17509_));
 sky130_as_sc_hs__inv_2 _49574_ (.Y(_17510_),
    .A(_17509_));
 sky130_as_sc_hs__nand3_2 _49575_ (.A(net799),
    .B(_17404_),
    .C(_17509_),
    .Y(_17511_));
 sky130_as_sc_hs__and2_2 _49576_ (.A(net97),
    .B(_17510_),
    .Y(_17512_));
 sky130_as_sc_hs__or2_2 _49577_ (.A(_16370_),
    .B(_17512_),
    .Y(_17513_));
 sky130_as_sc_hs__nand3_2 _49579_ (.A(_17264_),
    .B(net800),
    .C(_17514_),
    .Y(_17515_));
 sky130_as_sc_hs__and2_2 _49581_ (.A(net507),
    .B(_17516_),
    .Y(_17517_));
 sky130_as_sc_hs__and2_2 _49582_ (.A(net801),
    .B(_17517_),
    .Y(_01357_));
 sky130_as_sc_hs__nor2_2 _49584_ (.A(\tholin_riscv.tmr1[14] ),
    .B(_17518_),
    .Y(_17519_));
 sky130_as_sc_hs__and2_2 _49586_ (.A(net96),
    .B(_17518_),
    .Y(_17521_));
 sky130_as_sc_hs__or2_2 _49587_ (.A(_16370_),
    .B(_17521_),
    .Y(_17522_));
 sky130_as_sc_hs__nand3_2 _49589_ (.A(_17264_),
    .B(_17520_),
    .C(_17523_),
    .Y(_17524_));
 sky130_as_sc_hs__or2_2 _49590_ (.A(net1796),
    .B(_17264_),
    .Y(_17525_));
 sky130_as_sc_hs__and2_2 _49591_ (.A(net508),
    .B(_17525_),
    .Y(_17526_));
 sky130_as_sc_hs__and2_2 _49592_ (.A(_17524_),
    .B(_17526_),
    .Y(_01358_));
 sky130_as_sc_hs__nor2_2 _49593_ (.A(_19733_),
    .B(_17518_),
    .Y(_17527_));
 sky130_as_sc_hs__inv_2 _49594_ (.Y(_17528_),
    .A(_17527_));
 sky130_as_sc_hs__nand3_2 _49595_ (.A(net1252),
    .B(net81),
    .C(_17527_),
    .Y(_17529_));
 sky130_as_sc_hs__and2_2 _49596_ (.A(net96),
    .B(_17528_),
    .Y(_17530_));
 sky130_as_sc_hs__or2_2 _49597_ (.A(_16370_),
    .B(_17530_),
    .Y(_17531_));
 sky130_as_sc_hs__nand3_2 _49599_ (.A(_17264_),
    .B(net1253),
    .C(_17532_),
    .Y(_17533_));
 sky130_as_sc_hs__and2_2 _49601_ (.A(net507),
    .B(_17534_),
    .Y(_17535_));
 sky130_as_sc_hs__and2_2 _49602_ (.A(_17533_),
    .B(_17535_),
    .Y(_01359_));
 sky130_as_sc_hs__and2_2 _49603_ (.A(\tholin_riscv.tmr1[15] ),
    .B(_17527_),
    .Y(_17536_));
 sky130_as_sc_hs__inv_2 _49604_ (.Y(_17537_),
    .A(_17536_));
 sky130_as_sc_hs__nand3_2 _49605_ (.A(net831),
    .B(net81),
    .C(_17536_),
    .Y(_17538_));
 sky130_as_sc_hs__and2_2 _49606_ (.A(net96),
    .B(_17537_),
    .Y(_17539_));
 sky130_as_sc_hs__or2_2 _49607_ (.A(_16370_),
    .B(_17539_),
    .Y(_17540_));
 sky130_as_sc_hs__nand3_2 _49609_ (.A(_17264_),
    .B(net832),
    .C(_17541_),
    .Y(_17542_));
 sky130_as_sc_hs__and2_2 _49611_ (.A(net507),
    .B(_17543_),
    .Y(_17544_));
 sky130_as_sc_hs__and2_2 _49612_ (.A(net833),
    .B(_17544_),
    .Y(_01360_));
 sky130_as_sc_hs__nor2_2 _49614_ (.A(\tholin_riscv.tmr1[17] ),
    .B(_17545_),
    .Y(_17546_));
 sky130_as_sc_hs__and2_2 _49616_ (.A(net96),
    .B(_17545_),
    .Y(_17548_));
 sky130_as_sc_hs__or2_2 _49617_ (.A(_16370_),
    .B(_17548_),
    .Y(_17549_));
 sky130_as_sc_hs__nand3_2 _49619_ (.A(_17264_),
    .B(_17547_),
    .C(_17550_),
    .Y(_17551_));
 sky130_as_sc_hs__and2_2 _49621_ (.A(net507),
    .B(_17552_),
    .Y(_17553_));
 sky130_as_sc_hs__and2_2 _49622_ (.A(_17551_),
    .B(_17553_),
    .Y(_01361_));
 sky130_as_sc_hs__nor2_2 _49623_ (.A(_19730_),
    .B(_17545_),
    .Y(_17554_));
 sky130_as_sc_hs__inv_2 _49624_ (.Y(_17555_),
    .A(_17554_));
 sky130_as_sc_hs__nand3_2 _49625_ (.A(net1335),
    .B(net81),
    .C(_17554_),
    .Y(_17556_));
 sky130_as_sc_hs__and2_2 _49626_ (.A(net96),
    .B(_17555_),
    .Y(_17557_));
 sky130_as_sc_hs__or2_2 _49627_ (.A(_16370_),
    .B(_17557_),
    .Y(_17558_));
 sky130_as_sc_hs__nand3_2 _49629_ (.A(_17264_),
    .B(net1336),
    .C(_17559_),
    .Y(_17560_));
 sky130_as_sc_hs__and2_2 _49631_ (.A(net507),
    .B(_17561_),
    .Y(_17562_));
 sky130_as_sc_hs__and2_2 _49632_ (.A(_17560_),
    .B(_17562_),
    .Y(_01362_));
 sky130_as_sc_hs__and2_2 _49633_ (.A(\tholin_riscv.tmr1[18] ),
    .B(_17554_),
    .Y(_17563_));
 sky130_as_sc_hs__inv_2 _49634_ (.Y(_17564_),
    .A(_17563_));
 sky130_as_sc_hs__nand3_2 _49635_ (.A(net840),
    .B(net81),
    .C(_17563_),
    .Y(_17565_));
 sky130_as_sc_hs__and2_2 _49636_ (.A(net96),
    .B(_17564_),
    .Y(_17566_));
 sky130_as_sc_hs__or2_2 _49637_ (.A(_16370_),
    .B(_17566_),
    .Y(_17567_));
 sky130_as_sc_hs__nand3_2 _49639_ (.A(_17264_),
    .B(net841),
    .C(_17568_),
    .Y(_17569_));
 sky130_as_sc_hs__and2_2 _49641_ (.A(net507),
    .B(_17570_),
    .Y(_17571_));
 sky130_as_sc_hs__and2_2 _49642_ (.A(net842),
    .B(_17571_),
    .Y(_01363_));
 sky130_as_sc_hs__nor2_2 _49644_ (.A(\tholin_riscv.tmr1[20] ),
    .B(_17572_),
    .Y(_17573_));
 sky130_as_sc_hs__and2_2 _49646_ (.A(net96),
    .B(_17572_),
    .Y(_17575_));
 sky130_as_sc_hs__or2_2 _49647_ (.A(_16370_),
    .B(_17575_),
    .Y(_17576_));
 sky130_as_sc_hs__nand3_2 _49649_ (.A(_17264_),
    .B(_17574_),
    .C(_17577_),
    .Y(_17578_));
 sky130_as_sc_hs__or2_2 _49650_ (.A(\tholin_riscv.Iimm[0] ),
    .B(_17264_),
    .Y(_17579_));
 sky130_as_sc_hs__and2_2 _49651_ (.A(net508),
    .B(_17579_),
    .Y(_17580_));
 sky130_as_sc_hs__and2_2 _49652_ (.A(_17578_),
    .B(_17580_),
    .Y(_01364_));
 sky130_as_sc_hs__nor2_2 _49653_ (.A(_19683_),
    .B(_17572_),
    .Y(_17581_));
 sky130_as_sc_hs__inv_2 _49654_ (.Y(_17582_),
    .A(_17581_));
 sky130_as_sc_hs__nand3_2 _49655_ (.A(net1258),
    .B(_17404_),
    .C(_17581_),
    .Y(_17583_));
 sky130_as_sc_hs__and2_2 _49656_ (.A(net96),
    .B(_17582_),
    .Y(_17584_));
 sky130_as_sc_hs__or2_2 _49657_ (.A(_16370_),
    .B(_17584_),
    .Y(_17585_));
 sky130_as_sc_hs__nand3_2 _49659_ (.A(_17264_),
    .B(net1259),
    .C(_17586_),
    .Y(_17587_));
 sky130_as_sc_hs__and2_2 _49661_ (.A(net508),
    .B(_17588_),
    .Y(_17589_));
 sky130_as_sc_hs__and2_2 _49662_ (.A(_17587_),
    .B(_17589_),
    .Y(_01365_));
 sky130_as_sc_hs__and2_2 _49663_ (.A(\tholin_riscv.tmr1[21] ),
    .B(_17581_),
    .Y(_17590_));
 sky130_as_sc_hs__nand3_2 _49664_ (.A(net819),
    .B(_17404_),
    .C(_17590_),
    .Y(_17591_));
 sky130_as_sc_hs__nor2b_2 _49665_ (.A(_17590_),
    .Y(_17592_),
    .B(net96));
 sky130_as_sc_hs__or2_2 _49666_ (.A(_16370_),
    .B(_17592_),
    .Y(_17593_));
 sky130_as_sc_hs__nand3_2 _49668_ (.A(_17264_),
    .B(net820),
    .C(_17594_),
    .Y(_17595_));
 sky130_as_sc_hs__or2_2 _49669_ (.A(\tholin_riscv.Iimm[2] ),
    .B(_17264_),
    .Y(_17596_));
 sky130_as_sc_hs__and2_2 _49670_ (.A(net508),
    .B(_17596_),
    .Y(_17597_));
 sky130_as_sc_hs__and2_2 _49671_ (.A(net821),
    .B(_17597_),
    .Y(_01366_));
 sky130_as_sc_hs__nor2_2 _49673_ (.A(\tholin_riscv.tmr1[23] ),
    .B(_17598_),
    .Y(_17599_));
 sky130_as_sc_hs__and2_2 _49675_ (.A(net96),
    .B(_17598_),
    .Y(_17601_));
 sky130_as_sc_hs__or2_2 _49676_ (.A(_16370_),
    .B(_17601_),
    .Y(_17602_));
 sky130_as_sc_hs__nand3_2 _49678_ (.A(_17264_),
    .B(_17600_),
    .C(_17603_),
    .Y(_17604_));
 sky130_as_sc_hs__and2_2 _49680_ (.A(net507),
    .B(_17605_),
    .Y(_17606_));
 sky130_as_sc_hs__and2_2 _49681_ (.A(_17604_),
    .B(_17606_),
    .Y(_01367_));
 sky130_as_sc_hs__nor2_2 _49682_ (.A(_19689_),
    .B(_17598_),
    .Y(_17607_));
 sky130_as_sc_hs__nand3_2 _49683_ (.A(net1302),
    .B(net81),
    .C(_17607_),
    .Y(_17608_));
 sky130_as_sc_hs__nor2b_2 _49684_ (.A(_17607_),
    .Y(_17609_),
    .B(net96));
 sky130_as_sc_hs__or2_2 _49685_ (.A(_16370_),
    .B(_17609_),
    .Y(_17610_));
 sky130_as_sc_hs__nand3_2 _49687_ (.A(_17264_),
    .B(net1303),
    .C(_17611_),
    .Y(_17612_));
 sky130_as_sc_hs__and2_2 _49689_ (.A(net506),
    .B(_17613_),
    .Y(_17614_));
 sky130_as_sc_hs__and2_2 _49690_ (.A(_17612_),
    .B(_17614_),
    .Y(_01368_));
 sky130_as_sc_hs__and2_2 _49691_ (.A(\tholin_riscv.tmr1[24] ),
    .B(_17607_),
    .Y(_17615_));
 sky130_as_sc_hs__nand3_2 _49692_ (.A(net872),
    .B(net81),
    .C(_17615_),
    .Y(_17616_));
 sky130_as_sc_hs__nor2b_2 _49693_ (.A(_17615_),
    .Y(_17617_),
    .B(net96));
 sky130_as_sc_hs__or2_2 _49694_ (.A(_16370_),
    .B(_17617_),
    .Y(_17618_));
 sky130_as_sc_hs__nand3_2 _49696_ (.A(_17264_),
    .B(net873),
    .C(_17619_),
    .Y(_17620_));
 sky130_as_sc_hs__or2_2 _49697_ (.A(\tholin_riscv.Bimm[5] ),
    .B(_17264_),
    .Y(_17621_));
 sky130_as_sc_hs__and2_2 _49698_ (.A(net506),
    .B(_17621_),
    .Y(_17622_));
 sky130_as_sc_hs__and2_2 _49699_ (.A(net874),
    .B(_17622_),
    .Y(_01369_));
 sky130_as_sc_hs__nor2_2 _49701_ (.A(\tholin_riscv.tmr1[26] ),
    .B(_17623_),
    .Y(_17624_));
 sky130_as_sc_hs__and2_2 _49703_ (.A(net98),
    .B(_17623_),
    .Y(_17626_));
 sky130_as_sc_hs__or2_2 _49704_ (.A(_16370_),
    .B(_17626_),
    .Y(_17627_));
 sky130_as_sc_hs__nand3_2 _49706_ (.A(_17264_),
    .B(_17625_),
    .C(_17628_),
    .Y(_17629_));
 sky130_as_sc_hs__or2_2 _49707_ (.A(\tholin_riscv.Bimm[6] ),
    .B(_17264_),
    .Y(_17630_));
 sky130_as_sc_hs__and2_2 _49708_ (.A(net510),
    .B(_17630_),
    .Y(_17631_));
 sky130_as_sc_hs__and2_2 _49709_ (.A(_17629_),
    .B(_17631_),
    .Y(_01370_));
 sky130_as_sc_hs__nor2_2 _49710_ (.A(_19726_),
    .B(_17623_),
    .Y(_17632_));
 sky130_as_sc_hs__nand3_2 _49711_ (.A(net1163),
    .B(net81),
    .C(_17632_),
    .Y(_17633_));
 sky130_as_sc_hs__nor2b_2 _49712_ (.A(_17632_),
    .Y(_17634_),
    .B(net98));
 sky130_as_sc_hs__or2_2 _49713_ (.A(_16370_),
    .B(_17634_),
    .Y(_17635_));
 sky130_as_sc_hs__nand3_2 _49715_ (.A(_17264_),
    .B(net1164),
    .C(_17636_),
    .Y(_17637_));
 sky130_as_sc_hs__and2_2 _49717_ (.A(net510),
    .B(_17638_),
    .Y(_17639_));
 sky130_as_sc_hs__and2_2 _49718_ (.A(_17637_),
    .B(_17639_),
    .Y(_01371_));
 sky130_as_sc_hs__and2_2 _49719_ (.A(\tholin_riscv.tmr1[27] ),
    .B(_17632_),
    .Y(_17640_));
 sky130_as_sc_hs__nand3_2 _49720_ (.A(net952),
    .B(net81),
    .C(_17640_),
    .Y(_17641_));
 sky130_as_sc_hs__nor2b_2 _49721_ (.A(_17640_),
    .Y(_17642_),
    .B(net98));
 sky130_as_sc_hs__or2_2 _49722_ (.A(_16370_),
    .B(_17642_),
    .Y(_17643_));
 sky130_as_sc_hs__nand3_2 _49724_ (.A(_17264_),
    .B(net953),
    .C(_17644_),
    .Y(_17645_));
 sky130_as_sc_hs__and2_2 _49726_ (.A(net512),
    .B(_17646_),
    .Y(_17647_));
 sky130_as_sc_hs__and2_2 _49727_ (.A(net954),
    .B(_17647_),
    .Y(_01372_));
 sky130_as_sc_hs__nor2_2 _49729_ (.A(\tholin_riscv.tmr1[29] ),
    .B(_17648_),
    .Y(_17649_));
 sky130_as_sc_hs__and2_2 _49731_ (.A(net98),
    .B(_17648_),
    .Y(_17651_));
 sky130_as_sc_hs__or2_2 _49732_ (.A(_16370_),
    .B(_17651_),
    .Y(_17652_));
 sky130_as_sc_hs__nand3_2 _49734_ (.A(_17264_),
    .B(_17650_),
    .C(_17653_),
    .Y(_17654_));
 sky130_as_sc_hs__or2_2 _49735_ (.A(\tholin_riscv.Bimm[9] ),
    .B(_17264_),
    .Y(_17655_));
 sky130_as_sc_hs__and2_2 _49736_ (.A(net510),
    .B(_17655_),
    .Y(_17656_));
 sky130_as_sc_hs__and2_2 _49737_ (.A(_17654_),
    .B(_17656_),
    .Y(_01373_));
 sky130_as_sc_hs__nor2_2 _49738_ (.A(_19723_),
    .B(_17648_),
    .Y(_17657_));
 sky130_as_sc_hs__nand3_2 _49739_ (.A(net889),
    .B(net81),
    .C(_17657_),
    .Y(_17658_));
 sky130_as_sc_hs__nor2b_2 _49740_ (.A(_17657_),
    .Y(_17659_),
    .B(net98));
 sky130_as_sc_hs__or2_2 _49741_ (.A(_16370_),
    .B(_17659_),
    .Y(_17660_));
 sky130_as_sc_hs__nand3_2 _49743_ (.A(_17264_),
    .B(net890),
    .C(_17661_),
    .Y(_17662_));
 sky130_as_sc_hs__or2_2 _49744_ (.A(\tholin_riscv.Bimm[10] ),
    .B(_17264_),
    .Y(_17663_));
 sky130_as_sc_hs__and2_2 _49745_ (.A(net510),
    .B(_17663_),
    .Y(_17664_));
 sky130_as_sc_hs__and2_2 _49746_ (.A(_17662_),
    .B(_17664_),
    .Y(_01374_));
 sky130_as_sc_hs__nor2_2 _49748_ (.A(\tholin_riscv.tmr1[31] ),
    .B(_17665_),
    .Y(_17666_));
 sky130_as_sc_hs__and2_2 _49750_ (.A(net98),
    .B(_17665_),
    .Y(_17668_));
 sky130_as_sc_hs__or2_2 _49751_ (.A(_16370_),
    .B(_17668_),
    .Y(_17669_));
 sky130_as_sc_hs__nand3_2 _49753_ (.A(_17264_),
    .B(_17667_),
    .C(_17670_),
    .Y(_17671_));
 sky130_as_sc_hs__or2_2 _49754_ (.A(\tholin_riscv.Bimm[12] ),
    .B(_17264_),
    .Y(_17672_));
 sky130_as_sc_hs__and2_2 _49755_ (.A(net510),
    .B(_17672_),
    .Y(_17673_));
 sky130_as_sc_hs__and2_2 _49756_ (.A(_17671_),
    .B(_17673_),
    .Y(_01375_));
 sky130_as_sc_hs__nand3_2 _49759_ (.A(net506),
    .B(_17674_),
    .C(_17675_),
    .Y(_01376_));
 sky130_as_sc_hs__nand3_2 _49762_ (.A(net506),
    .B(_17676_),
    .C(_17677_),
    .Y(_01377_));
 sky130_as_sc_hs__nand3_2 _49765_ (.A(net506),
    .B(_17678_),
    .C(_17679_),
    .Y(_01378_));
 sky130_as_sc_hs__nand3_2 _49768_ (.A(net505),
    .B(_17680_),
    .C(_17681_),
    .Y(_01379_));
 sky130_as_sc_hs__nand3_2 _49771_ (.A(net505),
    .B(_17682_),
    .C(_17683_),
    .Y(_01380_));
 sky130_as_sc_hs__nand3_2 _49774_ (.A(net505),
    .B(_17684_),
    .C(_17685_),
    .Y(_01381_));
 sky130_as_sc_hs__nand3_2 _49777_ (.A(net505),
    .B(_17686_),
    .C(_17687_),
    .Y(_01382_));
 sky130_as_sc_hs__nand3_2 _49780_ (.A(net509),
    .B(_17688_),
    .C(_17689_),
    .Y(_01383_));
 sky130_as_sc_hs__nand3_2 _49783_ (.A(net512),
    .B(_17690_),
    .C(_17691_),
    .Y(_01384_));
 sky130_as_sc_hs__nand3_2 _49786_ (.A(net512),
    .B(_17692_),
    .C(_17693_),
    .Y(_01385_));
 sky130_as_sc_hs__nand3_2 _49789_ (.A(net512),
    .B(_17694_),
    .C(_17695_),
    .Y(_01386_));
 sky130_as_sc_hs__nand3_2 _49792_ (.A(net508),
    .B(_17696_),
    .C(_17697_),
    .Y(_01387_));
 sky130_as_sc_hs__nand3_2 _49795_ (.A(net508),
    .B(_17698_),
    .C(_17699_),
    .Y(_01388_));
 sky130_as_sc_hs__nand3_2 _49798_ (.A(net508),
    .B(_17700_),
    .C(_17701_),
    .Y(_01389_));
 sky130_as_sc_hs__nand3_2 _49801_ (.A(net507),
    .B(_17702_),
    .C(_17703_),
    .Y(_01390_));
 sky130_as_sc_hs__nand3_2 _49804_ (.A(net507),
    .B(_17704_),
    .C(_17705_),
    .Y(_01391_));
 sky130_as_sc_hs__nand3_2 _49807_ (.A(net507),
    .B(_17706_),
    .C(_17707_),
    .Y(_01392_));
 sky130_as_sc_hs__nand3_2 _49810_ (.A(net507),
    .B(_17708_),
    .C(_17709_),
    .Y(_01393_));
 sky130_as_sc_hs__nand3_2 _49813_ (.A(net507),
    .B(_17710_),
    .C(_17711_),
    .Y(_01394_));
 sky130_as_sc_hs__nand3_2 _49816_ (.A(net509),
    .B(_17712_),
    .C(_17713_),
    .Y(_01395_));
 sky130_as_sc_hs__nand3_2 _49819_ (.A(net508),
    .B(_17714_),
    .C(_17715_),
    .Y(_01396_));
 sky130_as_sc_hs__nand3_2 _49822_ (.A(net508),
    .B(_17716_),
    .C(_17717_),
    .Y(_01397_));
 sky130_as_sc_hs__nand3_2 _49825_ (.A(net508),
    .B(_17718_),
    .C(_17719_),
    .Y(_01398_));
 sky130_as_sc_hs__nand3_2 _49828_ (.A(net508),
    .B(_17720_),
    .C(_17721_),
    .Y(_01399_));
 sky130_as_sc_hs__nand3_2 _49831_ (.A(net506),
    .B(_17722_),
    .C(_17723_),
    .Y(_01400_));
 sky130_as_sc_hs__nand3_2 _49834_ (.A(net509),
    .B(_17724_),
    .C(_17725_),
    .Y(_01401_));
 sky130_as_sc_hs__nand3_2 _49837_ (.A(net510),
    .B(_17726_),
    .C(_17727_),
    .Y(_01402_));
 sky130_as_sc_hs__nand3_2 _49840_ (.A(net510),
    .B(_17728_),
    .C(_17729_),
    .Y(_01403_));
 sky130_as_sc_hs__nand3_2 _49843_ (.A(net512),
    .B(_17730_),
    .C(_17731_),
    .Y(_01404_));
 sky130_as_sc_hs__nand3_2 _49846_ (.A(net510),
    .B(_17732_),
    .C(_17733_),
    .Y(_01405_));
 sky130_as_sc_hs__nand3_2 _49849_ (.A(net509),
    .B(_17734_),
    .C(_17735_),
    .Y(_01406_));
 sky130_as_sc_hs__nand3_2 _49852_ (.A(net510),
    .B(_17736_),
    .C(_17737_),
    .Y(_01407_));
 sky130_as_sc_hs__nand3_2 _49855_ (.A(net491),
    .B(_17738_),
    .C(_17739_),
    .Y(_01408_));
 sky130_as_sc_hs__nand3_2 _49858_ (.A(net491),
    .B(_17740_),
    .C(_17741_),
    .Y(_01409_));
 sky130_as_sc_hs__nand3_2 _49861_ (.A(net491),
    .B(_17742_),
    .C(_17743_),
    .Y(_01410_));
 sky130_as_sc_hs__nand3_2 _49864_ (.A(net491),
    .B(_17744_),
    .C(_17745_),
    .Y(_01411_));
 sky130_as_sc_hs__nand3_2 _49867_ (.A(net490),
    .B(_17746_),
    .C(_17747_),
    .Y(_01412_));
 sky130_as_sc_hs__nand3_2 _49870_ (.A(net490),
    .B(_17748_),
    .C(_17749_),
    .Y(_01413_));
 sky130_as_sc_hs__nand3_2 _49873_ (.A(net490),
    .B(_17750_),
    .C(_17751_),
    .Y(_01414_));
 sky130_as_sc_hs__nand3_2 _49876_ (.A(net490),
    .B(_17752_),
    .C(_17753_),
    .Y(_01415_));
 sky130_as_sc_hs__nand3_2 _49879_ (.A(net510),
    .B(_17754_),
    .C(_17755_),
    .Y(_01416_));
 sky130_as_sc_hs__nand3_2 _49882_ (.A(net510),
    .B(_17756_),
    .C(_17757_),
    .Y(_01417_));
 sky130_as_sc_hs__nand3_2 _49885_ (.A(net506),
    .B(_17758_),
    .C(_17759_),
    .Y(_01418_));
 sky130_as_sc_hs__nand3_2 _49888_ (.A(net506),
    .B(_17760_),
    .C(_17761_),
    .Y(_01419_));
 sky130_as_sc_hs__nand3_2 _49891_ (.A(net506),
    .B(_17762_),
    .C(_17763_),
    .Y(_01420_));
 sky130_as_sc_hs__nand3_2 _49894_ (.A(net505),
    .B(_17764_),
    .C(_17765_),
    .Y(_01421_));
 sky130_as_sc_hs__nand3_2 _49897_ (.A(net492),
    .B(_17766_),
    .C(_17767_),
    .Y(_01422_));
 sky130_as_sc_hs__nand3_2 _49900_ (.A(net492),
    .B(_17768_),
    .C(_17769_),
    .Y(_01423_));
 sky130_as_sc_hs__nand3_2 _49903_ (.A(net505),
    .B(_17770_),
    .C(_17771_),
    .Y(_01424_));
 sky130_as_sc_hs__nand3_2 _49906_ (.A(net505),
    .B(_17772_),
    .C(_17773_),
    .Y(_01425_));
 sky130_as_sc_hs__nand3_2 _49909_ (.A(net505),
    .B(_17774_),
    .C(_17775_),
    .Y(_01426_));
 sky130_as_sc_hs__nand3_2 _49912_ (.A(net505),
    .B(_17776_),
    .C(_17777_),
    .Y(_01427_));
 sky130_as_sc_hs__nand3_2 _49915_ (.A(net491),
    .B(_17778_),
    .C(_17779_),
    .Y(_01428_));
 sky130_as_sc_hs__nand3_2 _49918_ (.A(net491),
    .B(_17780_),
    .C(_17781_),
    .Y(_01429_));
 sky130_as_sc_hs__nand3_2 _49921_ (.A(net491),
    .B(_17782_),
    .C(_17783_),
    .Y(_01430_));
 sky130_as_sc_hs__nand3_2 _49924_ (.A(net491),
    .B(_17784_),
    .C(_17785_),
    .Y(_01431_));
 sky130_as_sc_hs__nand3_2 _49927_ (.A(net491),
    .B(_17786_),
    .C(_17787_),
    .Y(_01432_));
 sky130_as_sc_hs__nand3_2 _49930_ (.A(net492),
    .B(_17788_),
    .C(_17789_),
    .Y(_01433_));
 sky130_as_sc_hs__nand3_2 _49933_ (.A(net493),
    .B(_17790_),
    .C(_17791_),
    .Y(_01434_));
 sky130_as_sc_hs__nand3_2 _49936_ (.A(net493),
    .B(_17792_),
    .C(_17793_),
    .Y(_01435_));
 sky130_as_sc_hs__nand3_2 _49939_ (.A(net492),
    .B(_17794_),
    .C(_17795_),
    .Y(_01436_));
 sky130_as_sc_hs__nand3_2 _49942_ (.A(net493),
    .B(_17796_),
    .C(_17797_),
    .Y(_01437_));
 sky130_as_sc_hs__nand3_2 _49945_ (.A(net493),
    .B(_17798_),
    .C(_17799_),
    .Y(_01438_));
 sky130_as_sc_hs__nand3_2 _49948_ (.A(net494),
    .B(_17800_),
    .C(_17801_),
    .Y(_01439_));
 sky130_as_sc_hs__or2_2 _49949_ (.A(net1185),
    .B(net103),
    .Y(_17802_));
 sky130_as_sc_hs__or2_2 _49950_ (.A(\tholin_riscv.instr[0] ),
    .B(_19962_),
    .Y(_17803_));
 sky130_as_sc_hs__and2_2 _49951_ (.A(net511),
    .B(net1186),
    .Y(_17804_));
 sky130_as_sc_hs__and2_2 _49952_ (.A(_17803_),
    .B(net1187),
    .Y(_01440_));
 sky130_as_sc_hs__or2_2 _49953_ (.A(net1376),
    .B(net104),
    .Y(_17805_));
 sky130_as_sc_hs__or2_2 _49954_ (.A(net1684),
    .B(_19962_),
    .Y(_17806_));
 sky130_as_sc_hs__and2_2 _49955_ (.A(net514),
    .B(net1377),
    .Y(_17807_));
 sky130_as_sc_hs__and2_2 _49956_ (.A(_17806_),
    .B(net1378),
    .Y(_01441_));
 sky130_as_sc_hs__or2_2 _49957_ (.A(net1392),
    .B(net104),
    .Y(_17808_));
 sky130_as_sc_hs__and2_2 _49959_ (.A(net514),
    .B(net1393),
    .Y(_17810_));
 sky130_as_sc_hs__and2_2 _49960_ (.A(_17809_),
    .B(net1394),
    .Y(_01442_));
 sky130_as_sc_hs__or2_2 _49961_ (.A(net1473),
    .B(net104),
    .Y(_17811_));
 sky130_as_sc_hs__and2_2 _49963_ (.A(net514),
    .B(net1474),
    .Y(_17813_));
 sky130_as_sc_hs__and2_2 _49964_ (.A(_17812_),
    .B(net1475),
    .Y(_01443_));
 sky130_as_sc_hs__or2_2 _49965_ (.A(net1506),
    .B(net104),
    .Y(_17814_));
 sky130_as_sc_hs__and2_2 _49967_ (.A(net514),
    .B(net1507),
    .Y(_17816_));
 sky130_as_sc_hs__and2_2 _49968_ (.A(_17815_),
    .B(net1508),
    .Y(_01444_));
 sky130_as_sc_hs__or2_2 _49969_ (.A(net1395),
    .B(net104),
    .Y(_17817_));
 sky130_as_sc_hs__and2_2 _49971_ (.A(net514),
    .B(net1396),
    .Y(_17819_));
 sky130_as_sc_hs__and2_2 _49972_ (.A(_17818_),
    .B(net1397),
    .Y(_01445_));
 sky130_as_sc_hs__or2_2 _49973_ (.A(net1490),
    .B(net104),
    .Y(_17820_));
 sky130_as_sc_hs__and2_2 _49975_ (.A(net512),
    .B(net1491),
    .Y(_17822_));
 sky130_as_sc_hs__and2_2 _49976_ (.A(_17821_),
    .B(net1492),
    .Y(_01446_));
 sky130_as_sc_hs__or2_2 _49977_ (.A(net1536),
    .B(net103),
    .Y(_17823_));
 sky130_as_sc_hs__or2_2 _49978_ (.A(\tholin_riscv.Bimm[11] ),
    .B(_19962_),
    .Y(_17824_));
 sky130_as_sc_hs__and2_2 _49979_ (.A(net512),
    .B(net1537),
    .Y(_17825_));
 sky130_as_sc_hs__and2_2 _49980_ (.A(_17824_),
    .B(net1538),
    .Y(_01447_));
 sky130_as_sc_hs__or2_2 _49981_ (.A(net1479),
    .B(net103),
    .Y(_17826_));
 sky130_as_sc_hs__or2_2 _49982_ (.A(net1260),
    .B(_19962_),
    .Y(_17827_));
 sky130_as_sc_hs__and2_2 _49983_ (.A(net513),
    .B(net1480),
    .Y(_17828_));
 sky130_as_sc_hs__and2_2 _49984_ (.A(_17827_),
    .B(net1481),
    .Y(_01448_));
 sky130_as_sc_hs__or2_2 _49985_ (.A(net1577),
    .B(net103),
    .Y(_17829_));
 sky130_as_sc_hs__or2_2 _49986_ (.A(net1168),
    .B(_19962_),
    .Y(_17830_));
 sky130_as_sc_hs__and2_2 _49987_ (.A(net513),
    .B(net1578),
    .Y(_17831_));
 sky130_as_sc_hs__and2_2 _49988_ (.A(_17830_),
    .B(net1579),
    .Y(_01449_));
 sky130_as_sc_hs__or2_2 _49989_ (.A(net1588),
    .B(net103),
    .Y(_17832_));
 sky130_as_sc_hs__or2_2 _49990_ (.A(net1374),
    .B(_19962_),
    .Y(_17833_));
 sky130_as_sc_hs__and2_2 _49991_ (.A(net513),
    .B(net1589),
    .Y(_17834_));
 sky130_as_sc_hs__and2_2 _49992_ (.A(_17833_),
    .B(_17834_),
    .Y(_01450_));
 sky130_as_sc_hs__or2_2 _49993_ (.A(net1493),
    .B(net103),
    .Y(_17835_));
 sky130_as_sc_hs__or2_2 _49994_ (.A(net1343),
    .B(_19962_),
    .Y(_17836_));
 sky130_as_sc_hs__and2_2 _49995_ (.A(net513),
    .B(net1494),
    .Y(_17837_));
 sky130_as_sc_hs__and2_2 _49996_ (.A(_17836_),
    .B(net1495),
    .Y(_01451_));
 sky130_as_sc_hs__nand3_2 _49999_ (.A(net513),
    .B(_17838_),
    .C(_17839_),
    .Y(_01452_));
 sky130_as_sc_hs__or2_2 _50000_ (.A(net1526),
    .B(net104),
    .Y(_17840_));
 sky130_as_sc_hs__and2_2 _50002_ (.A(net513),
    .B(net1527),
    .Y(_17842_));
 sky130_as_sc_hs__and2_2 _50003_ (.A(_17841_),
    .B(net1528),
    .Y(_01453_));
 sky130_as_sc_hs__or2_2 _50004_ (.A(net1383),
    .B(net104),
    .Y(_17843_));
 sky130_as_sc_hs__or2_2 _50005_ (.A(net1032),
    .B(_19962_),
    .Y(_17844_));
 sky130_as_sc_hs__and2_2 _50006_ (.A(net512),
    .B(net1384),
    .Y(_17845_));
 sky130_as_sc_hs__and2_2 _50007_ (.A(_17844_),
    .B(net1385),
    .Y(_01454_));
 sky130_as_sc_hs__or2_2 _50008_ (.A(net1431),
    .B(net104),
    .Y(_17846_));
 sky130_as_sc_hs__and2_2 _50010_ (.A(net514),
    .B(net1432),
    .Y(_17848_));
 sky130_as_sc_hs__and2_2 _50011_ (.A(_17847_),
    .B(net1433),
    .Y(_01455_));
 sky130_as_sc_hs__or2_2 _50012_ (.A(net1476),
    .B(net104),
    .Y(_17849_));
 sky130_as_sc_hs__and2_2 _50014_ (.A(net514),
    .B(net1477),
    .Y(_17851_));
 sky130_as_sc_hs__and2_2 _50015_ (.A(_17850_),
    .B(net1478),
    .Y(_01456_));
 sky130_as_sc_hs__or2_2 _50016_ (.A(net1349),
    .B(net104),
    .Y(_17852_));
 sky130_as_sc_hs__and2_2 _50018_ (.A(net514),
    .B(net1350),
    .Y(_17854_));
 sky130_as_sc_hs__and2_2 _50019_ (.A(_17853_),
    .B(net1351),
    .Y(_01457_));
 sky130_as_sc_hs__or2_2 _50020_ (.A(net1380),
    .B(net104),
    .Y(_17855_));
 sky130_as_sc_hs__and2_2 _50022_ (.A(net514),
    .B(net1381),
    .Y(_17857_));
 sky130_as_sc_hs__and2_2 _50023_ (.A(_17856_),
    .B(net1382),
    .Y(_01458_));
 sky130_as_sc_hs__or2_2 _50024_ (.A(net1419),
    .B(net104),
    .Y(_17858_));
 sky130_as_sc_hs__and2_2 _50026_ (.A(net512),
    .B(net1420),
    .Y(_17860_));
 sky130_as_sc_hs__and2_2 _50027_ (.A(_17859_),
    .B(net1421),
    .Y(_01459_));
 sky130_as_sc_hs__or2_2 _50028_ (.A(net1542),
    .B(net104),
    .Y(_17861_));
 sky130_as_sc_hs__or2_2 _50029_ (.A(\tholin_riscv.Iimm[0] ),
    .B(_19962_),
    .Y(_17862_));
 sky130_as_sc_hs__and2_2 _50030_ (.A(net512),
    .B(net1543),
    .Y(_17863_));
 sky130_as_sc_hs__and2_2 _50031_ (.A(_17862_),
    .B(net1544),
    .Y(_01460_));
 sky130_as_sc_hs__or2_2 _50032_ (.A(net1459),
    .B(net104),
    .Y(_17864_));
 sky130_as_sc_hs__and2_2 _50034_ (.A(net512),
    .B(net1460),
    .Y(_17866_));
 sky130_as_sc_hs__and2_2 _50035_ (.A(_17865_),
    .B(net1461),
    .Y(_01461_));
 sky130_as_sc_hs__or2_2 _50036_ (.A(net1361),
    .B(net103),
    .Y(_17867_));
 sky130_as_sc_hs__or2_2 _50037_ (.A(\tholin_riscv.Iimm[2] ),
    .B(_19962_),
    .Y(_17868_));
 sky130_as_sc_hs__and2_2 _50038_ (.A(net512),
    .B(net1362),
    .Y(_17869_));
 sky130_as_sc_hs__and2_2 _50039_ (.A(_17868_),
    .B(net1363),
    .Y(_01462_));
 sky130_as_sc_hs__or2_2 _50040_ (.A(net1509),
    .B(net103),
    .Y(_17870_));
 sky130_as_sc_hs__and2_2 _50042_ (.A(net512),
    .B(net1510),
    .Y(_17872_));
 sky130_as_sc_hs__and2_2 _50043_ (.A(_17871_),
    .B(net1511),
    .Y(_01463_));
 sky130_as_sc_hs__or2_2 _50044_ (.A(net1453),
    .B(net103),
    .Y(_17873_));
 sky130_as_sc_hs__and2_2 _50046_ (.A(net513),
    .B(net1454),
    .Y(_17875_));
 sky130_as_sc_hs__and2_2 _50047_ (.A(_17874_),
    .B(net1455),
    .Y(_01464_));
 sky130_as_sc_hs__or2_2 _50048_ (.A(net1415),
    .B(net103),
    .Y(_17876_));
 sky130_as_sc_hs__or2_2 _50049_ (.A(\tholin_riscv.Bimm[5] ),
    .B(_19962_),
    .Y(_17877_));
 sky130_as_sc_hs__and2_2 _50050_ (.A(net511),
    .B(net1416),
    .Y(_17878_));
 sky130_as_sc_hs__and2_2 _50051_ (.A(_17877_),
    .B(net1417),
    .Y(_01465_));
 sky130_as_sc_hs__or2_2 _50052_ (.A(net1580),
    .B(net103),
    .Y(_17879_));
 sky130_as_sc_hs__or2_2 _50053_ (.A(\tholin_riscv.Bimm[6] ),
    .B(_19962_),
    .Y(_17880_));
 sky130_as_sc_hs__and2_2 _50054_ (.A(net511),
    .B(net1581),
    .Y(_17881_));
 sky130_as_sc_hs__and2_2 _50055_ (.A(_17880_),
    .B(net1582),
    .Y(_01466_));
 sky130_as_sc_hs__or2_2 _50056_ (.A(net1441),
    .B(net103),
    .Y(_17882_));
 sky130_as_sc_hs__and2_2 _50058_ (.A(net511),
    .B(net1442),
    .Y(_17884_));
 sky130_as_sc_hs__and2_2 _50059_ (.A(_17883_),
    .B(net1443),
    .Y(_01467_));
 sky130_as_sc_hs__or2_2 _50060_ (.A(net1559),
    .B(net103),
    .Y(_17885_));
 sky130_as_sc_hs__and2_2 _50062_ (.A(net511),
    .B(net1560),
    .Y(_17887_));
 sky130_as_sc_hs__and2_2 _50063_ (.A(_17886_),
    .B(net1561),
    .Y(_01468_));
 sky130_as_sc_hs__or2_2 _50064_ (.A(net1555),
    .B(net103),
    .Y(_17888_));
 sky130_as_sc_hs__or2_2 _50065_ (.A(\tholin_riscv.Bimm[9] ),
    .B(_19962_),
    .Y(_17889_));
 sky130_as_sc_hs__and2_2 _50066_ (.A(net511),
    .B(net1556),
    .Y(_17890_));
 sky130_as_sc_hs__and2_2 _50067_ (.A(_17889_),
    .B(net1557),
    .Y(_01469_));
 sky130_as_sc_hs__or2_2 _50068_ (.A(net1469),
    .B(net103),
    .Y(_17891_));
 sky130_as_sc_hs__or2_2 _50069_ (.A(\tholin_riscv.Bimm[10] ),
    .B(_19962_),
    .Y(_17892_));
 sky130_as_sc_hs__and2_2 _50070_ (.A(net513),
    .B(net1470),
    .Y(_17893_));
 sky130_as_sc_hs__and2_2 _50071_ (.A(_17892_),
    .B(net1471),
    .Y(_01470_));
 sky130_as_sc_hs__or2_2 _50072_ (.A(net1502),
    .B(net103),
    .Y(_17894_));
 sky130_as_sc_hs__or2_2 _50073_ (.A(\tholin_riscv.Bimm[12] ),
    .B(_19962_),
    .Y(_17895_));
 sky130_as_sc_hs__and2_2 _50074_ (.A(net511),
    .B(net1503),
    .Y(_17896_));
 sky130_as_sc_hs__and2_2 _50075_ (.A(_17895_),
    .B(net1504),
    .Y(_01471_));
 sky130_as_sc_hs__and2_2 _50076_ (.A(_19901_),
    .B(_20000_),
    .Y(_17897_));
 sky130_as_sc_hs__or2_2 _50078_ (.A(net1131),
    .B(net95),
    .Y(_17899_));
 sky130_as_sc_hs__or2_2 _50079_ (.A(\tholin_riscv.instr[0] ),
    .B(_17898_),
    .Y(_17900_));
 sky130_as_sc_hs__and2_2 _50080_ (.A(net523),
    .B(net1132),
    .Y(_17901_));
 sky130_as_sc_hs__and2_2 _50081_ (.A(_17900_),
    .B(net1133),
    .Y(_01472_));
 sky130_as_sc_hs__or2_2 _50082_ (.A(net1462),
    .B(net95),
    .Y(_17902_));
 sky130_as_sc_hs__or2_2 _50083_ (.A(net1684),
    .B(_17898_),
    .Y(_17903_));
 sky130_as_sc_hs__and2_2 _50084_ (.A(net518),
    .B(net1463),
    .Y(_17904_));
 sky130_as_sc_hs__and2_2 _50085_ (.A(_17903_),
    .B(net1464),
    .Y(_01473_));
 sky130_as_sc_hs__or2_2 _50086_ (.A(net1499),
    .B(net95),
    .Y(_17905_));
 sky130_as_sc_hs__and2_2 _50088_ (.A(net523),
    .B(net1500),
    .Y(_17907_));
 sky130_as_sc_hs__and2_2 _50089_ (.A(_17906_),
    .B(net1501),
    .Y(_01474_));
 sky130_as_sc_hs__or2_2 _50090_ (.A(net1355),
    .B(net95),
    .Y(_17908_));
 sky130_as_sc_hs__and2_2 _50092_ (.A(net523),
    .B(net1356),
    .Y(_17910_));
 sky130_as_sc_hs__and2_2 _50093_ (.A(_17909_),
    .B(net1357),
    .Y(_01475_));
 sky130_as_sc_hs__or2_2 _50094_ (.A(net1450),
    .B(net95),
    .Y(_17911_));
 sky130_as_sc_hs__and2_2 _50096_ (.A(net518),
    .B(net1451),
    .Y(_17913_));
 sky130_as_sc_hs__and2_2 _50097_ (.A(_17912_),
    .B(net1452),
    .Y(_01476_));
 sky130_as_sc_hs__or2_2 _50098_ (.A(net1545),
    .B(net95),
    .Y(_17914_));
 sky130_as_sc_hs__and2_2 _50100_ (.A(net518),
    .B(net1546),
    .Y(_17916_));
 sky130_as_sc_hs__and2_2 _50101_ (.A(_17915_),
    .B(net1547),
    .Y(_01477_));
 sky130_as_sc_hs__or2_2 _50102_ (.A(net1444),
    .B(net94),
    .Y(_17917_));
 sky130_as_sc_hs__and2_2 _50104_ (.A(net518),
    .B(net1445),
    .Y(_17919_));
 sky130_as_sc_hs__and2_2 _50105_ (.A(_17918_),
    .B(net1446),
    .Y(_01478_));
 sky130_as_sc_hs__or2_2 _50106_ (.A(net1404),
    .B(net94),
    .Y(_17920_));
 sky130_as_sc_hs__or2_2 _50107_ (.A(\tholin_riscv.Bimm[11] ),
    .B(_17898_),
    .Y(_17921_));
 sky130_as_sc_hs__and2_2 _50108_ (.A(net522),
    .B(net1405),
    .Y(_17922_));
 sky130_as_sc_hs__and2_2 _50109_ (.A(_17921_),
    .B(net1406),
    .Y(_01479_));
 sky130_as_sc_hs__or2_2 _50110_ (.A(net1771),
    .B(net94),
    .Y(_17923_));
 sky130_as_sc_hs__or2_2 _50111_ (.A(net1260),
    .B(_17898_),
    .Y(_17924_));
 sky130_as_sc_hs__and2_2 _50112_ (.A(net522),
    .B(net1772),
    .Y(_17925_));
 sky130_as_sc_hs__and2_2 _50113_ (.A(net1261),
    .B(_17925_),
    .Y(_01480_));
 sky130_as_sc_hs__or2_2 _50114_ (.A(net1330),
    .B(net94),
    .Y(_17926_));
 sky130_as_sc_hs__or2_2 _50115_ (.A(net1168),
    .B(_17898_),
    .Y(_17927_));
 sky130_as_sc_hs__and2_2 _50116_ (.A(net522),
    .B(net1331),
    .Y(_17928_));
 sky130_as_sc_hs__and2_2 _50117_ (.A(_17927_),
    .B(net1332),
    .Y(_01481_));
 sky130_as_sc_hs__or2_2 _50118_ (.A(net1411),
    .B(net94),
    .Y(_17929_));
 sky130_as_sc_hs__or2_2 _50119_ (.A(net1374),
    .B(_17898_),
    .Y(_17930_));
 sky130_as_sc_hs__and2_2 _50120_ (.A(net518),
    .B(net1412),
    .Y(_17931_));
 sky130_as_sc_hs__and2_2 _50121_ (.A(_17930_),
    .B(net1413),
    .Y(_01482_));
 sky130_as_sc_hs__or2_2 _50122_ (.A(net1486),
    .B(net94),
    .Y(_17932_));
 sky130_as_sc_hs__or2_2 _50123_ (.A(net1343),
    .B(_17898_),
    .Y(_17933_));
 sky130_as_sc_hs__and2_2 _50124_ (.A(net518),
    .B(net1487),
    .Y(_17934_));
 sky130_as_sc_hs__and2_2 _50125_ (.A(_17933_),
    .B(net1488),
    .Y(_01483_));
 sky130_as_sc_hs__or2_2 _50126_ (.A(net1422),
    .B(net95),
    .Y(_17935_));
 sky130_as_sc_hs__and2_2 _50128_ (.A(net518),
    .B(net1423),
    .Y(_17937_));
 sky130_as_sc_hs__and2_2 _50129_ (.A(_17936_),
    .B(net1424),
    .Y(_01484_));
 sky130_as_sc_hs__or2_2 _50130_ (.A(net1438),
    .B(net95),
    .Y(_17938_));
 sky130_as_sc_hs__and2_2 _50132_ (.A(net523),
    .B(net1439),
    .Y(_17940_));
 sky130_as_sc_hs__and2_2 _50133_ (.A(_17939_),
    .B(net1440),
    .Y(_01485_));
 sky130_as_sc_hs__or2_2 _50134_ (.A(net1529),
    .B(net95),
    .Y(_17941_));
 sky130_as_sc_hs__or2_2 _50135_ (.A(net1032),
    .B(_17898_),
    .Y(_17942_));
 sky130_as_sc_hs__and2_2 _50136_ (.A(net518),
    .B(net1530),
    .Y(_17943_));
 sky130_as_sc_hs__and2_2 _50137_ (.A(_17942_),
    .B(net1531),
    .Y(_01486_));
 sky130_as_sc_hs__nand3_2 _50140_ (.A(net523),
    .B(_17944_),
    .C(_17945_),
    .Y(_01487_));
 sky130_as_sc_hs__or2_2 _50141_ (.A(net1346),
    .B(net95),
    .Y(_17946_));
 sky130_as_sc_hs__and2_2 _50143_ (.A(net523),
    .B(net1347),
    .Y(_17948_));
 sky130_as_sc_hs__and2_2 _50144_ (.A(_17947_),
    .B(net1348),
    .Y(_01488_));
 sky130_as_sc_hs__or2_2 _50145_ (.A(net1371),
    .B(net95),
    .Y(_17949_));
 sky130_as_sc_hs__and2_2 _50147_ (.A(net523),
    .B(net1372),
    .Y(_17951_));
 sky130_as_sc_hs__and2_2 _50148_ (.A(_17950_),
    .B(net1373),
    .Y(_01489_));
 sky130_as_sc_hs__or2_2 _50149_ (.A(net1466),
    .B(net95),
    .Y(_17952_));
 sky130_as_sc_hs__and2_2 _50151_ (.A(net523),
    .B(net1467),
    .Y(_17954_));
 sky130_as_sc_hs__and2_2 _50152_ (.A(_17953_),
    .B(net1468),
    .Y(_01490_));
 sky130_as_sc_hs__or2_2 _50153_ (.A(net1447),
    .B(net95),
    .Y(_17955_));
 sky130_as_sc_hs__and2_2 _50155_ (.A(net513),
    .B(net1448),
    .Y(_17957_));
 sky130_as_sc_hs__and2_2 _50156_ (.A(_17956_),
    .B(net1449),
    .Y(_01491_));
 sky130_as_sc_hs__or2_2 _50157_ (.A(net1521),
    .B(net95),
    .Y(_17958_));
 sky130_as_sc_hs__or2_2 _50158_ (.A(\tholin_riscv.Iimm[0] ),
    .B(_17898_),
    .Y(_17959_));
 sky130_as_sc_hs__and2_2 _50159_ (.A(net518),
    .B(net1522),
    .Y(_17960_));
 sky130_as_sc_hs__and2_2 _50160_ (.A(_17959_),
    .B(net1523),
    .Y(_01492_));
 sky130_as_sc_hs__or2_2 _50161_ (.A(net1515),
    .B(net95),
    .Y(_17961_));
 sky130_as_sc_hs__and2_2 _50163_ (.A(net513),
    .B(net1516),
    .Y(_17963_));
 sky130_as_sc_hs__and2_2 _50164_ (.A(_17962_),
    .B(net1517),
    .Y(_01493_));
 sky130_as_sc_hs__or2_2 _50165_ (.A(net1568),
    .B(net94),
    .Y(_17964_));
 sky130_as_sc_hs__or2_2 _50166_ (.A(\tholin_riscv.Iimm[2] ),
    .B(_17898_),
    .Y(_17965_));
 sky130_as_sc_hs__and2_2 _50167_ (.A(net518),
    .B(net1569),
    .Y(_17966_));
 sky130_as_sc_hs__and2_2 _50168_ (.A(_17965_),
    .B(net1570),
    .Y(_01494_));
 sky130_as_sc_hs__or2_2 _50169_ (.A(net1389),
    .B(net94),
    .Y(_17967_));
 sky130_as_sc_hs__and2_2 _50171_ (.A(net513),
    .B(net1390),
    .Y(_17969_));
 sky130_as_sc_hs__and2_2 _50172_ (.A(_17968_),
    .B(net1391),
    .Y(_01495_));
 sky130_as_sc_hs__or2_2 _50173_ (.A(net1352),
    .B(net94),
    .Y(_17970_));
 sky130_as_sc_hs__and2_2 _50175_ (.A(net513),
    .B(net1353),
    .Y(_17972_));
 sky130_as_sc_hs__and2_2 _50176_ (.A(_17971_),
    .B(net1354),
    .Y(_01496_));
 sky130_as_sc_hs__or2_2 _50177_ (.A(net1364),
    .B(net94),
    .Y(_17973_));
 sky130_as_sc_hs__or2_2 _50178_ (.A(\tholin_riscv.Bimm[5] ),
    .B(_17898_),
    .Y(_17974_));
 sky130_as_sc_hs__and2_2 _50179_ (.A(net517),
    .B(net1365),
    .Y(_17975_));
 sky130_as_sc_hs__and2_2 _50180_ (.A(_17974_),
    .B(net1366),
    .Y(_01497_));
 sky130_as_sc_hs__or2_2 _50181_ (.A(net1584),
    .B(net94),
    .Y(_17976_));
 sky130_as_sc_hs__or2_2 _50182_ (.A(net1781),
    .B(_17898_),
    .Y(_17977_));
 sky130_as_sc_hs__and2_2 _50183_ (.A(net517),
    .B(net1585),
    .Y(_17978_));
 sky130_as_sc_hs__and2_2 _50184_ (.A(_17977_),
    .B(net1586),
    .Y(_01498_));
 sky130_as_sc_hs__or2_2 _50185_ (.A(net1533),
    .B(net94),
    .Y(_17979_));
 sky130_as_sc_hs__and2_2 _50187_ (.A(net518),
    .B(net1534),
    .Y(_17981_));
 sky130_as_sc_hs__and2_2 _50188_ (.A(_17980_),
    .B(net1535),
    .Y(_01499_));
 sky130_as_sc_hs__or2_2 _50189_ (.A(net1368),
    .B(net94),
    .Y(_17982_));
 sky130_as_sc_hs__and2_2 _50191_ (.A(net517),
    .B(net1369),
    .Y(_17984_));
 sky130_as_sc_hs__and2_2 _50192_ (.A(_17983_),
    .B(net1370),
    .Y(_01500_));
 sky130_as_sc_hs__or2_2 _50193_ (.A(net1551),
    .B(net94),
    .Y(_17985_));
 sky130_as_sc_hs__or2_2 _50194_ (.A(net1779),
    .B(_17898_),
    .Y(_17986_));
 sky130_as_sc_hs__and2_2 _50195_ (.A(net517),
    .B(net1552),
    .Y(_17987_));
 sky130_as_sc_hs__and2_2 _50196_ (.A(_17986_),
    .B(net1553),
    .Y(_01501_));
 sky130_as_sc_hs__or2_2 _50197_ (.A(net1434),
    .B(net94),
    .Y(_17988_));
 sky130_as_sc_hs__or2_2 _50198_ (.A(\tholin_riscv.Bimm[10] ),
    .B(_17898_),
    .Y(_17989_));
 sky130_as_sc_hs__and2_2 _50199_ (.A(net522),
    .B(net1435),
    .Y(_17990_));
 sky130_as_sc_hs__and2_2 _50200_ (.A(_17989_),
    .B(net1436),
    .Y(_01502_));
 sky130_as_sc_hs__or2_2 _50201_ (.A(net1456),
    .B(net94),
    .Y(_17991_));
 sky130_as_sc_hs__or2_2 _50202_ (.A(net334),
    .B(_17898_),
    .Y(_17992_));
 sky130_as_sc_hs__and2_2 _50203_ (.A(net517),
    .B(net1457),
    .Y(_17993_));
 sky130_as_sc_hs__and2_2 _50204_ (.A(_17992_),
    .B(net1458),
    .Y(_01503_));
 sky130_as_sc_hs__and2_2 _50205_ (.A(_19901_),
    .B(_20028_),
    .Y(_17994_));
 sky130_as_sc_hs__nor2_2 _50210_ (.A(\tholin_riscv.tmr0_top[30] ),
    .B(_19695_),
    .Y(_17999_));
 sky130_as_sc_hs__nor2_2 _50211_ (.A(\tholin_riscv.tmr0_top[31] ),
    .B(_19694_),
    .Y(_18000_));
 sky130_as_sc_hs__nor2_2 _50212_ (.A(_17999_),
    .B(_18000_),
    .Y(_18001_));
 sky130_as_sc_hs__nor2_2 _50213_ (.A(\tholin_riscv.tmr0_top[29] ),
    .B(_19696_),
    .Y(_18002_));
 sky130_as_sc_hs__nor2_2 _50214_ (.A(\tholin_riscv.tmr0_top[28] ),
    .B(_19697_),
    .Y(_18003_));
 sky130_as_sc_hs__nor2_2 _50215_ (.A(_18002_),
    .B(_18003_),
    .Y(_18004_));
 sky130_as_sc_hs__nor2_2 _50216_ (.A(\tholin_riscv.tmr0_top[27] ),
    .B(_19698_),
    .Y(_18005_));
 sky130_as_sc_hs__nor2_2 _50217_ (.A(\tholin_riscv.tmr0_top[26] ),
    .B(_19699_),
    .Y(_18006_));
 sky130_as_sc_hs__nor2_2 _50218_ (.A(_18005_),
    .B(_18006_),
    .Y(_18007_));
 sky130_as_sc_hs__nor2_2 _50219_ (.A(\tholin_riscv.tmr0_top[24] ),
    .B(_19692_),
    .Y(_18008_));
 sky130_as_sc_hs__nor2_2 _50220_ (.A(\tholin_riscv.tmr0_top[25] ),
    .B(_19700_),
    .Y(_18009_));
 sky130_as_sc_hs__or2_2 _50221_ (.A(_18008_),
    .B(_18009_),
    .Y(_18010_));
 sky130_as_sc_hs__and2_2 _50224_ (.A(_18011_),
    .B(_18012_),
    .Y(_18013_));
 sky130_as_sc_hs__and2_2 _50229_ (.A(_18016_),
    .B(_18017_),
    .Y(_18018_));
 sky130_as_sc_hs__and2_2 _50234_ (.A(_18021_),
    .B(_18022_),
    .Y(_18023_));
 sky130_as_sc_hs__nor2_2 _50239_ (.A(\tholin_riscv.tmr0_top[22] ),
    .B(_19688_),
    .Y(_18028_));
 sky130_as_sc_hs__nor2_2 _50240_ (.A(\tholin_riscv.tmr0_top[23] ),
    .B(_19690_),
    .Y(_18029_));
 sky130_as_sc_hs__nor2_2 _50241_ (.A(_18028_),
    .B(_18029_),
    .Y(_18030_));
 sky130_as_sc_hs__nor2_2 _50242_ (.A(\tholin_riscv.tmr0_top[21] ),
    .B(_19686_),
    .Y(_18031_));
 sky130_as_sc_hs__nor2_2 _50243_ (.A(\tholin_riscv.tmr0_top[20] ),
    .B(_19684_),
    .Y(_18032_));
 sky130_as_sc_hs__nor2_2 _50244_ (.A(_18031_),
    .B(_18032_),
    .Y(_18033_));
 sky130_as_sc_hs__nor2_2 _50245_ (.A(\tholin_riscv.tmr0_top[19] ),
    .B(_19701_),
    .Y(_18034_));
 sky130_as_sc_hs__nor2_2 _50246_ (.A(\tholin_riscv.tmr0_top[18] ),
    .B(_19702_),
    .Y(_18035_));
 sky130_as_sc_hs__nor2_2 _50247_ (.A(_18034_),
    .B(_18035_),
    .Y(_18036_));
 sky130_as_sc_hs__nor2_2 _50248_ (.A(\tholin_riscv.tmr0_top[16] ),
    .B(_19704_),
    .Y(_18037_));
 sky130_as_sc_hs__nor2_2 _50249_ (.A(\tholin_riscv.tmr0_top[17] ),
    .B(_19703_),
    .Y(_18038_));
 sky130_as_sc_hs__or2_2 _50250_ (.A(_18037_),
    .B(_18038_),
    .Y(_18039_));
 sky130_as_sc_hs__and2_2 _50253_ (.A(_18040_),
    .B(_18041_),
    .Y(_18042_));
 sky130_as_sc_hs__and2_2 _50258_ (.A(_18045_),
    .B(_18046_),
    .Y(_18047_));
 sky130_as_sc_hs__and2_2 _50263_ (.A(_18050_),
    .B(_18051_),
    .Y(_18052_));
 sky130_as_sc_hs__nor2_2 _50267_ (.A(\tholin_riscv.tmr0_top[14] ),
    .B(_19706_),
    .Y(_18056_));
 sky130_as_sc_hs__nor2_2 _50268_ (.A(\tholin_riscv.tmr0_top[15] ),
    .B(_19705_),
    .Y(_18057_));
 sky130_as_sc_hs__or2_2 _50269_ (.A(_18056_),
    .B(_18057_),
    .Y(_18058_));
 sky130_as_sc_hs__or2_2 _50272_ (.A(\tholin_riscv.tmr0_top[13] ),
    .B(_19707_),
    .Y(_18061_));
 sky130_as_sc_hs__or2_2 _50273_ (.A(\tholin_riscv.tmr0_top[12] ),
    .B(_19708_),
    .Y(_18062_));
 sky130_as_sc_hs__nor2_2 _50275_ (.A(\tholin_riscv.tmr0_top[11] ),
    .B(_19709_),
    .Y(_18064_));
 sky130_as_sc_hs__nor2_2 _50276_ (.A(\tholin_riscv.tmr0_top[10] ),
    .B(_19710_),
    .Y(_18065_));
 sky130_as_sc_hs__or2_2 _50277_ (.A(_18064_),
    .B(_18065_),
    .Y(_18066_));
 sky130_as_sc_hs__or2_2 _50280_ (.A(\tholin_riscv.tmr0_top[8] ),
    .B(_19712_),
    .Y(_18069_));
 sky130_as_sc_hs__or2_2 _50281_ (.A(\tholin_riscv.tmr0_top[9] ),
    .B(_19711_),
    .Y(_18070_));
 sky130_as_sc_hs__or2_2 _50283_ (.A(\tholin_riscv.tmr0_top[1] ),
    .B(_19719_),
    .Y(_18072_));
 sky130_as_sc_hs__nand3_2 _50285_ (.A(\tholin_riscv.tmr0_top[0] ),
    .B(_19720_),
    .C(_18072_),
    .Y(_18074_));
 sky130_as_sc_hs__nand3_2 _50286_ (.A(_18071_),
    .B(_18073_),
    .C(_18074_),
    .Y(_18075_));
 sky130_as_sc_hs__or2_2 _50287_ (.A(\tholin_riscv.tmr0_top[3] ),
    .B(_19717_),
    .Y(_18076_));
 sky130_as_sc_hs__or2_2 _50288_ (.A(\tholin_riscv.tmr0_top[2] ),
    .B(_19718_),
    .Y(_18077_));
 sky130_as_sc_hs__nand3_2 _50289_ (.A(_18075_),
    .B(_18076_),
    .C(_18077_),
    .Y(_18078_));
 sky130_as_sc_hs__nand3_2 _50292_ (.A(_18078_),
    .B(_18079_),
    .C(_18080_),
    .Y(_18081_));
 sky130_as_sc_hs__or2_2 _50293_ (.A(\tholin_riscv.tmr0_top[5] ),
    .B(_19715_),
    .Y(_18082_));
 sky130_as_sc_hs__or2_2 _50294_ (.A(\tholin_riscv.tmr0_top[4] ),
    .B(_19716_),
    .Y(_18083_));
 sky130_as_sc_hs__nand3_2 _50295_ (.A(_18081_),
    .B(_18082_),
    .C(_18083_),
    .Y(_18084_));
 sky130_as_sc_hs__or2_2 _50296_ (.A(\tholin_riscv.tmr0_top[6] ),
    .B(_19714_),
    .Y(_18085_));
 sky130_as_sc_hs__and2_2 _50298_ (.A(_18085_),
    .B(_18086_),
    .Y(_18087_));
 sky130_as_sc_hs__and2_2 _50301_ (.A(_18088_),
    .B(_18089_),
    .Y(_18090_));
 sky130_as_sc_hs__nand3_2 _50302_ (.A(_18084_),
    .B(_18087_),
    .C(_18090_),
    .Y(_18091_));
 sky130_as_sc_hs__nand2b_2 _50303_ (.B(_18086_),
    .Y(_18092_),
    .A(_18085_));
 sky130_as_sc_hs__or2_2 _50304_ (.A(\tholin_riscv.tmr0_top[7] ),
    .B(_19713_),
    .Y(_18093_));
 sky130_as_sc_hs__nand3_2 _50305_ (.A(_18091_),
    .B(_18092_),
    .C(_18093_),
    .Y(_18094_));
 sky130_as_sc_hs__nand3_2 _50308_ (.A(_18069_),
    .B(_18070_),
    .C(_18096_),
    .Y(_18097_));
 sky130_as_sc_hs__nand3_2 _50311_ (.A(_18067_),
    .B(_18098_),
    .C(_18099_),
    .Y(_18100_));
 sky130_as_sc_hs__nor2_2 _50312_ (.A(_18066_),
    .B(_18100_),
    .Y(_18101_));
 sky130_as_sc_hs__nand3_2 _50316_ (.A(_18061_),
    .B(_18062_),
    .C(_18104_),
    .Y(_18105_));
 sky130_as_sc_hs__nand3_2 _50319_ (.A(_18059_),
    .B(_18106_),
    .C(_18107_),
    .Y(_18108_));
 sky130_as_sc_hs__nor2_2 _50320_ (.A(_18058_),
    .B(_18108_),
    .Y(_18109_));
 sky130_as_sc_hs__nand2b_2 _50323_ (.B(_18042_),
    .Y(_18112_),
    .A(_18039_));
 sky130_as_sc_hs__nor2_2 _50325_ (.A(_18112_),
    .B(_18113_),
    .Y(_18114_));
 sky130_as_sc_hs__nand3_2 _50327_ (.A(_18027_),
    .B(_18030_),
    .C(_18115_),
    .Y(_18116_));
 sky130_as_sc_hs__nor2_2 _50329_ (.A(_18116_),
    .B(_18117_),
    .Y(_18118_));
 sky130_as_sc_hs__nand3_2 _50330_ (.A(_18111_),
    .B(_18114_),
    .C(_18118_),
    .Y(_18119_));
 sky130_as_sc_hs__nand2b_2 _50332_ (.B(_18013_),
    .Y(_18121_),
    .A(_18010_));
 sky130_as_sc_hs__nor2_2 _50334_ (.A(_18121_),
    .B(_18122_),
    .Y(_18123_));
 sky130_as_sc_hs__nand3_2 _50336_ (.A(_17998_),
    .B(_18001_),
    .C(_18124_),
    .Y(_18125_));
 sky130_as_sc_hs__nor2_2 _50338_ (.A(_18125_),
    .B(_18126_),
    .Y(_18127_));
 sky130_as_sc_hs__nand3_2 _50339_ (.A(_18120_),
    .B(_18123_),
    .C(_18127_),
    .Y(_18128_));
 sky130_as_sc_hs__and2_2 _50340_ (.A(_18026_),
    .B(_18128_),
    .Y(_18129_));
 sky130_as_sc_hs__and2_2 _50341_ (.A(_19720_),
    .B(net93),
    .Y(_18130_));
 sky130_as_sc_hs__nor2_2 _50342_ (.A(_17260_),
    .B(_18130_),
    .Y(_18131_));
 sky130_as_sc_hs__nor2_2 _50343_ (.A(_17994_),
    .B(_18131_),
    .Y(_18132_));
 sky130_as_sc_hs__and2_2 _50346_ (.A(net493),
    .B(_18134_),
    .Y(_01504_));
 sky130_as_sc_hs__nor2b_2 _50347_ (.A(_17260_),
    .Y(_18135_),
    .B(net92));
 sky130_as_sc_hs__nand3_2 _50348_ (.A(_19719_),
    .B(net779),
    .C(net80),
    .Y(_18136_));
 sky130_as_sc_hs__or2_2 _50349_ (.A(_19719_),
    .B(_18131_),
    .Y(_18137_));
 sky130_as_sc_hs__nand3_2 _50350_ (.A(_17995_),
    .B(net780),
    .C(_18137_),
    .Y(_18138_));
 sky130_as_sc_hs__or2_2 _50351_ (.A(\tholin_riscv.instr[1] ),
    .B(_17995_),
    .Y(_18139_));
 sky130_as_sc_hs__and2_2 _50352_ (.A(net493),
    .B(_18139_),
    .Y(_18140_));
 sky130_as_sc_hs__and2_2 _50353_ (.A(net781),
    .B(_18140_),
    .Y(_01505_));
 sky130_as_sc_hs__nor2_2 _50355_ (.A(\tholin_riscv.tmr0[2] ),
    .B(_18141_),
    .Y(_18142_));
 sky130_as_sc_hs__and2_2 _50357_ (.A(net92),
    .B(_18141_),
    .Y(_18144_));
 sky130_as_sc_hs__or2_2 _50358_ (.A(_17260_),
    .B(_18144_),
    .Y(_18145_));
 sky130_as_sc_hs__nand3_2 _50360_ (.A(_17995_),
    .B(_18143_),
    .C(_18146_),
    .Y(_18147_));
 sky130_as_sc_hs__and2_2 _50362_ (.A(net491),
    .B(_18148_),
    .Y(_18149_));
 sky130_as_sc_hs__and2_2 _50363_ (.A(_18147_),
    .B(_18149_),
    .Y(_01506_));
 sky130_as_sc_hs__nor2_2 _50364_ (.A(_19718_),
    .B(_18141_),
    .Y(_18150_));
 sky130_as_sc_hs__inv_2 _50365_ (.Y(_18151_),
    .A(_18150_));
 sky130_as_sc_hs__nand3_2 _50366_ (.A(net1074),
    .B(net80),
    .C(_18150_),
    .Y(_18152_));
 sky130_as_sc_hs__and2_2 _50367_ (.A(net92),
    .B(_18151_),
    .Y(_18153_));
 sky130_as_sc_hs__or2_2 _50368_ (.A(_17260_),
    .B(_18153_),
    .Y(_18154_));
 sky130_as_sc_hs__nand3_2 _50370_ (.A(_17995_),
    .B(net1075),
    .C(_18155_),
    .Y(_18156_));
 sky130_as_sc_hs__and2_2 _50372_ (.A(net491),
    .B(_18157_),
    .Y(_18158_));
 sky130_as_sc_hs__and2_2 _50373_ (.A(_18156_),
    .B(_18158_),
    .Y(_01507_));
 sky130_as_sc_hs__and2_2 _50374_ (.A(\tholin_riscv.tmr0[3] ),
    .B(_18150_),
    .Y(_18159_));
 sky130_as_sc_hs__inv_2 _50375_ (.Y(_18160_),
    .A(_18159_));
 sky130_as_sc_hs__nand3_2 _50376_ (.A(net807),
    .B(net80),
    .C(_18159_),
    .Y(_18161_));
 sky130_as_sc_hs__and2_2 _50377_ (.A(net92),
    .B(_18160_),
    .Y(_18162_));
 sky130_as_sc_hs__or2_2 _50378_ (.A(_17260_),
    .B(_18162_),
    .Y(_18163_));
 sky130_as_sc_hs__nand3_2 _50380_ (.A(_17995_),
    .B(net808),
    .C(_18164_),
    .Y(_18165_));
 sky130_as_sc_hs__and2_2 _50382_ (.A(net490),
    .B(_18166_),
    .Y(_18167_));
 sky130_as_sc_hs__and2_2 _50383_ (.A(net809),
    .B(_18167_),
    .Y(_01508_));
 sky130_as_sc_hs__nor2_2 _50385_ (.A(\tholin_riscv.tmr0[5] ),
    .B(_18168_),
    .Y(_18169_));
 sky130_as_sc_hs__and2_2 _50387_ (.A(net92),
    .B(_18168_),
    .Y(_18171_));
 sky130_as_sc_hs__or2_2 _50388_ (.A(_17260_),
    .B(_18171_),
    .Y(_18172_));
 sky130_as_sc_hs__nand3_2 _50390_ (.A(_17995_),
    .B(_18170_),
    .C(_18173_),
    .Y(_18174_));
 sky130_as_sc_hs__and2_2 _50392_ (.A(net490),
    .B(_18175_),
    .Y(_18176_));
 sky130_as_sc_hs__and2_2 _50393_ (.A(_18174_),
    .B(_18176_),
    .Y(_01509_));
 sky130_as_sc_hs__nor2_2 _50394_ (.A(_19715_),
    .B(_18168_),
    .Y(_18177_));
 sky130_as_sc_hs__inv_2 _50395_ (.Y(_18178_),
    .A(_18177_));
 sky130_as_sc_hs__nand3_2 _50396_ (.A(net1083),
    .B(net80),
    .C(_18177_),
    .Y(_18179_));
 sky130_as_sc_hs__and2_2 _50397_ (.A(net92),
    .B(_18178_),
    .Y(_18180_));
 sky130_as_sc_hs__or2_2 _50398_ (.A(_17260_),
    .B(_18180_),
    .Y(_18181_));
 sky130_as_sc_hs__nand3_2 _50400_ (.A(_17995_),
    .B(net1084),
    .C(_18182_),
    .Y(_18183_));
 sky130_as_sc_hs__and2_2 _50402_ (.A(net492),
    .B(_18184_),
    .Y(_18185_));
 sky130_as_sc_hs__and2_2 _50403_ (.A(net1085),
    .B(_18185_),
    .Y(_01510_));
 sky130_as_sc_hs__and2_2 _50404_ (.A(\tholin_riscv.tmr0[6] ),
    .B(_18177_),
    .Y(_18186_));
 sky130_as_sc_hs__inv_2 _50405_ (.Y(_18187_),
    .A(_18186_));
 sky130_as_sc_hs__nand3_2 _50406_ (.A(net791),
    .B(net80),
    .C(_18186_),
    .Y(_18188_));
 sky130_as_sc_hs__and2_2 _50407_ (.A(net92),
    .B(_18187_),
    .Y(_18189_));
 sky130_as_sc_hs__or2_2 _50408_ (.A(_17260_),
    .B(_18189_),
    .Y(_18190_));
 sky130_as_sc_hs__nand3_2 _50410_ (.A(_17995_),
    .B(net792),
    .C(_18191_),
    .Y(_18192_));
 sky130_as_sc_hs__or2_2 _50411_ (.A(\tholin_riscv.Bimm[11] ),
    .B(_17995_),
    .Y(_18193_));
 sky130_as_sc_hs__and2_2 _50412_ (.A(net492),
    .B(_18193_),
    .Y(_18194_));
 sky130_as_sc_hs__and2_2 _50413_ (.A(net793),
    .B(_18194_),
    .Y(_01511_));
 sky130_as_sc_hs__nor2_2 _50415_ (.A(\tholin_riscv.tmr0[8] ),
    .B(_18195_),
    .Y(_18196_));
 sky130_as_sc_hs__and2_2 _50417_ (.A(net93),
    .B(_18195_),
    .Y(_18198_));
 sky130_as_sc_hs__or2_2 _50418_ (.A(_17260_),
    .B(_18198_),
    .Y(_18199_));
 sky130_as_sc_hs__nand3_2 _50420_ (.A(_17995_),
    .B(_18197_),
    .C(_18200_),
    .Y(_18201_));
 sky130_as_sc_hs__or2_2 _50421_ (.A(net1260),
    .B(_17995_),
    .Y(_18202_));
 sky130_as_sc_hs__and2_2 _50422_ (.A(net510),
    .B(_18202_),
    .Y(_18203_));
 sky130_as_sc_hs__and2_2 _50423_ (.A(_18201_),
    .B(_18203_),
    .Y(_01512_));
 sky130_as_sc_hs__nor2_2 _50424_ (.A(_19712_),
    .B(_18195_),
    .Y(_18204_));
 sky130_as_sc_hs__inv_2 _50425_ (.Y(_18205_),
    .A(_18204_));
 sky130_as_sc_hs__nand3_2 _50426_ (.A(net1101),
    .B(_18135_),
    .C(_18204_),
    .Y(_18206_));
 sky130_as_sc_hs__and2_2 _50427_ (.A(net93),
    .B(_18205_),
    .Y(_18207_));
 sky130_as_sc_hs__or2_2 _50428_ (.A(_17260_),
    .B(_18207_),
    .Y(_18208_));
 sky130_as_sc_hs__nand3_2 _50430_ (.A(_17995_),
    .B(net1102),
    .C(_18209_),
    .Y(_18210_));
 sky130_as_sc_hs__or2_2 _50431_ (.A(net1780),
    .B(_17995_),
    .Y(_18211_));
 sky130_as_sc_hs__and2_2 _50432_ (.A(net510),
    .B(_18211_),
    .Y(_18212_));
 sky130_as_sc_hs__and2_2 _50433_ (.A(_18210_),
    .B(_18212_),
    .Y(_01513_));
 sky130_as_sc_hs__and2_2 _50434_ (.A(\tholin_riscv.tmr0[9] ),
    .B(_18204_),
    .Y(_18213_));
 sky130_as_sc_hs__inv_2 _50435_ (.Y(_18214_),
    .A(_18213_));
 sky130_as_sc_hs__nand3_2 _50436_ (.A(net848),
    .B(_18135_),
    .C(_18213_),
    .Y(_18215_));
 sky130_as_sc_hs__and2_2 _50437_ (.A(net93),
    .B(_18214_),
    .Y(_18216_));
 sky130_as_sc_hs__or2_2 _50438_ (.A(_17260_),
    .B(_18216_),
    .Y(_18217_));
 sky130_as_sc_hs__nand3_2 _50440_ (.A(_17995_),
    .B(net849),
    .C(_18218_),
    .Y(_18219_));
 sky130_as_sc_hs__or2_2 _50441_ (.A(net1791),
    .B(_17995_),
    .Y(_18220_));
 sky130_as_sc_hs__and2_2 _50442_ (.A(net510),
    .B(_18220_),
    .Y(_18221_));
 sky130_as_sc_hs__and2_2 _50443_ (.A(net850),
    .B(_18221_),
    .Y(_01514_));
 sky130_as_sc_hs__nor2_2 _50445_ (.A(\tholin_riscv.tmr0[11] ),
    .B(_18222_),
    .Y(_18223_));
 sky130_as_sc_hs__and2_2 _50447_ (.A(_18129_),
    .B(_18222_),
    .Y(_18225_));
 sky130_as_sc_hs__or2_2 _50448_ (.A(_17260_),
    .B(_18225_),
    .Y(_18226_));
 sky130_as_sc_hs__nand3_2 _50450_ (.A(_17995_),
    .B(_18224_),
    .C(_18227_),
    .Y(_18228_));
 sky130_as_sc_hs__or2_2 _50451_ (.A(net1792),
    .B(_17995_),
    .Y(_18229_));
 sky130_as_sc_hs__and2_2 _50452_ (.A(net506),
    .B(_18229_),
    .Y(_18230_));
 sky130_as_sc_hs__and2_2 _50453_ (.A(_18228_),
    .B(_18230_),
    .Y(_01515_));
 sky130_as_sc_hs__nor2_2 _50454_ (.A(_19709_),
    .B(_18222_),
    .Y(_18231_));
 sky130_as_sc_hs__inv_2 _50455_ (.Y(_18232_),
    .A(_18231_));
 sky130_as_sc_hs__nand3_2 _50456_ (.A(net1171),
    .B(_18135_),
    .C(_18231_),
    .Y(_18233_));
 sky130_as_sc_hs__and2_2 _50457_ (.A(net92),
    .B(_18232_),
    .Y(_18234_));
 sky130_as_sc_hs__or2_2 _50458_ (.A(_17260_),
    .B(_18234_),
    .Y(_18235_));
 sky130_as_sc_hs__nand3_2 _50460_ (.A(_17995_),
    .B(net1172),
    .C(_18236_),
    .Y(_18237_));
 sky130_as_sc_hs__and2_2 _50462_ (.A(net506),
    .B(_18238_),
    .Y(_18239_));
 sky130_as_sc_hs__and2_2 _50463_ (.A(_18237_),
    .B(_18239_),
    .Y(_01516_));
 sky130_as_sc_hs__and2_2 _50464_ (.A(\tholin_riscv.tmr0[12] ),
    .B(_18231_),
    .Y(_18240_));
 sky130_as_sc_hs__inv_2 _50465_ (.Y(_18241_),
    .A(_18240_));
 sky130_as_sc_hs__nand3_2 _50466_ (.A(net795),
    .B(net80),
    .C(_18240_),
    .Y(_18242_));
 sky130_as_sc_hs__and2_2 _50467_ (.A(net92),
    .B(_18241_),
    .Y(_18243_));
 sky130_as_sc_hs__or2_2 _50468_ (.A(_17260_),
    .B(_18243_),
    .Y(_18244_));
 sky130_as_sc_hs__nand3_2 _50470_ (.A(_17995_),
    .B(net796),
    .C(_18245_),
    .Y(_18246_));
 sky130_as_sc_hs__and2_2 _50472_ (.A(net505),
    .B(_18247_),
    .Y(_18248_));
 sky130_as_sc_hs__and2_2 _50473_ (.A(net797),
    .B(_18248_),
    .Y(_01517_));
 sky130_as_sc_hs__nor2_2 _50475_ (.A(\tholin_riscv.tmr0[14] ),
    .B(_18249_),
    .Y(_18250_));
 sky130_as_sc_hs__and2_2 _50477_ (.A(net92),
    .B(_18249_),
    .Y(_18252_));
 sky130_as_sc_hs__or2_2 _50478_ (.A(_17260_),
    .B(_18252_),
    .Y(_18253_));
 sky130_as_sc_hs__nand3_2 _50480_ (.A(_17995_),
    .B(_18251_),
    .C(_18254_),
    .Y(_18255_));
 sky130_as_sc_hs__or2_2 _50481_ (.A(net1796),
    .B(_17995_),
    .Y(_18256_));
 sky130_as_sc_hs__and2_2 _50482_ (.A(net492),
    .B(_18256_),
    .Y(_18257_));
 sky130_as_sc_hs__and2_2 _50483_ (.A(_18255_),
    .B(_18257_),
    .Y(_01518_));
 sky130_as_sc_hs__nor2_2 _50484_ (.A(_19706_),
    .B(_18249_),
    .Y(_18258_));
 sky130_as_sc_hs__inv_2 _50485_ (.Y(_18259_),
    .A(_18258_));
 sky130_as_sc_hs__nand3_2 _50486_ (.A(net1212),
    .B(net80),
    .C(_18258_),
    .Y(_18260_));
 sky130_as_sc_hs__and2_2 _50487_ (.A(net93),
    .B(_18259_),
    .Y(_18261_));
 sky130_as_sc_hs__or2_2 _50488_ (.A(_17260_),
    .B(_18261_),
    .Y(_18262_));
 sky130_as_sc_hs__nand3_2 _50490_ (.A(_17995_),
    .B(net1213),
    .C(_18263_),
    .Y(_18264_));
 sky130_as_sc_hs__and2_2 _50492_ (.A(net492),
    .B(_18265_),
    .Y(_18266_));
 sky130_as_sc_hs__and2_2 _50493_ (.A(_18264_),
    .B(_18266_),
    .Y(_01519_));
 sky130_as_sc_hs__and2_2 _50494_ (.A(\tholin_riscv.tmr0[15] ),
    .B(_18258_),
    .Y(_18267_));
 sky130_as_sc_hs__inv_2 _50495_ (.Y(_18268_),
    .A(_18267_));
 sky130_as_sc_hs__nand3_2 _50496_ (.A(net876),
    .B(net80),
    .C(_18267_),
    .Y(_18269_));
 sky130_as_sc_hs__and2_2 _50497_ (.A(net92),
    .B(_18268_),
    .Y(_18270_));
 sky130_as_sc_hs__or2_2 _50498_ (.A(_17260_),
    .B(_18270_),
    .Y(_18271_));
 sky130_as_sc_hs__nand3_2 _50500_ (.A(_17995_),
    .B(net877),
    .C(_18272_),
    .Y(_18273_));
 sky130_as_sc_hs__and2_2 _50502_ (.A(net505),
    .B(_18274_),
    .Y(_18275_));
 sky130_as_sc_hs__and2_2 _50503_ (.A(net878),
    .B(_18275_),
    .Y(_01520_));
 sky130_as_sc_hs__nor2_2 _50505_ (.A(\tholin_riscv.tmr0[17] ),
    .B(_18276_),
    .Y(_18277_));
 sky130_as_sc_hs__and2_2 _50507_ (.A(net93),
    .B(_18276_),
    .Y(_18279_));
 sky130_as_sc_hs__or2_2 _50508_ (.A(_17260_),
    .B(_18279_),
    .Y(_18280_));
 sky130_as_sc_hs__nand3_2 _50510_ (.A(_17995_),
    .B(_18278_),
    .C(_18281_),
    .Y(_18282_));
 sky130_as_sc_hs__and2_2 _50512_ (.A(net505),
    .B(_18283_),
    .Y(_18284_));
 sky130_as_sc_hs__and2_2 _50513_ (.A(_18282_),
    .B(_18284_),
    .Y(_01521_));
 sky130_as_sc_hs__nor2_2 _50514_ (.A(_19703_),
    .B(_18276_),
    .Y(_18285_));
 sky130_as_sc_hs__inv_2 _50515_ (.Y(_18286_),
    .A(_18285_));
 sky130_as_sc_hs__nand3_2 _50516_ (.A(net1327),
    .B(net80),
    .C(_18285_),
    .Y(_18287_));
 sky130_as_sc_hs__and2_2 _50517_ (.A(net92),
    .B(_18286_),
    .Y(_18288_));
 sky130_as_sc_hs__or2_2 _50518_ (.A(_17260_),
    .B(_18288_),
    .Y(_18289_));
 sky130_as_sc_hs__nand3_2 _50520_ (.A(_17995_),
    .B(net1328),
    .C(_18290_),
    .Y(_18291_));
 sky130_as_sc_hs__and2_2 _50522_ (.A(net505),
    .B(_18292_),
    .Y(_18293_));
 sky130_as_sc_hs__and2_2 _50523_ (.A(net1329),
    .B(_18293_),
    .Y(_01522_));
 sky130_as_sc_hs__and2_2 _50524_ (.A(\tholin_riscv.tmr0[18] ),
    .B(_18285_),
    .Y(_18294_));
 sky130_as_sc_hs__inv_2 _50525_ (.Y(_18295_),
    .A(_18294_));
 sky130_as_sc_hs__nand3_2 _50526_ (.A(net836),
    .B(net80),
    .C(_18294_),
    .Y(_18296_));
 sky130_as_sc_hs__and2_2 _50527_ (.A(net92),
    .B(_18295_),
    .Y(_18297_));
 sky130_as_sc_hs__or2_2 _50528_ (.A(_17260_),
    .B(_18297_),
    .Y(_18298_));
 sky130_as_sc_hs__nand3_2 _50530_ (.A(_17995_),
    .B(net837),
    .C(_18299_),
    .Y(_18300_));
 sky130_as_sc_hs__and2_2 _50532_ (.A(net509),
    .B(_18301_),
    .Y(_18302_));
 sky130_as_sc_hs__and2_2 _50533_ (.A(net838),
    .B(_18302_),
    .Y(_01523_));
 sky130_as_sc_hs__nor2_2 _50535_ (.A(\tholin_riscv.tmr0[20] ),
    .B(_18303_),
    .Y(_18304_));
 sky130_as_sc_hs__and2_2 _50537_ (.A(net93),
    .B(_18303_),
    .Y(_18306_));
 sky130_as_sc_hs__or2_2 _50538_ (.A(_17260_),
    .B(_18306_),
    .Y(_18307_));
 sky130_as_sc_hs__nand3_2 _50540_ (.A(_17995_),
    .B(_18305_),
    .C(_18308_),
    .Y(_18309_));
 sky130_as_sc_hs__or2_2 _50541_ (.A(\tholin_riscv.Iimm[0] ),
    .B(_17995_),
    .Y(_18310_));
 sky130_as_sc_hs__and2_2 _50542_ (.A(net492),
    .B(_18310_),
    .Y(_18311_));
 sky130_as_sc_hs__and2_2 _50543_ (.A(_18309_),
    .B(_18311_),
    .Y(_01524_));
 sky130_as_sc_hs__nor2_2 _50544_ (.A(_19684_),
    .B(_18303_),
    .Y(_18312_));
 sky130_as_sc_hs__inv_2 _50545_ (.Y(_18313_),
    .A(_18312_));
 sky130_as_sc_hs__nand3_2 _50546_ (.A(net1287),
    .B(_18135_),
    .C(_18312_),
    .Y(_18314_));
 sky130_as_sc_hs__and2_2 _50547_ (.A(net93),
    .B(_18313_),
    .Y(_18315_));
 sky130_as_sc_hs__or2_2 _50548_ (.A(_17260_),
    .B(_18315_),
    .Y(_18316_));
 sky130_as_sc_hs__nand3_2 _50550_ (.A(_17995_),
    .B(net1288),
    .C(_18317_),
    .Y(_18318_));
 sky130_as_sc_hs__and2_2 _50552_ (.A(net492),
    .B(_18319_),
    .Y(_18320_));
 sky130_as_sc_hs__and2_2 _50553_ (.A(_18318_),
    .B(_18320_),
    .Y(_01525_));
 sky130_as_sc_hs__and2_2 _50554_ (.A(\tholin_riscv.tmr0[21] ),
    .B(_18312_),
    .Y(_18321_));
 sky130_as_sc_hs__nand3_2 _50555_ (.A(net972),
    .B(net80),
    .C(_18321_),
    .Y(_18322_));
 sky130_as_sc_hs__nor2b_2 _50556_ (.A(_18321_),
    .Y(_18323_),
    .B(net92));
 sky130_as_sc_hs__or2_2 _50557_ (.A(_17260_),
    .B(_18323_),
    .Y(_18324_));
 sky130_as_sc_hs__nand3_2 _50559_ (.A(_17995_),
    .B(net973),
    .C(_18325_),
    .Y(_18326_));
 sky130_as_sc_hs__or2_2 _50560_ (.A(\tholin_riscv.Iimm[2] ),
    .B(_17995_),
    .Y(_18327_));
 sky130_as_sc_hs__and2_2 _50561_ (.A(net492),
    .B(_18327_),
    .Y(_18328_));
 sky130_as_sc_hs__and2_2 _50562_ (.A(net974),
    .B(_18328_),
    .Y(_01526_));
 sky130_as_sc_hs__nor2_2 _50564_ (.A(\tholin_riscv.tmr0[23] ),
    .B(_18329_),
    .Y(_18330_));
 sky130_as_sc_hs__and2_2 _50566_ (.A(net92),
    .B(_18329_),
    .Y(_18332_));
 sky130_as_sc_hs__or2_2 _50567_ (.A(_17260_),
    .B(_18332_),
    .Y(_18333_));
 sky130_as_sc_hs__nand3_2 _50569_ (.A(_17995_),
    .B(_18331_),
    .C(_18334_),
    .Y(_18335_));
 sky130_as_sc_hs__and2_2 _50571_ (.A(net492),
    .B(_18336_),
    .Y(_18337_));
 sky130_as_sc_hs__and2_2 _50572_ (.A(_18335_),
    .B(_18337_),
    .Y(_01527_));
 sky130_as_sc_hs__nor2_2 _50573_ (.A(_19690_),
    .B(_18329_),
    .Y(_18338_));
 sky130_as_sc_hs__nand3_2 _50574_ (.A(net1324),
    .B(net80),
    .C(_18338_),
    .Y(_18339_));
 sky130_as_sc_hs__nor2b_2 _50575_ (.A(_18338_),
    .Y(_18340_),
    .B(net93));
 sky130_as_sc_hs__or2_2 _50576_ (.A(_17260_),
    .B(_18340_),
    .Y(_18341_));
 sky130_as_sc_hs__nand3_2 _50578_ (.A(_17995_),
    .B(net1325),
    .C(_18342_),
    .Y(_18343_));
 sky130_as_sc_hs__and2_2 _50580_ (.A(net506),
    .B(_18344_),
    .Y(_18345_));
 sky130_as_sc_hs__and2_2 _50581_ (.A(_18343_),
    .B(_18345_),
    .Y(_01528_));
 sky130_as_sc_hs__and2_2 _50582_ (.A(\tholin_riscv.tmr0[24] ),
    .B(_18338_),
    .Y(_18346_));
 sky130_as_sc_hs__nand3_2 _50583_ (.A(net827),
    .B(net80),
    .C(_18346_),
    .Y(_18347_));
 sky130_as_sc_hs__nor2b_2 _50584_ (.A(_18346_),
    .Y(_18348_),
    .B(net92));
 sky130_as_sc_hs__or2_2 _50585_ (.A(_17260_),
    .B(_18348_),
    .Y(_18349_));
 sky130_as_sc_hs__nand3_2 _50587_ (.A(_17995_),
    .B(net828),
    .C(_18350_),
    .Y(_18351_));
 sky130_as_sc_hs__or2_2 _50588_ (.A(\tholin_riscv.Bimm[5] ),
    .B(_17995_),
    .Y(_18352_));
 sky130_as_sc_hs__and2_2 _50589_ (.A(net506),
    .B(_18352_),
    .Y(_18353_));
 sky130_as_sc_hs__and2_2 _50590_ (.A(net829),
    .B(_18353_),
    .Y(_01529_));
 sky130_as_sc_hs__nor2_2 _50592_ (.A(\tholin_riscv.tmr0[26] ),
    .B(_18354_),
    .Y(_18355_));
 sky130_as_sc_hs__and2_2 _50594_ (.A(net93),
    .B(_18354_),
    .Y(_18357_));
 sky130_as_sc_hs__or2_2 _50595_ (.A(_17260_),
    .B(_18357_),
    .Y(_18358_));
 sky130_as_sc_hs__nand3_2 _50597_ (.A(_17995_),
    .B(_18356_),
    .C(_18359_),
    .Y(_18360_));
 sky130_as_sc_hs__or2_2 _50598_ (.A(\tholin_riscv.Bimm[6] ),
    .B(_17995_),
    .Y(_18361_));
 sky130_as_sc_hs__and2_2 _50599_ (.A(net494),
    .B(_18361_),
    .Y(_18362_));
 sky130_as_sc_hs__and2_2 _50600_ (.A(_18360_),
    .B(_18362_),
    .Y(_01530_));
 sky130_as_sc_hs__nor2_2 _50601_ (.A(_19699_),
    .B(_18354_),
    .Y(_18363_));
 sky130_as_sc_hs__nand3_2 _50602_ (.A(net1199),
    .B(net80),
    .C(_18363_),
    .Y(_18364_));
 sky130_as_sc_hs__nor2b_2 _50603_ (.A(_18363_),
    .Y(_18365_),
    .B(net93));
 sky130_as_sc_hs__or2_2 _50604_ (.A(_17260_),
    .B(_18365_),
    .Y(_18366_));
 sky130_as_sc_hs__nand3_2 _50606_ (.A(_17995_),
    .B(net1200),
    .C(_18367_),
    .Y(_18368_));
 sky130_as_sc_hs__and2_2 _50608_ (.A(net494),
    .B(_18369_),
    .Y(_18370_));
 sky130_as_sc_hs__and2_2 _50609_ (.A(_18368_),
    .B(_18370_),
    .Y(_01531_));
 sky130_as_sc_hs__and2_2 _50610_ (.A(\tholin_riscv.tmr0[27] ),
    .B(_18363_),
    .Y(_18371_));
 sky130_as_sc_hs__nand3_2 _50611_ (.A(net924),
    .B(net80),
    .C(_18371_),
    .Y(_18372_));
 sky130_as_sc_hs__nor2b_2 _50612_ (.A(_18371_),
    .Y(_18373_),
    .B(net93));
 sky130_as_sc_hs__or2_2 _50613_ (.A(_17260_),
    .B(_18373_),
    .Y(_18374_));
 sky130_as_sc_hs__nand3_2 _50615_ (.A(_17995_),
    .B(net925),
    .C(_18375_),
    .Y(_18376_));
 sky130_as_sc_hs__and2_2 _50617_ (.A(net492),
    .B(_18377_),
    .Y(_18378_));
 sky130_as_sc_hs__and2_2 _50618_ (.A(net926),
    .B(_18378_),
    .Y(_01532_));
 sky130_as_sc_hs__nor2_2 _50620_ (.A(\tholin_riscv.tmr0[29] ),
    .B(_18379_),
    .Y(_18380_));
 sky130_as_sc_hs__and2_2 _50622_ (.A(net93),
    .B(_18379_),
    .Y(_18382_));
 sky130_as_sc_hs__or2_2 _50623_ (.A(_17260_),
    .B(_18382_),
    .Y(_18383_));
 sky130_as_sc_hs__nand3_2 _50625_ (.A(_17995_),
    .B(_18381_),
    .C(_18384_),
    .Y(_18385_));
 sky130_as_sc_hs__or2_2 _50626_ (.A(\tholin_riscv.Bimm[9] ),
    .B(_17995_),
    .Y(_18386_));
 sky130_as_sc_hs__and2_2 _50627_ (.A(net494),
    .B(_18386_),
    .Y(_18387_));
 sky130_as_sc_hs__and2_2 _50628_ (.A(_18385_),
    .B(_18387_),
    .Y(_01533_));
 sky130_as_sc_hs__nor2_2 _50629_ (.A(_19696_),
    .B(_18379_),
    .Y(_18388_));
 sky130_as_sc_hs__nand3_2 _50630_ (.A(net1043),
    .B(net80),
    .C(_18388_),
    .Y(_18389_));
 sky130_as_sc_hs__nor2b_2 _50631_ (.A(_18388_),
    .Y(_18390_),
    .B(net93));
 sky130_as_sc_hs__or2_2 _50632_ (.A(_17260_),
    .B(_18390_),
    .Y(_18391_));
 sky130_as_sc_hs__nand3_2 _50634_ (.A(_17995_),
    .B(net1044),
    .C(_18392_),
    .Y(_18393_));
 sky130_as_sc_hs__or2_2 _50635_ (.A(\tholin_riscv.Bimm[10] ),
    .B(_17995_),
    .Y(_18394_));
 sky130_as_sc_hs__and2_2 _50636_ (.A(net510),
    .B(_18394_),
    .Y(_18395_));
 sky130_as_sc_hs__and2_2 _50637_ (.A(_18393_),
    .B(_18395_),
    .Y(_01534_));
 sky130_as_sc_hs__nor2_2 _50639_ (.A(\tholin_riscv.tmr0[31] ),
    .B(_18396_),
    .Y(_18397_));
 sky130_as_sc_hs__and2_2 _50641_ (.A(net93),
    .B(_18396_),
    .Y(_18399_));
 sky130_as_sc_hs__or2_2 _50642_ (.A(_17260_),
    .B(_18399_),
    .Y(_18400_));
 sky130_as_sc_hs__nand3_2 _50644_ (.A(_17995_),
    .B(_18398_),
    .C(_18401_),
    .Y(_18402_));
 sky130_as_sc_hs__or2_2 _50645_ (.A(\tholin_riscv.Bimm[12] ),
    .B(_17995_),
    .Y(_18403_));
 sky130_as_sc_hs__and2_2 _50646_ (.A(net510),
    .B(_18403_),
    .Y(_18404_));
 sky130_as_sc_hs__and2_2 _50647_ (.A(_18402_),
    .B(_18404_),
    .Y(_01535_));
 sky130_as_sc_hs__nand3_2 _50650_ (.A(net487),
    .B(_16398_),
    .C(_18406_),
    .Y(_18407_));
 sky130_as_sc_hs__and2_2 _50653_ (.A(_18408_),
    .B(_18409_),
    .Y(_18410_));
 sky130_as_sc_hs__or2_2 _50654_ (.A(net146),
    .B(_18410_),
    .Y(_18411_));
 sky130_as_sc_hs__and2_2 _50659_ (.A(_18413_),
    .B(_18414_),
    .Y(_18415_));
 sky130_as_sc_hs__or2_2 _50660_ (.A(net147),
    .B(_18415_),
    .Y(_18416_));
 sky130_as_sc_hs__and2_2 _50665_ (.A(_18418_),
    .B(_18419_),
    .Y(_18420_));
 sky130_as_sc_hs__or2_2 _50666_ (.A(net146),
    .B(_18420_),
    .Y(_18421_));
 sky130_as_sc_hs__and2_2 _50671_ (.A(_18423_),
    .B(_18424_),
    .Y(_18425_));
 sky130_as_sc_hs__or2_2 _50672_ (.A(net146),
    .B(_18425_),
    .Y(_18426_));
 sky130_as_sc_hs__and2_2 _50677_ (.A(_18428_),
    .B(_18429_),
    .Y(_18430_));
 sky130_as_sc_hs__or2_2 _50678_ (.A(net148),
    .B(_18430_),
    .Y(_18431_));
 sky130_as_sc_hs__and2_2 _50683_ (.A(_18433_),
    .B(_18434_),
    .Y(_18435_));
 sky130_as_sc_hs__or2_2 _50684_ (.A(net146),
    .B(_18435_),
    .Y(_18436_));
 sky130_as_sc_hs__and2_2 _50689_ (.A(_18438_),
    .B(_18439_),
    .Y(_18440_));
 sky130_as_sc_hs__or2_2 _50690_ (.A(net148),
    .B(_18440_),
    .Y(_18441_));
 sky130_as_sc_hs__and2_2 _50695_ (.A(_18443_),
    .B(_18444_),
    .Y(_18445_));
 sky130_as_sc_hs__or2_2 _50696_ (.A(net148),
    .B(_18445_),
    .Y(_18446_));
 sky130_as_sc_hs__and2_2 _50701_ (.A(_18448_),
    .B(_18449_),
    .Y(_18450_));
 sky130_as_sc_hs__or2_2 _50702_ (.A(net146),
    .B(_18450_),
    .Y(_18451_));
 sky130_as_sc_hs__and2_2 _50707_ (.A(_18453_),
    .B(_18454_),
    .Y(_18455_));
 sky130_as_sc_hs__or2_2 _50708_ (.A(net146),
    .B(_18455_),
    .Y(_18456_));
 sky130_as_sc_hs__and2_2 _50713_ (.A(_18458_),
    .B(_18459_),
    .Y(_18460_));
 sky130_as_sc_hs__or2_2 _50714_ (.A(net146),
    .B(_18460_),
    .Y(_18461_));
 sky130_as_sc_hs__and2_2 _50719_ (.A(_18463_),
    .B(_18464_),
    .Y(_18465_));
 sky130_as_sc_hs__or2_2 _50720_ (.A(net146),
    .B(_18465_),
    .Y(_18466_));
 sky130_as_sc_hs__and2_2 _50725_ (.A(_18468_),
    .B(_18469_),
    .Y(_18470_));
 sky130_as_sc_hs__or2_2 _50726_ (.A(net148),
    .B(_18470_),
    .Y(_18471_));
 sky130_as_sc_hs__and2_2 _50731_ (.A(_18473_),
    .B(_18474_),
    .Y(_18475_));
 sky130_as_sc_hs__or2_2 _50732_ (.A(net146),
    .B(_18475_),
    .Y(_18476_));
 sky130_as_sc_hs__and2_2 _50737_ (.A(_18478_),
    .B(_18479_),
    .Y(_18480_));
 sky130_as_sc_hs__or2_2 _50738_ (.A(net147),
    .B(_18480_),
    .Y(_18481_));
 sky130_as_sc_hs__and2_2 _50743_ (.A(_18483_),
    .B(_18484_),
    .Y(_18485_));
 sky130_as_sc_hs__or2_2 _50744_ (.A(net146),
    .B(_18485_),
    .Y(_18486_));
 sky130_as_sc_hs__and2_2 _50749_ (.A(_18488_),
    .B(_18489_),
    .Y(_18490_));
 sky130_as_sc_hs__or2_2 _50750_ (.A(net148),
    .B(_18490_),
    .Y(_18491_));
 sky130_as_sc_hs__and2_2 _50755_ (.A(_18493_),
    .B(_18494_),
    .Y(_18495_));
 sky130_as_sc_hs__or2_2 _50756_ (.A(net148),
    .B(_18495_),
    .Y(_18496_));
 sky130_as_sc_hs__and2_2 _50761_ (.A(_18498_),
    .B(_18499_),
    .Y(_18500_));
 sky130_as_sc_hs__or2_2 _50762_ (.A(net147),
    .B(_18500_),
    .Y(_18501_));
 sky130_as_sc_hs__and2_2 _50767_ (.A(_18503_),
    .B(_18504_),
    .Y(_18505_));
 sky130_as_sc_hs__or2_2 _50768_ (.A(net147),
    .B(_18505_),
    .Y(_18506_));
 sky130_as_sc_hs__and2_2 _50773_ (.A(_18508_),
    .B(_18509_),
    .Y(_18510_));
 sky130_as_sc_hs__or2_2 _50774_ (.A(net146),
    .B(_18510_),
    .Y(_18511_));
 sky130_as_sc_hs__and2_2 _50779_ (.A(_18513_),
    .B(_18514_),
    .Y(_18515_));
 sky130_as_sc_hs__or2_2 _50780_ (.A(net147),
    .B(_18515_),
    .Y(_18516_));
 sky130_as_sc_hs__and2_2 _50785_ (.A(_18518_),
    .B(_18519_),
    .Y(_18520_));
 sky130_as_sc_hs__or2_2 _50786_ (.A(net147),
    .B(_18520_),
    .Y(_18521_));
 sky130_as_sc_hs__and2_2 _50791_ (.A(_18523_),
    .B(_18524_),
    .Y(_18525_));
 sky130_as_sc_hs__or2_2 _50792_ (.A(net146),
    .B(_18525_),
    .Y(_18526_));
 sky130_as_sc_hs__and2_2 _50797_ (.A(_18528_),
    .B(_18529_),
    .Y(_18530_));
 sky130_as_sc_hs__or2_2 _50798_ (.A(net146),
    .B(_18530_),
    .Y(_18531_));
 sky130_as_sc_hs__and2_2 _50803_ (.A(_18533_),
    .B(_18534_),
    .Y(_18535_));
 sky130_as_sc_hs__or2_2 _50804_ (.A(net148),
    .B(_18535_),
    .Y(_18536_));
 sky130_as_sc_hs__and2_2 _50809_ (.A(_18538_),
    .B(_18539_),
    .Y(_18540_));
 sky130_as_sc_hs__or2_2 _50810_ (.A(net148),
    .B(_18540_),
    .Y(_18541_));
 sky130_as_sc_hs__and2_2 _50815_ (.A(_18543_),
    .B(_18544_),
    .Y(_18545_));
 sky130_as_sc_hs__or2_2 _50816_ (.A(net146),
    .B(_18545_),
    .Y(_18546_));
 sky130_as_sc_hs__and2_2 _50821_ (.A(_18548_),
    .B(_18549_),
    .Y(_18550_));
 sky130_as_sc_hs__or2_2 _50822_ (.A(net146),
    .B(_18550_),
    .Y(_18551_));
 sky130_as_sc_hs__and2_2 _50827_ (.A(_18553_),
    .B(_18554_),
    .Y(_18555_));
 sky130_as_sc_hs__or2_2 _50828_ (.A(net147),
    .B(_18555_),
    .Y(_18556_));
 sky130_as_sc_hs__and2_2 _50833_ (.A(_18558_),
    .B(_18559_),
    .Y(_18560_));
 sky130_as_sc_hs__or2_2 _50834_ (.A(net148),
    .B(_18560_),
    .Y(_18561_));
 sky130_as_sc_hs__and2_2 _50839_ (.A(_18563_),
    .B(_18564_),
    .Y(_18565_));
 sky130_as_sc_hs__or2_2 _50840_ (.A(net146),
    .B(_18565_),
    .Y(_18566_));
 sky130_as_sc_hs__and2_2 _50843_ (.A(net500),
    .B(net14),
    .Y(_01568_));
 sky130_as_sc_hs__and2_2 _50844_ (.A(_19529_),
    .B(\tholin_riscv.irqs[0] ),
    .Y(_18568_));
 sky130_as_sc_hs__nor2_2 _50845_ (.A(\tholin_riscv.irqs[2] ),
    .B(_18568_),
    .Y(_18569_));
 sky130_as_sc_hs__or2_2 _50846_ (.A(net602),
    .B(_19941_),
    .Y(_18570_));
 sky130_as_sc_hs__and2_2 _50848_ (.A(net500),
    .B(_18571_),
    .Y(_18572_));
 sky130_as_sc_hs__and2_2 _50849_ (.A(net603),
    .B(_18572_),
    .Y(_01569_));
 sky130_as_sc_hs__and2_2 _50853_ (.A(net526),
    .B(_18575_),
    .Y(_01570_));
 sky130_as_sc_hs__and2_2 _50854_ (.A(_19901_),
    .B(_20725_),
    .Y(_18576_));
 sky130_as_sc_hs__nor2b_2 _50855_ (.A(\tholin_riscv.last_io_state ),
    .Y(_18577_),
    .B(net14));
 sky130_as_sc_hs__or2_2 _50856_ (.A(net1795),
    .B(_18577_),
    .Y(_18578_));
 sky130_as_sc_hs__nand3_2 _50857_ (.A(net548),
    .B(net494),
    .C(_18578_),
    .Y(_18579_));
 sky130_as_sc_hs__nor2_2 _50858_ (.A(_18576_),
    .B(net549),
    .Y(_01571_));
 sky130_as_sc_hs__and2_2 _50859_ (.A(net1722),
    .B(net98),
    .Y(_18580_));
 sky130_as_sc_hs__nand3_2 _50860_ (.A(_19901_),
    .B(_19908_),
    .C(_19921_),
    .Y(_18581_));
 sky130_as_sc_hs__nand3_2 _50861_ (.A(net551),
    .B(net495),
    .C(_18581_),
    .Y(_18582_));
 sky130_as_sc_hs__nor2_2 _50862_ (.A(_18580_),
    .B(net552),
    .Y(_01572_));
 sky130_as_sc_hs__and2_2 _50863_ (.A(net1496),
    .B(net500),
    .Y(_18583_));
 sky130_as_sc_hs__and2_2 _50864_ (.A(net1718),
    .B(_18583_),
    .Y(_01573_));
 sky130_as_sc_hs__and2_2 _50865_ (.A(_19901_),
    .B(_19913_),
    .Y(_18584_));
 sky130_as_sc_hs__or2_2 _50867_ (.A(net551),
    .B(_18584_),
    .Y(_18586_));
 sky130_as_sc_hs__or2_2 _50868_ (.A(net1597),
    .B(_18585_),
    .Y(_18587_));
 sky130_as_sc_hs__and2_2 _50869_ (.A(net495),
    .B(_18586_),
    .Y(_18588_));
 sky130_as_sc_hs__and2_2 _50870_ (.A(_18587_),
    .B(_18588_),
    .Y(_01574_));
 sky130_as_sc_hs__or2_2 _50871_ (.A(net1496),
    .B(_18584_),
    .Y(_18589_));
 sky130_as_sc_hs__and2_2 _50873_ (.A(net500),
    .B(net1497),
    .Y(_18591_));
 sky130_as_sc_hs__and2_2 _50874_ (.A(_18590_),
    .B(net1498),
    .Y(_01575_));
 sky130_as_sc_hs__or2_2 _50875_ (.A(net548),
    .B(_18584_),
    .Y(_18592_));
 sky130_as_sc_hs__or2_2 _50876_ (.A(\tholin_riscv.instr[0] ),
    .B(_18585_),
    .Y(_18593_));
 sky130_as_sc_hs__and2_2 _50877_ (.A(net495),
    .B(_18592_),
    .Y(_18594_));
 sky130_as_sc_hs__and2_2 _50878_ (.A(_18593_),
    .B(_18594_),
    .Y(_01576_));
 sky130_as_sc_hs__and2_2 _50879_ (.A(_19901_),
    .B(_20736_),
    .Y(_18595_));
 sky130_as_sc_hs__or2_2 _50881_ (.A(net1655),
    .B(_18595_),
    .Y(_18597_));
 sky130_as_sc_hs__or2_2 _50882_ (.A(\tholin_riscv.instr[0] ),
    .B(_18596_),
    .Y(_18598_));
 sky130_as_sc_hs__and2_2 _50883_ (.A(net514),
    .B(net1656),
    .Y(_18599_));
 sky130_as_sc_hs__and2_2 _50884_ (.A(_18598_),
    .B(_18599_),
    .Y(_01577_));
 sky130_as_sc_hs__or2_2 _50885_ (.A(net1650),
    .B(_18595_),
    .Y(_18600_));
 sky130_as_sc_hs__or2_2 _50886_ (.A(net1597),
    .B(_18596_),
    .Y(_18601_));
 sky130_as_sc_hs__and2_2 _50887_ (.A(net514),
    .B(net1651),
    .Y(_18602_));
 sky130_as_sc_hs__and2_2 _50888_ (.A(_18601_),
    .B(_18602_),
    .Y(_01578_));
 sky130_as_sc_hs__or2_2 _50889_ (.A(net1652),
    .B(_18595_),
    .Y(_18603_));
 sky130_as_sc_hs__and2_2 _50891_ (.A(net514),
    .B(net1653),
    .Y(_18605_));
 sky130_as_sc_hs__and2_2 _50892_ (.A(_18604_),
    .B(_18605_),
    .Y(_01579_));
 sky130_as_sc_hs__or2_2 _50893_ (.A(net1657),
    .B(_18595_),
    .Y(_18606_));
 sky130_as_sc_hs__and2_2 _50895_ (.A(net524),
    .B(net1658),
    .Y(_18608_));
 sky130_as_sc_hs__and2_2 _50896_ (.A(_18607_),
    .B(_18608_),
    .Y(_01580_));
 sky130_as_sc_hs__or2_2 _50897_ (.A(net1659),
    .B(_18595_),
    .Y(_18609_));
 sky130_as_sc_hs__and2_2 _50899_ (.A(net524),
    .B(net1660),
    .Y(_18611_));
 sky130_as_sc_hs__and2_2 _50900_ (.A(_18610_),
    .B(_18611_),
    .Y(_01581_));
 sky130_as_sc_hs__or2_2 _50901_ (.A(net1671),
    .B(_18595_),
    .Y(_18612_));
 sky130_as_sc_hs__and2_2 _50903_ (.A(net524),
    .B(net1672),
    .Y(_18614_));
 sky130_as_sc_hs__and2_2 _50904_ (.A(_18613_),
    .B(_18614_),
    .Y(_01582_));
 sky130_as_sc_hs__and2_2 _50905_ (.A(_19901_),
    .B(_20723_),
    .Y(_18615_));
 sky130_as_sc_hs__or2_2 _50908_ (.A(\tholin_riscv.instr[0] ),
    .B(_18616_),
    .Y(_18618_));
 sky130_as_sc_hs__and2_2 _50909_ (.A(net523),
    .B(_18617_),
    .Y(_18619_));
 sky130_as_sc_hs__and2_2 _50910_ (.A(_18618_),
    .B(_18619_),
    .Y(_01583_));
 sky130_as_sc_hs__or2_2 _50912_ (.A(net1597),
    .B(_18616_),
    .Y(_18621_));
 sky130_as_sc_hs__and2_2 _50913_ (.A(net523),
    .B(_18620_),
    .Y(_18622_));
 sky130_as_sc_hs__and2_2 _50914_ (.A(_18621_),
    .B(_18622_),
    .Y(_01584_));
 sky130_as_sc_hs__and2_2 _50917_ (.A(net22),
    .B(_18623_),
    .Y(_18625_));
 sky130_as_sc_hs__and2_2 _50918_ (.A(_18624_),
    .B(_18625_),
    .Y(_01585_));
 sky130_as_sc_hs__and2_2 _50921_ (.A(net527),
    .B(_18626_),
    .Y(_18628_));
 sky130_as_sc_hs__and2_2 _50922_ (.A(_18627_),
    .B(_18628_),
    .Y(_01586_));
 sky130_as_sc_hs__and2_2 _50925_ (.A(net527),
    .B(_18629_),
    .Y(_18631_));
 sky130_as_sc_hs__and2_2 _50926_ (.A(_18630_),
    .B(_18631_),
    .Y(_01587_));
 sky130_as_sc_hs__and2_2 _50929_ (.A(net527),
    .B(_18632_),
    .Y(_18634_));
 sky130_as_sc_hs__and2_2 _50930_ (.A(_18633_),
    .B(_18634_),
    .Y(_01588_));
 sky130_as_sc_hs__and2_2 _50931_ (.A(_12816_),
    .B(_13146_),
    .Y(_18635_));
 sky130_as_sc_hs__or2_2 _50934_ (.A(net678),
    .B(_18635_),
    .Y(_18638_));
 sky130_as_sc_hs__and2_2 _50935_ (.A(_18637_),
    .B(net679),
    .Y(_01589_));
 sky130_as_sc_hs__and2_2 _51032_ (.A(net495),
    .B(_18703_),
    .Y(_18704_));
 sky130_as_sc_hs__or2_2 _51033_ (.A(_19496_),
    .B(net596),
    .Y(_18705_));
 sky130_as_sc_hs__and2_2 _51034_ (.A(_18704_),
    .B(_18705_),
    .Y(_18706_));
 sky130_as_sc_hs__nor2_2 _51035_ (.A(net596),
    .B(_18704_),
    .Y(_18707_));
 sky130_as_sc_hs__nor2_2 _51036_ (.A(_18706_),
    .B(net597),
    .Y(_01621_));
 sky130_as_sc_hs__and2_2 _51037_ (.A(_13146_),
    .B(_13478_),
    .Y(_18708_));
 sky130_as_sc_hs__and2_2 _51038_ (.A(_06178_),
    .B(_18708_),
    .Y(_18709_));
 sky130_as_sc_hs__nor2_2 _51039_ (.A(_19528_),
    .B(_18708_),
    .Y(_18710_));
 sky130_as_sc_hs__and2_2 _51040_ (.A(net723),
    .B(_18710_),
    .Y(_18711_));
 sky130_as_sc_hs__or2_2 _51041_ (.A(_18709_),
    .B(net724),
    .Y(_01622_));
 sky130_as_sc_hs__and2_2 _51135_ (.A(_19948_),
    .B(_13045_),
    .Y(_18774_));
 sky130_as_sc_hs__or2_2 _51137_ (.A(\tholin_riscv.Iimm[2] ),
    .B(_05519_),
    .Y(_18776_));
 sky130_as_sc_hs__or2_2 _51138_ (.A(\tholin_riscv.Bimm[2] ),
    .B(net127),
    .Y(_18777_));
 sky130_as_sc_hs__or2_2 _51140_ (.A(_19471_),
    .B(_18778_),
    .Y(_18779_));
 sky130_as_sc_hs__or2_2 _51143_ (.A(_13051_),
    .B(_18781_),
    .Y(_18782_));
 sky130_as_sc_hs__nand3_2 _51145_ (.A(_13046_),
    .B(_18782_),
    .C(_18783_),
    .Y(_18784_));
 sky130_as_sc_hs__or2_2 _51146_ (.A(_06873_),
    .B(_13065_),
    .Y(_18785_));
 sky130_as_sc_hs__and2_2 _51147_ (.A(_19990_),
    .B(_18785_),
    .Y(_18786_));
 sky130_as_sc_hs__nand3_2 _51148_ (.A(_18775_),
    .B(_18784_),
    .C(_18786_),
    .Y(_18787_));
 sky130_as_sc_hs__nand3_2 _51151_ (.A(net135),
    .B(_18788_),
    .C(_18789_),
    .Y(_18790_));
 sky130_as_sc_hs__nand3_2 _51152_ (.A(_19942_),
    .B(_18787_),
    .C(_18790_),
    .Y(_18791_));
 sky130_as_sc_hs__nand3_2 _51154_ (.A(_19944_),
    .B(_18791_),
    .C(_18792_),
    .Y(_18793_));
 sky130_as_sc_hs__and2_2 _51156_ (.A(net503),
    .B(_18794_),
    .Y(_18795_));
 sky130_as_sc_hs__and2_2 _51157_ (.A(_18793_),
    .B(_18795_),
    .Y(_01654_));
 sky130_as_sc_hs__or2_2 _51160_ (.A(\tholin_riscv.Bimm[3] ),
    .B(net127),
    .Y(_18798_));
 sky130_as_sc_hs__and2_2 _51161_ (.A(_18797_),
    .B(_18798_),
    .Y(_18799_));
 sky130_as_sc_hs__or2_2 _51163_ (.A(\tholin_riscv.PC[3] ),
    .B(_18799_),
    .Y(_18801_));
 sky130_as_sc_hs__or2_2 _51168_ (.A(_18802_),
    .B(_18803_),
    .Y(_18806_));
 sky130_as_sc_hs__nand3_2 _51169_ (.A(_13046_),
    .B(_18805_),
    .C(_18806_),
    .Y(_18807_));
 sky130_as_sc_hs__nand3_2 _51171_ (.A(_18796_),
    .B(_18807_),
    .C(_18808_),
    .Y(_18809_));
 sky130_as_sc_hs__nand3_2 _51175_ (.A(net135),
    .B(_18811_),
    .C(_18812_),
    .Y(_18813_));
 sky130_as_sc_hs__nand3_2 _51176_ (.A(_19942_),
    .B(_18810_),
    .C(_18813_),
    .Y(_18814_));
 sky130_as_sc_hs__nand3_2 _51178_ (.A(_19944_),
    .B(_18814_),
    .C(_18815_),
    .Y(_18816_));
 sky130_as_sc_hs__or2_2 _51179_ (.A(net1680),
    .B(_19944_),
    .Y(_18817_));
 sky130_as_sc_hs__and2_2 _51180_ (.A(net503),
    .B(_18817_),
    .Y(_18818_));
 sky130_as_sc_hs__and2_2 _51181_ (.A(_18816_),
    .B(_18818_),
    .Y(_01655_));
 sky130_as_sc_hs__or2_2 _51184_ (.A(\tholin_riscv.Bimm[4] ),
    .B(net127),
    .Y(_18821_));
 sky130_as_sc_hs__and2_2 _51185_ (.A(_18820_),
    .B(_18821_),
    .Y(_18822_));
 sky130_as_sc_hs__or2_2 _51187_ (.A(\tholin_riscv.PC[4] ),
    .B(_18822_),
    .Y(_18824_));
 sky130_as_sc_hs__and2_2 _51188_ (.A(_18823_),
    .B(_18824_),
    .Y(_18825_));
 sky130_as_sc_hs__or2_2 _51191_ (.A(_18825_),
    .B(_18826_),
    .Y(_18828_));
 sky130_as_sc_hs__nand3_2 _51195_ (.A(_18819_),
    .B(_18830_),
    .C(_18831_),
    .Y(_18832_));
 sky130_as_sc_hs__nand3_2 _51199_ (.A(net135),
    .B(_18834_),
    .C(_18835_),
    .Y(_18836_));
 sky130_as_sc_hs__nand3_2 _51200_ (.A(_19942_),
    .B(_18833_),
    .C(_18836_),
    .Y(_18837_));
 sky130_as_sc_hs__nand3_2 _51202_ (.A(_19944_),
    .B(_18837_),
    .C(_18838_),
    .Y(_18839_));
 sky130_as_sc_hs__or2_2 _51203_ (.A(net1667),
    .B(_19944_),
    .Y(_18840_));
 sky130_as_sc_hs__and2_2 _51204_ (.A(net503),
    .B(net1668),
    .Y(_18841_));
 sky130_as_sc_hs__and2_2 _51205_ (.A(_18839_),
    .B(_18841_),
    .Y(_01656_));
 sky130_as_sc_hs__or2_2 _51206_ (.A(\tholin_riscv.PCE[5] ),
    .B(_13062_),
    .Y(_18842_));
 sky130_as_sc_hs__or2_2 _51207_ (.A(_07848_),
    .B(_13061_),
    .Y(_18843_));
 sky130_as_sc_hs__nand3_2 _51208_ (.A(net136),
    .B(_18842_),
    .C(_18843_),
    .Y(_18844_));
 sky130_as_sc_hs__or2_2 _51209_ (.A(\tholin_riscv.PC[5] ),
    .B(\tholin_riscv.Bimm[5] ),
    .Y(_18845_));
 sky130_as_sc_hs__and2_2 _51211_ (.A(_18845_),
    .B(_18846_),
    .Y(_18847_));
 sky130_as_sc_hs__or2_2 _51213_ (.A(_18847_),
    .B(_18848_),
    .Y(_18849_));
 sky130_as_sc_hs__nand3_2 _51215_ (.A(_13046_),
    .B(_18849_),
    .C(_18850_),
    .Y(_18851_));
 sky130_as_sc_hs__or2_2 _51217_ (.A(_07795_),
    .B(_13065_),
    .Y(_18853_));
 sky130_as_sc_hs__nand3_2 _51218_ (.A(_18851_),
    .B(_18852_),
    .C(_18853_),
    .Y(_18854_));
 sky130_as_sc_hs__nand3_2 _51223_ (.A(_19944_),
    .B(_18857_),
    .C(_18858_),
    .Y(_18859_));
 sky130_as_sc_hs__or2_2 _51224_ (.A(net1661),
    .B(_19944_),
    .Y(_18860_));
 sky130_as_sc_hs__and2_2 _51225_ (.A(net503),
    .B(net1662),
    .Y(_18861_));
 sky130_as_sc_hs__and2_2 _51226_ (.A(_18859_),
    .B(_18861_),
    .Y(_01657_));
 sky130_as_sc_hs__or2_2 _51228_ (.A(\tholin_riscv.PC[6] ),
    .B(\tholin_riscv.Bimm[6] ),
    .Y(_18863_));
 sky130_as_sc_hs__or2_2 _51234_ (.A(_18865_),
    .B(_18867_),
    .Y(_18869_));
 sky130_as_sc_hs__nand3_2 _51235_ (.A(_13046_),
    .B(_18868_),
    .C(_18869_),
    .Y(_18870_));
 sky130_as_sc_hs__nand3_2 _51237_ (.A(_18862_),
    .B(_18870_),
    .C(_18871_),
    .Y(_18872_));
 sky130_as_sc_hs__nand3_2 _51241_ (.A(net136),
    .B(_18874_),
    .C(_18875_),
    .Y(_18876_));
 sky130_as_sc_hs__nand3_2 _51242_ (.A(_19942_),
    .B(_18873_),
    .C(_18876_),
    .Y(_18877_));
 sky130_as_sc_hs__nand3_2 _51244_ (.A(_19944_),
    .B(_18877_),
    .C(_18878_),
    .Y(_18879_));
 sky130_as_sc_hs__or2_2 _51245_ (.A(net1673),
    .B(_19944_),
    .Y(_18880_));
 sky130_as_sc_hs__and2_2 _51246_ (.A(net503),
    .B(_18880_),
    .Y(_18881_));
 sky130_as_sc_hs__and2_2 _51247_ (.A(_18879_),
    .B(_18881_),
    .Y(_01658_));
 sky130_as_sc_hs__or2_2 _51249_ (.A(\tholin_riscv.PC[7] ),
    .B(\tholin_riscv.Bimm[7] ),
    .Y(_18883_));
 sky130_as_sc_hs__or2_2 _51255_ (.A(_18885_),
    .B(_18887_),
    .Y(_18889_));
 sky130_as_sc_hs__nand3_2 _51256_ (.A(_13046_),
    .B(_18888_),
    .C(_18889_),
    .Y(_18890_));
 sky130_as_sc_hs__nand3_2 _51258_ (.A(_18882_),
    .B(_18890_),
    .C(_18891_),
    .Y(_18892_));
 sky130_as_sc_hs__nand3_2 _51262_ (.A(net135),
    .B(_18894_),
    .C(_18895_),
    .Y(_18896_));
 sky130_as_sc_hs__nand3_2 _51263_ (.A(_19942_),
    .B(_18893_),
    .C(_18896_),
    .Y(_18897_));
 sky130_as_sc_hs__nand3_2 _51265_ (.A(_19944_),
    .B(_18897_),
    .C(_18898_),
    .Y(_18899_));
 sky130_as_sc_hs__or2_2 _51266_ (.A(net1687),
    .B(_19944_),
    .Y(_18900_));
 sky130_as_sc_hs__and2_2 _51267_ (.A(net503),
    .B(_18900_),
    .Y(_18901_));
 sky130_as_sc_hs__and2_2 _51268_ (.A(_18899_),
    .B(_18901_),
    .Y(_01659_));
 sky130_as_sc_hs__or2_2 _51270_ (.A(\tholin_riscv.PC[8] ),
    .B(\tholin_riscv.Bimm[8] ),
    .Y(_18903_));
 sky130_as_sc_hs__or2_2 _51276_ (.A(_18905_),
    .B(_18907_),
    .Y(_18909_));
 sky130_as_sc_hs__nand3_2 _51277_ (.A(_13046_),
    .B(_18908_),
    .C(_18909_),
    .Y(_18910_));
 sky130_as_sc_hs__nand3_2 _51279_ (.A(_18902_),
    .B(_18910_),
    .C(_18911_),
    .Y(_18912_));
 sky130_as_sc_hs__nand3_2 _51283_ (.A(net135),
    .B(_18914_),
    .C(_18915_),
    .Y(_18916_));
 sky130_as_sc_hs__nand3_2 _51284_ (.A(_19942_),
    .B(_18913_),
    .C(_18916_),
    .Y(_18917_));
 sky130_as_sc_hs__nand3_2 _51286_ (.A(_19944_),
    .B(_18917_),
    .C(_18918_),
    .Y(_18919_));
 sky130_as_sc_hs__or2_2 _51287_ (.A(net1669),
    .B(_19944_),
    .Y(_18920_));
 sky130_as_sc_hs__and2_2 _51288_ (.A(net502),
    .B(net1670),
    .Y(_18921_));
 sky130_as_sc_hs__and2_2 _51289_ (.A(_18919_),
    .B(_18921_),
    .Y(_01660_));
 sky130_as_sc_hs__or2_2 _51290_ (.A(_08943_),
    .B(_13061_),
    .Y(_18922_));
 sky130_as_sc_hs__or2_2 _51291_ (.A(\tholin_riscv.PCE[9] ),
    .B(_13062_),
    .Y(_18923_));
 sky130_as_sc_hs__nand3_2 _51292_ (.A(net136),
    .B(_18922_),
    .C(_18923_),
    .Y(_18924_));
 sky130_as_sc_hs__or2_2 _51294_ (.A(\tholin_riscv.PC[9] ),
    .B(\tholin_riscv.Bimm[9] ),
    .Y(_18926_));
 sky130_as_sc_hs__and2_2 _51295_ (.A(_18925_),
    .B(_18926_),
    .Y(_18927_));
 sky130_as_sc_hs__or2_2 _51298_ (.A(_18927_),
    .B(_18929_),
    .Y(_18930_));
 sky130_as_sc_hs__nand3_2 _51300_ (.A(_13046_),
    .B(_18930_),
    .C(_18931_),
    .Y(_18932_));
 sky130_as_sc_hs__or2_2 _51302_ (.A(_08902_),
    .B(_13065_),
    .Y(_18934_));
 sky130_as_sc_hs__nand3_2 _51303_ (.A(_18932_),
    .B(_18933_),
    .C(_18934_),
    .Y(_18935_));
 sky130_as_sc_hs__nand3_2 _51308_ (.A(_19944_),
    .B(_18938_),
    .C(_18939_),
    .Y(_18940_));
 sky130_as_sc_hs__or2_2 _51309_ (.A(net1676),
    .B(_19944_),
    .Y(_18941_));
 sky130_as_sc_hs__and2_2 _51310_ (.A(net502),
    .B(net1677),
    .Y(_18942_));
 sky130_as_sc_hs__and2_2 _51311_ (.A(_18940_),
    .B(_18942_),
    .Y(_01661_));
 sky130_as_sc_hs__or2_2 _51313_ (.A(\tholin_riscv.PC[10] ),
    .B(\tholin_riscv.Bimm[10] ),
    .Y(_18944_));
 sky130_as_sc_hs__or2_2 _51319_ (.A(_18946_),
    .B(_18948_),
    .Y(_18950_));
 sky130_as_sc_hs__nand3_2 _51320_ (.A(_13046_),
    .B(_18949_),
    .C(_18950_),
    .Y(_18951_));
 sky130_as_sc_hs__nand3_2 _51322_ (.A(_18943_),
    .B(_18951_),
    .C(_18952_),
    .Y(_18953_));
 sky130_as_sc_hs__nand3_2 _51326_ (.A(net135),
    .B(_18955_),
    .C(_18956_),
    .Y(_18957_));
 sky130_as_sc_hs__nand3_2 _51327_ (.A(_19942_),
    .B(_18954_),
    .C(_18957_),
    .Y(_18958_));
 sky130_as_sc_hs__nand3_2 _51329_ (.A(_19944_),
    .B(_18958_),
    .C(_18959_),
    .Y(_18960_));
 sky130_as_sc_hs__or2_2 _51330_ (.A(net1663),
    .B(_19944_),
    .Y(_18961_));
 sky130_as_sc_hs__and2_2 _51331_ (.A(net502),
    .B(net1664),
    .Y(_18962_));
 sky130_as_sc_hs__and2_2 _51332_ (.A(_18960_),
    .B(_18962_),
    .Y(_01662_));
 sky130_as_sc_hs__or2_2 _51334_ (.A(\tholin_riscv.Iimm[0] ),
    .B(_05519_),
    .Y(_18964_));
 sky130_as_sc_hs__or2_2 _51335_ (.A(\tholin_riscv.Bimm[11] ),
    .B(net127),
    .Y(_18965_));
 sky130_as_sc_hs__and2_2 _51336_ (.A(_18964_),
    .B(_18965_),
    .Y(_18966_));
 sky130_as_sc_hs__or2_2 _51338_ (.A(\tholin_riscv.PC[11] ),
    .B(_18966_),
    .Y(_18968_));
 sky130_as_sc_hs__or2_2 _51342_ (.A(_18969_),
    .B(_18971_),
    .Y(_18972_));
 sky130_as_sc_hs__nand3_2 _51344_ (.A(_13046_),
    .B(_18972_),
    .C(_18973_),
    .Y(_18974_));
 sky130_as_sc_hs__nand3_2 _51346_ (.A(_18963_),
    .B(_18974_),
    .C(_18975_),
    .Y(_18976_));
 sky130_as_sc_hs__nand3_2 _51350_ (.A(net135),
    .B(_18978_),
    .C(_18979_),
    .Y(_18980_));
 sky130_as_sc_hs__nand3_2 _51351_ (.A(_19942_),
    .B(_18977_),
    .C(_18980_),
    .Y(_18981_));
 sky130_as_sc_hs__nand3_2 _51353_ (.A(_19944_),
    .B(_18981_),
    .C(_18982_),
    .Y(_18983_));
 sky130_as_sc_hs__or2_2 _51354_ (.A(net1674),
    .B(_19944_),
    .Y(_18984_));
 sky130_as_sc_hs__and2_2 _51355_ (.A(net502),
    .B(net1675),
    .Y(_18985_));
 sky130_as_sc_hs__and2_2 _51356_ (.A(_18983_),
    .B(_18985_),
    .Y(_01663_));
 sky130_as_sc_hs__or2_2 _51358_ (.A(net334),
    .B(net127),
    .Y(_18987_));
 sky130_as_sc_hs__and2_2 _51360_ (.A(_18987_),
    .B(_18988_),
    .Y(_18989_));
 sky130_as_sc_hs__or2_2 _51362_ (.A(\tholin_riscv.PC[12] ),
    .B(_18989_),
    .Y(_18991_));
 sky130_as_sc_hs__and2_2 _51363_ (.A(_18990_),
    .B(_18991_),
    .Y(_18992_));
 sky130_as_sc_hs__or2_2 _51367_ (.A(_18992_),
    .B(_18994_),
    .Y(_18996_));
 sky130_as_sc_hs__nand3_2 _51371_ (.A(_18986_),
    .B(_18998_),
    .C(_18999_),
    .Y(_19000_));
 sky130_as_sc_hs__or2_2 _51373_ (.A(_09674_),
    .B(net125),
    .Y(_19002_));
 sky130_as_sc_hs__nand3_2 _51375_ (.A(net135),
    .B(_19002_),
    .C(_19003_),
    .Y(_19004_));
 sky130_as_sc_hs__nand3_2 _51376_ (.A(_19942_),
    .B(_19001_),
    .C(_19004_),
    .Y(_19005_));
 sky130_as_sc_hs__nand3_2 _51378_ (.A(_19944_),
    .B(_19005_),
    .C(_19006_),
    .Y(_19007_));
 sky130_as_sc_hs__or2_2 _51379_ (.A(net1706),
    .B(_19944_),
    .Y(_19008_));
 sky130_as_sc_hs__and2_2 _51380_ (.A(net497),
    .B(_19008_),
    .Y(_19009_));
 sky130_as_sc_hs__and2_2 _51381_ (.A(_19007_),
    .B(_19009_),
    .Y(_01664_));
 sky130_as_sc_hs__and2_2 _51384_ (.A(_18987_),
    .B(_19011_),
    .Y(_19012_));
 sky130_as_sc_hs__or2_2 _51386_ (.A(\tholin_riscv.PC[13] ),
    .B(_19012_),
    .Y(_19014_));
 sky130_as_sc_hs__or2_2 _51390_ (.A(_19015_),
    .B(_19016_),
    .Y(_19018_));
 sky130_as_sc_hs__nand3_2 _51391_ (.A(_13046_),
    .B(_19017_),
    .C(_19018_),
    .Y(_19019_));
 sky130_as_sc_hs__nand3_2 _51393_ (.A(_19010_),
    .B(_19019_),
    .C(_19020_),
    .Y(_19021_));
 sky130_as_sc_hs__or2_2 _51395_ (.A(_09896_),
    .B(net125),
    .Y(_19023_));
 sky130_as_sc_hs__nand3_2 _51397_ (.A(net135),
    .B(_19023_),
    .C(_19024_),
    .Y(_19025_));
 sky130_as_sc_hs__nand3_2 _51398_ (.A(_19942_),
    .B(_19022_),
    .C(_19025_),
    .Y(_19026_));
 sky130_as_sc_hs__nand3_2 _51400_ (.A(_19944_),
    .B(_19026_),
    .C(_19027_),
    .Y(_19028_));
 sky130_as_sc_hs__or2_2 _51401_ (.A(net1679),
    .B(_19944_),
    .Y(_19029_));
 sky130_as_sc_hs__and2_2 _51402_ (.A(net497),
    .B(_19029_),
    .Y(_19030_));
 sky130_as_sc_hs__and2_2 _51403_ (.A(_19028_),
    .B(_19030_),
    .Y(_01665_));
 sky130_as_sc_hs__or2_2 _51405_ (.A(net411),
    .B(_05519_),
    .Y(_19032_));
 sky130_as_sc_hs__and2_2 _51406_ (.A(_18987_),
    .B(_19032_),
    .Y(_19033_));
 sky130_as_sc_hs__or2_2 _51408_ (.A(\tholin_riscv.PC[14] ),
    .B(_19033_),
    .Y(_19035_));
 sky130_as_sc_hs__and2_2 _51409_ (.A(_19034_),
    .B(_19035_),
    .Y(_19036_));
 sky130_as_sc_hs__or2_2 _51413_ (.A(_19036_),
    .B(_19038_),
    .Y(_19040_));
 sky130_as_sc_hs__nand3_2 _51417_ (.A(_19031_),
    .B(_19042_),
    .C(_19043_),
    .Y(_19044_));
 sky130_as_sc_hs__or2_2 _51419_ (.A(_10122_),
    .B(net125),
    .Y(_19046_));
 sky130_as_sc_hs__nand3_2 _51421_ (.A(net135),
    .B(_19046_),
    .C(_19047_),
    .Y(_19048_));
 sky130_as_sc_hs__nand3_2 _51422_ (.A(_19942_),
    .B(_19045_),
    .C(_19048_),
    .Y(_19049_));
 sky130_as_sc_hs__nand3_2 _51424_ (.A(_19944_),
    .B(_19049_),
    .C(_19050_),
    .Y(_19051_));
 sky130_as_sc_hs__or2_2 _51425_ (.A(net1681),
    .B(_19944_),
    .Y(_19052_));
 sky130_as_sc_hs__and2_2 _51426_ (.A(net499),
    .B(_19052_),
    .Y(_19053_));
 sky130_as_sc_hs__and2_2 _51427_ (.A(_19051_),
    .B(_19053_),
    .Y(_01666_));
 sky130_as_sc_hs__and2_2 _51430_ (.A(_18987_),
    .B(_19055_),
    .Y(_19056_));
 sky130_as_sc_hs__or2_2 _51432_ (.A(\tholin_riscv.PC[15] ),
    .B(_19056_),
    .Y(_19058_));
 sky130_as_sc_hs__or2_2 _51436_ (.A(_19059_),
    .B(_19060_),
    .Y(_19062_));
 sky130_as_sc_hs__nand3_2 _51437_ (.A(_13046_),
    .B(_19061_),
    .C(_19062_),
    .Y(_19063_));
 sky130_as_sc_hs__nand3_2 _51439_ (.A(_19054_),
    .B(_19063_),
    .C(_19064_),
    .Y(_19065_));
 sky130_as_sc_hs__or2_2 _51441_ (.A(_10334_),
    .B(net125),
    .Y(_19067_));
 sky130_as_sc_hs__nand3_2 _51443_ (.A(net135),
    .B(_19067_),
    .C(_19068_),
    .Y(_19069_));
 sky130_as_sc_hs__nand3_2 _51444_ (.A(_19942_),
    .B(_19066_),
    .C(_19069_),
    .Y(_19070_));
 sky130_as_sc_hs__nand3_2 _51446_ (.A(_19944_),
    .B(_19070_),
    .C(_19071_),
    .Y(_19072_));
 sky130_as_sc_hs__or2_2 _51447_ (.A(net1692),
    .B(_19944_),
    .Y(_19073_));
 sky130_as_sc_hs__and2_2 _51448_ (.A(net498),
    .B(_19073_),
    .Y(_19074_));
 sky130_as_sc_hs__and2_2 _51449_ (.A(_19072_),
    .B(_19074_),
    .Y(_01667_));
 sky130_as_sc_hs__and2_2 _51452_ (.A(_18987_),
    .B(_19076_),
    .Y(_19077_));
 sky130_as_sc_hs__or2_2 _51454_ (.A(\tholin_riscv.PC[16] ),
    .B(_19077_),
    .Y(_19079_));
 sky130_as_sc_hs__and2_2 _51455_ (.A(_19078_),
    .B(_19079_),
    .Y(_19080_));
 sky130_as_sc_hs__or2_2 _51459_ (.A(_19080_),
    .B(_19082_),
    .Y(_19084_));
 sky130_as_sc_hs__nand3_2 _51463_ (.A(_19075_),
    .B(_19086_),
    .C(_19087_),
    .Y(_19088_));
 sky130_as_sc_hs__or2_2 _51465_ (.A(_10549_),
    .B(net125),
    .Y(_19090_));
 sky130_as_sc_hs__nand3_2 _51467_ (.A(net135),
    .B(_19090_),
    .C(_19091_),
    .Y(_19092_));
 sky130_as_sc_hs__nand3_2 _51468_ (.A(_19942_),
    .B(_19089_),
    .C(_19092_),
    .Y(_19093_));
 sky130_as_sc_hs__nand3_2 _51470_ (.A(_19944_),
    .B(_19093_),
    .C(_19094_),
    .Y(_19095_));
 sky130_as_sc_hs__or2_2 _51471_ (.A(net1701),
    .B(_19944_),
    .Y(_19096_));
 sky130_as_sc_hs__and2_2 _51472_ (.A(net499),
    .B(_19096_),
    .Y(_19097_));
 sky130_as_sc_hs__and2_2 _51473_ (.A(_19095_),
    .B(_19097_),
    .Y(_01668_));
 sky130_as_sc_hs__and2_2 _51476_ (.A(_18987_),
    .B(_19099_),
    .Y(_19100_));
 sky130_as_sc_hs__or2_2 _51478_ (.A(\tholin_riscv.PC[17] ),
    .B(_19100_),
    .Y(_19102_));
 sky130_as_sc_hs__or2_2 _51482_ (.A(_19103_),
    .B(_19104_),
    .Y(_19106_));
 sky130_as_sc_hs__nand3_2 _51483_ (.A(_13046_),
    .B(_19105_),
    .C(_19106_),
    .Y(_19107_));
 sky130_as_sc_hs__nand3_2 _51485_ (.A(_19098_),
    .B(_19107_),
    .C(_19108_),
    .Y(_19109_));
 sky130_as_sc_hs__or2_2 _51487_ (.A(_10740_),
    .B(net125),
    .Y(_19111_));
 sky130_as_sc_hs__nand3_2 _51489_ (.A(net135),
    .B(_19111_),
    .C(_19112_),
    .Y(_19113_));
 sky130_as_sc_hs__nand3_2 _51490_ (.A(_19942_),
    .B(_19110_),
    .C(_19113_),
    .Y(_19114_));
 sky130_as_sc_hs__nand3_2 _51492_ (.A(_19944_),
    .B(_19114_),
    .C(_19115_),
    .Y(_19116_));
 sky130_as_sc_hs__or2_2 _51493_ (.A(net1700),
    .B(_19944_),
    .Y(_19117_));
 sky130_as_sc_hs__and2_2 _51494_ (.A(net499),
    .B(_19117_),
    .Y(_19118_));
 sky130_as_sc_hs__and2_2 _51495_ (.A(_19116_),
    .B(_19118_),
    .Y(_01669_));
 sky130_as_sc_hs__and2_2 _51498_ (.A(_18987_),
    .B(_19120_),
    .Y(_19121_));
 sky130_as_sc_hs__or2_2 _51499_ (.A(\tholin_riscv.PC[18] ),
    .B(_19121_),
    .Y(_19122_));
 sky130_as_sc_hs__and2_2 _51501_ (.A(_19122_),
    .B(_19123_),
    .Y(_19124_));
 sky130_as_sc_hs__and2_2 _51503_ (.A(_19101_),
    .B(_19125_),
    .Y(_19126_));
 sky130_as_sc_hs__or2_2 _51504_ (.A(_19124_),
    .B(_19126_),
    .Y(_19127_));
 sky130_as_sc_hs__nand3_2 _51506_ (.A(_13046_),
    .B(_19127_),
    .C(_19128_),
    .Y(_19129_));
 sky130_as_sc_hs__nand3_2 _51508_ (.A(_19119_),
    .B(_19129_),
    .C(_19130_),
    .Y(_19131_));
 sky130_as_sc_hs__or2_2 _51510_ (.A(_10930_),
    .B(net125),
    .Y(_19133_));
 sky130_as_sc_hs__nand3_2 _51512_ (.A(net135),
    .B(_19133_),
    .C(_19134_),
    .Y(_19135_));
 sky130_as_sc_hs__nand3_2 _51513_ (.A(_19942_),
    .B(_19132_),
    .C(_19135_),
    .Y(_19136_));
 sky130_as_sc_hs__nand3_2 _51515_ (.A(_19944_),
    .B(_19136_),
    .C(_19137_),
    .Y(_19138_));
 sky130_as_sc_hs__or2_2 _51516_ (.A(net1698),
    .B(_19944_),
    .Y(_19139_));
 sky130_as_sc_hs__and2_2 _51517_ (.A(net499),
    .B(_19139_),
    .Y(_19140_));
 sky130_as_sc_hs__and2_2 _51518_ (.A(_19138_),
    .B(_19140_),
    .Y(_01670_));
 sky130_as_sc_hs__and2_2 _51521_ (.A(_18987_),
    .B(_19142_),
    .Y(_19143_));
 sky130_as_sc_hs__or2_2 _51522_ (.A(\tholin_riscv.PC[19] ),
    .B(_19143_),
    .Y(_19144_));
 sky130_as_sc_hs__and2_2 _51524_ (.A(_19144_),
    .B(_19145_),
    .Y(_19146_));
 sky130_as_sc_hs__or2_2 _51527_ (.A(_19146_),
    .B(_19148_),
    .Y(_19149_));
 sky130_as_sc_hs__nand3_2 _51529_ (.A(_13046_),
    .B(_19149_),
    .C(_19150_),
    .Y(_19151_));
 sky130_as_sc_hs__nand3_2 _51531_ (.A(_19141_),
    .B(_19151_),
    .C(_19152_),
    .Y(_19153_));
 sky130_as_sc_hs__nand3_2 _51535_ (.A(net135),
    .B(_19155_),
    .C(_19156_),
    .Y(_19157_));
 sky130_as_sc_hs__nand3_2 _51536_ (.A(_19942_),
    .B(_19154_),
    .C(_19157_),
    .Y(_19158_));
 sky130_as_sc_hs__nand3_2 _51538_ (.A(_19944_),
    .B(_19158_),
    .C(_19159_),
    .Y(_19160_));
 sky130_as_sc_hs__or2_2 _51539_ (.A(net1708),
    .B(_19944_),
    .Y(_19161_));
 sky130_as_sc_hs__and2_2 _51540_ (.A(net504),
    .B(_19161_),
    .Y(_19162_));
 sky130_as_sc_hs__and2_2 _51541_ (.A(_19160_),
    .B(_19162_),
    .Y(_01671_));
 sky130_as_sc_hs__or2_2 _51543_ (.A(\tholin_riscv.PC[20] ),
    .B(net334),
    .Y(_19164_));
 sky130_as_sc_hs__and2_2 _51545_ (.A(_19164_),
    .B(_19165_),
    .Y(_19166_));
 sky130_as_sc_hs__or2_2 _51548_ (.A(_19166_),
    .B(_19168_),
    .Y(_19169_));
 sky130_as_sc_hs__nand3_2 _51550_ (.A(_13046_),
    .B(_19169_),
    .C(_19170_),
    .Y(_19171_));
 sky130_as_sc_hs__nand3_2 _51552_ (.A(_19163_),
    .B(_19171_),
    .C(_19172_),
    .Y(_19173_));
 sky130_as_sc_hs__or2_2 _51554_ (.A(_11288_),
    .B(net125),
    .Y(_19175_));
 sky130_as_sc_hs__nand3_2 _51556_ (.A(net136),
    .B(_19175_),
    .C(_19176_),
    .Y(_19177_));
 sky130_as_sc_hs__nand3_2 _51557_ (.A(_19942_),
    .B(_19174_),
    .C(_19177_),
    .Y(_19178_));
 sky130_as_sc_hs__nand3_2 _51559_ (.A(_19944_),
    .B(_19178_),
    .C(_19179_),
    .Y(_19180_));
 sky130_as_sc_hs__or2_2 _51560_ (.A(net1702),
    .B(_19944_),
    .Y(_19181_));
 sky130_as_sc_hs__and2_2 _51561_ (.A(net504),
    .B(_19181_),
    .Y(_19182_));
 sky130_as_sc_hs__and2_2 _51562_ (.A(_19180_),
    .B(_19182_),
    .Y(_01672_));
 sky130_as_sc_hs__or2_2 _51564_ (.A(\tholin_riscv.PC[21] ),
    .B(net334),
    .Y(_19184_));
 sky130_as_sc_hs__and2_2 _51566_ (.A(_19184_),
    .B(_19185_),
    .Y(_19186_));
 sky130_as_sc_hs__and2_2 _51568_ (.A(_19164_),
    .B(_19187_),
    .Y(_19188_));
 sky130_as_sc_hs__nor2_2 _51569_ (.A(_19186_),
    .B(_19188_),
    .Y(_19189_));
 sky130_as_sc_hs__and2_2 _51570_ (.A(_19186_),
    .B(_19188_),
    .Y(_19190_));
 sky130_as_sc_hs__or2_2 _51571_ (.A(_19189_),
    .B(_19190_),
    .Y(_19191_));
 sky130_as_sc_hs__nand3_2 _51574_ (.A(_19183_),
    .B(_19192_),
    .C(_19193_),
    .Y(_19194_));
 sky130_as_sc_hs__or2_2 _51576_ (.A(_11457_),
    .B(net125),
    .Y(_19196_));
 sky130_as_sc_hs__nand3_2 _51578_ (.A(_19989_),
    .B(_19196_),
    .C(_19197_),
    .Y(_19198_));
 sky130_as_sc_hs__nand3_2 _51579_ (.A(_19942_),
    .B(_19195_),
    .C(_19198_),
    .Y(_19199_));
 sky130_as_sc_hs__nand3_2 _51581_ (.A(_19944_),
    .B(_19199_),
    .C(_19200_),
    .Y(_19201_));
 sky130_as_sc_hs__or2_2 _51582_ (.A(net1707),
    .B(_19944_),
    .Y(_19202_));
 sky130_as_sc_hs__and2_2 _51583_ (.A(net504),
    .B(_19202_),
    .Y(_19203_));
 sky130_as_sc_hs__and2_2 _51584_ (.A(_19201_),
    .B(_19203_),
    .Y(_01673_));
 sky130_as_sc_hs__or2_2 _51586_ (.A(\tholin_riscv.PC[22] ),
    .B(net334),
    .Y(_19205_));
 sky130_as_sc_hs__and2_2 _51588_ (.A(_19205_),
    .B(_19206_),
    .Y(_19207_));
 sky130_as_sc_hs__and2_2 _51590_ (.A(_19185_),
    .B(_19208_),
    .Y(_19209_));
 sky130_as_sc_hs__or2_2 _51591_ (.A(_19207_),
    .B(_19209_),
    .Y(_19210_));
 sky130_as_sc_hs__nand3_2 _51593_ (.A(_13046_),
    .B(_19210_),
    .C(_19211_),
    .Y(_19212_));
 sky130_as_sc_hs__nand3_2 _51595_ (.A(_19204_),
    .B(_19212_),
    .C(_19213_),
    .Y(_19214_));
 sky130_as_sc_hs__or2_2 _51597_ (.A(_11616_),
    .B(net125),
    .Y(_19216_));
 sky130_as_sc_hs__nand3_2 _51599_ (.A(net136),
    .B(_19216_),
    .C(_19217_),
    .Y(_19218_));
 sky130_as_sc_hs__nand3_2 _51600_ (.A(_19942_),
    .B(_19215_),
    .C(_19218_),
    .Y(_19219_));
 sky130_as_sc_hs__nand3_2 _51602_ (.A(_19944_),
    .B(_19219_),
    .C(_19220_),
    .Y(_19221_));
 sky130_as_sc_hs__or2_2 _51603_ (.A(net1704),
    .B(_19944_),
    .Y(_19222_));
 sky130_as_sc_hs__and2_2 _51604_ (.A(net504),
    .B(_19222_),
    .Y(_19223_));
 sky130_as_sc_hs__and2_2 _51605_ (.A(_19221_),
    .B(_19223_),
    .Y(_01674_));
 sky130_as_sc_hs__or2_2 _51607_ (.A(\tholin_riscv.PC[23] ),
    .B(net334),
    .Y(_19225_));
 sky130_as_sc_hs__inv_2 _51610_ (.Y(_19228_),
    .A(_19227_));
 sky130_as_sc_hs__and2_2 _51611_ (.A(_19185_),
    .B(_19206_),
    .Y(_19229_));
 sky130_as_sc_hs__and2_2 _51612_ (.A(_19190_),
    .B(_19207_),
    .Y(_19230_));
 sky130_as_sc_hs__nand2b_2 _51613_ (.B(_19229_),
    .Y(_19231_),
    .A(_19230_));
 sky130_as_sc_hs__or2_2 _51615_ (.A(_19227_),
    .B(_19231_),
    .Y(_19233_));
 sky130_as_sc_hs__nand3_2 _51616_ (.A(_13046_),
    .B(_19232_),
    .C(_19233_),
    .Y(_19234_));
 sky130_as_sc_hs__nand3_2 _51618_ (.A(_19224_),
    .B(_19234_),
    .C(_19235_),
    .Y(_19236_));
 sky130_as_sc_hs__nand3_2 _51622_ (.A(net136),
    .B(_19238_),
    .C(_19239_),
    .Y(_19240_));
 sky130_as_sc_hs__nand3_2 _51623_ (.A(_19942_),
    .B(_19237_),
    .C(_19240_),
    .Y(_19241_));
 sky130_as_sc_hs__nand3_2 _51625_ (.A(_19944_),
    .B(_19241_),
    .C(_19242_),
    .Y(_19243_));
 sky130_as_sc_hs__or2_2 _51626_ (.A(net1686),
    .B(_19944_),
    .Y(_19244_));
 sky130_as_sc_hs__and2_2 _51627_ (.A(net504),
    .B(_19244_),
    .Y(_19245_));
 sky130_as_sc_hs__and2_2 _51628_ (.A(_19243_),
    .B(_19245_),
    .Y(_01675_));
 sky130_as_sc_hs__or2_2 _51630_ (.A(\tholin_riscv.PC[24] ),
    .B(net334),
    .Y(_19247_));
 sky130_as_sc_hs__and2_2 _51632_ (.A(_19247_),
    .B(_19248_),
    .Y(_19249_));
 sky130_as_sc_hs__and2_2 _51634_ (.A(_19226_),
    .B(_19250_),
    .Y(_19251_));
 sky130_as_sc_hs__or2_2 _51635_ (.A(_19249_),
    .B(_19251_),
    .Y(_19252_));
 sky130_as_sc_hs__nand3_2 _51637_ (.A(_13046_),
    .B(_19252_),
    .C(_19253_),
    .Y(_19254_));
 sky130_as_sc_hs__nand3_2 _51639_ (.A(_19246_),
    .B(_19254_),
    .C(_19255_),
    .Y(_19256_));
 sky130_as_sc_hs__or2_2 _51641_ (.A(_11911_),
    .B(net125),
    .Y(_19258_));
 sky130_as_sc_hs__nand3_2 _51643_ (.A(net136),
    .B(_19258_),
    .C(_19259_),
    .Y(_19260_));
 sky130_as_sc_hs__nand3_2 _51644_ (.A(_19942_),
    .B(_19257_),
    .C(_19260_),
    .Y(_19261_));
 sky130_as_sc_hs__nand3_2 _51646_ (.A(_19944_),
    .B(_19261_),
    .C(_19262_),
    .Y(_19263_));
 sky130_as_sc_hs__or2_2 _51647_ (.A(net1689),
    .B(_19944_),
    .Y(_19264_));
 sky130_as_sc_hs__and2_2 _51648_ (.A(net504),
    .B(_19264_),
    .Y(_19265_));
 sky130_as_sc_hs__and2_2 _51649_ (.A(_19263_),
    .B(_19265_),
    .Y(_01676_));
 sky130_as_sc_hs__or2_2 _51651_ (.A(\tholin_riscv.PC[25] ),
    .B(net334),
    .Y(_19267_));
 sky130_as_sc_hs__and2_2 _51653_ (.A(_19267_),
    .B(_19268_),
    .Y(_19269_));
 sky130_as_sc_hs__nand3_2 _51654_ (.A(_19228_),
    .B(_19230_),
    .C(_19249_),
    .Y(_19270_));
 sky130_as_sc_hs__and2_2 _51655_ (.A(_19226_),
    .B(_19248_),
    .Y(_19271_));
 sky130_as_sc_hs__nand3_2 _51656_ (.A(_19229_),
    .B(_19270_),
    .C(_19271_),
    .Y(_19272_));
 sky130_as_sc_hs__and2_2 _51657_ (.A(_19269_),
    .B(_19272_),
    .Y(_19273_));
 sky130_as_sc_hs__nor2_2 _51658_ (.A(_19269_),
    .B(_19272_),
    .Y(_19274_));
 sky130_as_sc_hs__or2_2 _51659_ (.A(_19273_),
    .B(_19274_),
    .Y(_19275_));
 sky130_as_sc_hs__nand3_2 _51662_ (.A(_19266_),
    .B(_19276_),
    .C(_19277_),
    .Y(_19278_));
 sky130_as_sc_hs__nand3_2 _51666_ (.A(net136),
    .B(_19280_),
    .C(_19281_),
    .Y(_19282_));
 sky130_as_sc_hs__nand3_2 _51667_ (.A(_19942_),
    .B(_19279_),
    .C(_19282_),
    .Y(_19283_));
 sky130_as_sc_hs__nand3_2 _51669_ (.A(_19944_),
    .B(_19283_),
    .C(_19284_),
    .Y(_19285_));
 sky130_as_sc_hs__or2_2 _51670_ (.A(net1695),
    .B(_19944_),
    .Y(_19286_));
 sky130_as_sc_hs__and2_2 _51671_ (.A(net504),
    .B(_19286_),
    .Y(_19287_));
 sky130_as_sc_hs__and2_2 _51672_ (.A(_19285_),
    .B(_19287_),
    .Y(_01677_));
 sky130_as_sc_hs__or2_2 _51674_ (.A(\tholin_riscv.PC[26] ),
    .B(net334),
    .Y(_19289_));
 sky130_as_sc_hs__and2_2 _51676_ (.A(_19289_),
    .B(_19290_),
    .Y(_19291_));
 sky130_as_sc_hs__and2_2 _51678_ (.A(_19268_),
    .B(_19292_),
    .Y(_19293_));
 sky130_as_sc_hs__or2_2 _51679_ (.A(_19291_),
    .B(_19293_),
    .Y(_19294_));
 sky130_as_sc_hs__nand3_2 _51681_ (.A(_13046_),
    .B(_19294_),
    .C(_19295_),
    .Y(_19296_));
 sky130_as_sc_hs__nand3_2 _51683_ (.A(_19288_),
    .B(_19296_),
    .C(_19297_),
    .Y(_19298_));
 sky130_as_sc_hs__or2_2 _51685_ (.A(_12170_),
    .B(net125),
    .Y(_19300_));
 sky130_as_sc_hs__nand3_2 _51687_ (.A(net136),
    .B(_19300_),
    .C(_19301_),
    .Y(_19302_));
 sky130_as_sc_hs__nand3_2 _51688_ (.A(_19942_),
    .B(_19299_),
    .C(_19302_),
    .Y(_19303_));
 sky130_as_sc_hs__nand3_2 _51690_ (.A(_19944_),
    .B(_19303_),
    .C(_19304_),
    .Y(_19305_));
 sky130_as_sc_hs__or2_2 _51691_ (.A(net1693),
    .B(_19944_),
    .Y(_19306_));
 sky130_as_sc_hs__and2_2 _51692_ (.A(net504),
    .B(_19306_),
    .Y(_19307_));
 sky130_as_sc_hs__and2_2 _51693_ (.A(_19305_),
    .B(_19307_),
    .Y(_01678_));
 sky130_as_sc_hs__or2_2 _51695_ (.A(\tholin_riscv.PC[27] ),
    .B(net334),
    .Y(_19309_));
 sky130_as_sc_hs__inv_2 _51698_ (.Y(_19312_),
    .A(_19311_));
 sky130_as_sc_hs__and2_2 _51699_ (.A(_19273_),
    .B(_19291_),
    .Y(_19313_));
 sky130_as_sc_hs__and2_2 _51700_ (.A(_19268_),
    .B(_19290_),
    .Y(_19314_));
 sky130_as_sc_hs__nand2b_2 _51701_ (.B(_19314_),
    .Y(_19315_),
    .A(_19313_));
 sky130_as_sc_hs__or2_2 _51703_ (.A(_19311_),
    .B(_19315_),
    .Y(_19317_));
 sky130_as_sc_hs__nand3_2 _51704_ (.A(_13046_),
    .B(_19316_),
    .C(_19317_),
    .Y(_19318_));
 sky130_as_sc_hs__nand3_2 _51706_ (.A(_19308_),
    .B(_19318_),
    .C(_19319_),
    .Y(_19320_));
 sky130_as_sc_hs__or2_2 _51708_ (.A(_12291_),
    .B(_13061_),
    .Y(_19322_));
 sky130_as_sc_hs__nand3_2 _51710_ (.A(net136),
    .B(_19322_),
    .C(_19323_),
    .Y(_19324_));
 sky130_as_sc_hs__nand3_2 _51711_ (.A(_19942_),
    .B(_19321_),
    .C(_19324_),
    .Y(_19325_));
 sky130_as_sc_hs__nand3_2 _51713_ (.A(_19944_),
    .B(_19325_),
    .C(_19326_),
    .Y(_19327_));
 sky130_as_sc_hs__or2_2 _51714_ (.A(net1683),
    .B(_19944_),
    .Y(_19328_));
 sky130_as_sc_hs__and2_2 _51715_ (.A(net503),
    .B(_19328_),
    .Y(_19329_));
 sky130_as_sc_hs__and2_2 _51716_ (.A(_19327_),
    .B(_19329_),
    .Y(_01679_));
 sky130_as_sc_hs__or2_2 _51718_ (.A(\tholin_riscv.PC[28] ),
    .B(\tholin_riscv.Bimm[12] ),
    .Y(_19331_));
 sky130_as_sc_hs__and2_2 _51720_ (.A(_19331_),
    .B(_19332_),
    .Y(_19333_));
 sky130_as_sc_hs__and2_2 _51722_ (.A(_19310_),
    .B(_19334_),
    .Y(_19335_));
 sky130_as_sc_hs__or2_2 _51723_ (.A(_19333_),
    .B(_19335_),
    .Y(_19336_));
 sky130_as_sc_hs__nand3_2 _51725_ (.A(_13046_),
    .B(_19336_),
    .C(_19337_),
    .Y(_19338_));
 sky130_as_sc_hs__nand3_2 _51727_ (.A(_19330_),
    .B(_19338_),
    .C(_19339_),
    .Y(_19340_));
 sky130_as_sc_hs__or2_2 _51729_ (.A(_12403_),
    .B(net125),
    .Y(_19342_));
 sky130_as_sc_hs__nand3_2 _51731_ (.A(net136),
    .B(_19342_),
    .C(_19343_),
    .Y(_19344_));
 sky130_as_sc_hs__nand3_2 _51732_ (.A(_19942_),
    .B(_19341_),
    .C(_19344_),
    .Y(_19345_));
 sky130_as_sc_hs__nand3_2 _51734_ (.A(_19944_),
    .B(_19345_),
    .C(_19346_),
    .Y(_19347_));
 sky130_as_sc_hs__or2_2 _51735_ (.A(net1696),
    .B(_19944_),
    .Y(_19348_));
 sky130_as_sc_hs__and2_2 _51736_ (.A(net504),
    .B(_19348_),
    .Y(_19349_));
 sky130_as_sc_hs__and2_2 _51737_ (.A(_19347_),
    .B(_19349_),
    .Y(_01680_));
 sky130_as_sc_hs__or2_2 _51739_ (.A(\tholin_riscv.PC[29] ),
    .B(\tholin_riscv.Bimm[12] ),
    .Y(_19351_));
 sky130_as_sc_hs__and2_2 _51741_ (.A(_19351_),
    .B(_19352_),
    .Y(_19353_));
 sky130_as_sc_hs__nand3_2 _51742_ (.A(_19312_),
    .B(_19313_),
    .C(_19333_),
    .Y(_19354_));
 sky130_as_sc_hs__and2_2 _51743_ (.A(_19310_),
    .B(_19332_),
    .Y(_19355_));
 sky130_as_sc_hs__nand3_2 _51744_ (.A(_19314_),
    .B(_19354_),
    .C(_19355_),
    .Y(_19356_));
 sky130_as_sc_hs__and2_2 _51745_ (.A(_19353_),
    .B(_19356_),
    .Y(_19357_));
 sky130_as_sc_hs__nor2_2 _51746_ (.A(_19353_),
    .B(_19356_),
    .Y(_19358_));
 sky130_as_sc_hs__or2_2 _51747_ (.A(_19357_),
    .B(_19358_),
    .Y(_19359_));
 sky130_as_sc_hs__nand3_2 _51750_ (.A(_19350_),
    .B(_19360_),
    .C(_19361_),
    .Y(_19362_));
 sky130_as_sc_hs__or2_2 _51752_ (.A(_12499_),
    .B(net125),
    .Y(_19364_));
 sky130_as_sc_hs__nand3_2 _51754_ (.A(net136),
    .B(_19364_),
    .C(_19365_),
    .Y(_19366_));
 sky130_as_sc_hs__nand3_2 _51755_ (.A(_19942_),
    .B(_19363_),
    .C(_19366_),
    .Y(_19367_));
 sky130_as_sc_hs__nand3_2 _51757_ (.A(_19944_),
    .B(_19367_),
    .C(_19368_),
    .Y(_19369_));
 sky130_as_sc_hs__or2_2 _51758_ (.A(net1697),
    .B(_19944_),
    .Y(_19370_));
 sky130_as_sc_hs__and2_2 _51759_ (.A(net504),
    .B(_19370_),
    .Y(_19371_));
 sky130_as_sc_hs__and2_2 _51760_ (.A(_19369_),
    .B(_19371_),
    .Y(_01681_));
 sky130_as_sc_hs__or2_2 _51763_ (.A(\tholin_riscv.PC[30] ),
    .B(net334),
    .Y(_19374_));
 sky130_as_sc_hs__and2_2 _51765_ (.A(_19374_),
    .B(_19375_),
    .Y(_19376_));
 sky130_as_sc_hs__or2_2 _51769_ (.A(_19376_),
    .B(_19378_),
    .Y(_19380_));
 sky130_as_sc_hs__nand3_2 _51770_ (.A(_13046_),
    .B(_19379_),
    .C(_19380_),
    .Y(_19381_));
 sky130_as_sc_hs__and2_2 _51772_ (.A(_19990_),
    .B(_19382_),
    .Y(_19383_));
 sky130_as_sc_hs__nand3_2 _51773_ (.A(_19373_),
    .B(_19381_),
    .C(_19383_),
    .Y(_19384_));
 sky130_as_sc_hs__nand3_2 _51776_ (.A(net136),
    .B(_19385_),
    .C(_19386_),
    .Y(_19387_));
 sky130_as_sc_hs__nand3_2 _51777_ (.A(net145),
    .B(_19384_),
    .C(_19387_),
    .Y(_19388_));
 sky130_as_sc_hs__and2_2 _51779_ (.A(net501),
    .B(_19389_),
    .Y(_01682_));
 sky130_as_sc_hs__nand3_2 _51782_ (.A(_19352_),
    .B(_19375_),
    .C(_19391_),
    .Y(_19392_));
 sky130_as_sc_hs__or2_2 _51784_ (.A(_12661_),
    .B(_19392_),
    .Y(_19394_));
 sky130_as_sc_hs__nand3_2 _51785_ (.A(_13046_),
    .B(_19393_),
    .C(_19394_),
    .Y(_19395_));
 sky130_as_sc_hs__or2_2 _51787_ (.A(_12620_),
    .B(_13065_),
    .Y(_19397_));
 sky130_as_sc_hs__and2_2 _51788_ (.A(_19990_),
    .B(_19397_),
    .Y(_19398_));
 sky130_as_sc_hs__nand3_2 _51789_ (.A(_19395_),
    .B(_19396_),
    .C(_19398_),
    .Y(_19399_));
 sky130_as_sc_hs__nand3_2 _51792_ (.A(net136),
    .B(_19400_),
    .C(_19401_),
    .Y(_19402_));
 sky130_as_sc_hs__nand3_2 _51793_ (.A(net145),
    .B(_19399_),
    .C(_19402_),
    .Y(_19403_));
 sky130_as_sc_hs__and2_2 _51795_ (.A(net501),
    .B(_19404_),
    .Y(_01683_));
 sky130_as_sc_hs__and2_2 _51796_ (.A(_21560_),
    .B(_13146_),
    .Y(_19405_));
 sky130_as_sc_hs__or2_2 _51799_ (.A(net669),
    .B(_19405_),
    .Y(_19408_));
 sky130_as_sc_hs__and2_2 _51800_ (.A(_19407_),
    .B(net670),
    .Y(_01689_));
 sky130_as_sc_hs__and2_2 _51894_ (.A(net524),
    .B(_16551_),
    .Y(_01684_));
 sky130_as_sc_hs__and2_2 _51895_ (.A(_16570_),
    .B(_16572_),
    .Y(_01685_));
 sky130_as_sc_hs__and2_2 _51896_ (.A(net520),
    .B(_16593_),
    .Y(_01686_));
 sky130_as_sc_hs__and2_2 _51897_ (.A(_16612_),
    .B(_16614_),
    .Y(_01687_));
 sky130_as_sc_hs__and2_2 _51898_ (.A(_16633_),
    .B(_16635_),
    .Y(_01688_));
 sky130_as_sc_hs__dfxtp_2 _51899_ (.CLK(clknet_leaf_203_wb_clk_i),
    .Q(\tholin_riscv.Bimm[1] ),
    .D(_00005_));
 sky130_as_sc_hs__dfxtp_2 _51900_ (.CLK(clknet_leaf_1_wb_clk_i),
    .Q(\tholin_riscv.Bimm[2] ),
    .D(_00006_));
 sky130_as_sc_hs__dfxtp_2 _51901_ (.CLK(clknet_leaf_203_wb_clk_i),
    .Q(\tholin_riscv.Bimm[3] ),
    .D(_00007_));
 sky130_as_sc_hs__dfxtp_2 _51902_ (.CLK(clknet_leaf_191_wb_clk_i),
    .Q(\tholin_riscv.Bimm[4] ),
    .D(_00008_));
 sky130_as_sc_hs__dfxtp_2 _51903_ (.CLK(clknet_leaf_203_wb_clk_i),
    .Q(\tholin_riscv.Jimm[12] ),
    .D(_00009_));
 sky130_as_sc_hs__dfxtp_2 _51904_ (.CLK(clknet_leaf_1_wb_clk_i),
    .Q(\tholin_riscv.Jimm[13] ),
    .D(_00010_));
 sky130_as_sc_hs__dfxtp_2 _51905_ (.CLK(clknet_leaf_1_wb_clk_i),
    .Q(\tholin_riscv.Jimm[14] ),
    .D(_00011_));
 sky130_as_sc_hs__dfxtp_2 _51906_ (.CLK(clknet_leaf_1_wb_clk_i),
    .Q(\tholin_riscv.Jimm[15] ),
    .D(_00012_));
 sky130_as_sc_hs__dfxtp_2 _51907_ (.CLK(clknet_leaf_187_wb_clk_i),
    .Q(\tholin_riscv.instr[0] ),
    .D(_00013_));
 sky130_as_sc_hs__dfxtp_2 _51908_ (.CLK(clknet_leaf_189_wb_clk_i),
    .Q(\tholin_riscv.instr[1] ),
    .D(_00014_));
 sky130_as_sc_hs__dfxtp_2 _51909_ (.CLK(clknet_leaf_190_wb_clk_i),
    .Q(\tholin_riscv.instr[2] ),
    .D(_00015_));
 sky130_as_sc_hs__dfxtp_2 _51910_ (.CLK(clknet_leaf_189_wb_clk_i),
    .Q(\tholin_riscv.instr[3] ),
    .D(_00016_));
 sky130_as_sc_hs__dfxtp_2 _51911_ (.CLK(clknet_leaf_189_wb_clk_i),
    .Q(\tholin_riscv.instr[4] ),
    .D(_00017_));
 sky130_as_sc_hs__dfxtp_2 _51912_ (.CLK(clknet_leaf_189_wb_clk_i),
    .Q(\tholin_riscv.instr[5] ),
    .D(_00018_));
 sky130_as_sc_hs__dfxtp_2 _51913_ (.CLK(clknet_leaf_190_wb_clk_i),
    .Q(\tholin_riscv.instr[6] ),
    .D(net1430));
 sky130_as_sc_hs__dfxtp_2 _51914_ (.CLK(clknet_leaf_188_wb_clk_i),
    .Q(\tholin_riscv.Bimm[11] ),
    .D(_00020_));
 sky130_as_sc_hs__dfxtp_2 _51915_ (.CLK(clknet_leaf_132_wb_clk_i),
    .Q(\tholin_riscv.regs[31][0] ),
    .D(net737));
 sky130_as_sc_hs__dfxtp_2 _51916_ (.CLK(clknet_leaf_126_wb_clk_i),
    .Q(\tholin_riscv.regs[31][1] ),
    .D(_00022_));
 sky130_as_sc_hs__dfxtp_2 _51917_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[31][2] ),
    .D(_00023_));
 sky130_as_sc_hs__dfxtp_2 _51918_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[31][3] ),
    .D(_00024_));
 sky130_as_sc_hs__dfxtp_2 _51919_ (.CLK(clknet_leaf_111_wb_clk_i),
    .Q(\tholin_riscv.regs[31][4] ),
    .D(_00025_));
 sky130_as_sc_hs__dfxtp_2 _51920_ (.CLK(clknet_leaf_54_wb_clk_i),
    .Q(\tholin_riscv.regs[31][5] ),
    .D(_00026_));
 sky130_as_sc_hs__dfxtp_2 _51921_ (.CLK(clknet_leaf_62_wb_clk_i),
    .Q(\tholin_riscv.regs[31][6] ),
    .D(_00027_));
 sky130_as_sc_hs__dfxtp_2 _51922_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[31][7] ),
    .D(_00028_));
 sky130_as_sc_hs__dfxtp_2 _51923_ (.CLK(clknet_leaf_80_wb_clk_i),
    .Q(\tholin_riscv.regs[31][8] ),
    .D(_00029_));
 sky130_as_sc_hs__dfxtp_2 _51924_ (.CLK(clknet_leaf_44_wb_clk_i),
    .Q(\tholin_riscv.regs[31][9] ),
    .D(_00030_));
 sky130_as_sc_hs__dfxtp_2 _51925_ (.CLK(clknet_leaf_42_wb_clk_i),
    .Q(\tholin_riscv.regs[31][10] ),
    .D(_00031_));
 sky130_as_sc_hs__dfxtp_2 _51926_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[31][11] ),
    .D(_00032_));
 sky130_as_sc_hs__dfxtp_2 _51927_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[31][12] ),
    .D(_00033_));
 sky130_as_sc_hs__dfxtp_2 _51928_ (.CLK(clknet_leaf_29_wb_clk_i),
    .Q(\tholin_riscv.regs[31][13] ),
    .D(_00034_));
 sky130_as_sc_hs__dfxtp_2 _51929_ (.CLK(clknet_leaf_19_wb_clk_i),
    .Q(\tholin_riscv.regs[31][14] ),
    .D(_00035_));
 sky130_as_sc_hs__dfxtp_2 _51930_ (.CLK(clknet_leaf_18_wb_clk_i),
    .Q(\tholin_riscv.regs[31][15] ),
    .D(_00036_));
 sky130_as_sc_hs__dfxtp_2 _51931_ (.CLK(clknet_leaf_103_wb_clk_i),
    .Q(\tholin_riscv.regs[31][16] ),
    .D(_00037_));
 sky130_as_sc_hs__dfxtp_2 _51932_ (.CLK(clknet_leaf_147_wb_clk_i),
    .Q(\tholin_riscv.regs[31][17] ),
    .D(_00038_));
 sky130_as_sc_hs__dfxtp_2 _51933_ (.CLK(clknet_leaf_115_wb_clk_i),
    .Q(\tholin_riscv.regs[31][18] ),
    .D(_00039_));
 sky130_as_sc_hs__dfxtp_2 _51934_ (.CLK(clknet_leaf_114_wb_clk_i),
    .Q(\tholin_riscv.regs[31][19] ),
    .D(_00040_));
 sky130_as_sc_hs__dfxtp_2 _51935_ (.CLK(clknet_leaf_113_wb_clk_i),
    .Q(\tholin_riscv.regs[31][20] ),
    .D(_00041_));
 sky130_as_sc_hs__dfxtp_2 _51936_ (.CLK(clknet_leaf_118_wb_clk_i),
    .Q(\tholin_riscv.regs[31][21] ),
    .D(_00042_));
 sky130_as_sc_hs__dfxtp_2 _51937_ (.CLK(clknet_leaf_107_wb_clk_i),
    .Q(\tholin_riscv.regs[31][22] ),
    .D(_00043_));
 sky130_as_sc_hs__dfxtp_2 _51938_ (.CLK(clknet_leaf_106_wb_clk_i),
    .Q(\tholin_riscv.regs[31][23] ),
    .D(_00044_));
 sky130_as_sc_hs__dfxtp_2 _51939_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[31][24] ),
    .D(_00045_));
 sky130_as_sc_hs__dfxtp_2 _51940_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[31][25] ),
    .D(_00046_));
 sky130_as_sc_hs__dfxtp_2 _51941_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[31][26] ),
    .D(_00047_));
 sky130_as_sc_hs__dfxtp_2 _51942_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[31][27] ),
    .D(_00048_));
 sky130_as_sc_hs__dfxtp_2 _51943_ (.CLK(clknet_leaf_91_wb_clk_i),
    .Q(\tholin_riscv.regs[31][28] ),
    .D(_00049_));
 sky130_as_sc_hs__dfxtp_2 _51944_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[31][29] ),
    .D(_00050_));
 sky130_as_sc_hs__dfxtp_2 _51945_ (.CLK(clknet_leaf_99_wb_clk_i),
    .Q(\tholin_riscv.regs[31][30] ),
    .D(_00051_));
 sky130_as_sc_hs__dfxtp_2 _51946_ (.CLK(clknet_leaf_150_wb_clk_i),
    .Q(\tholin_riscv.regs[31][31] ),
    .D(_00052_));
 sky130_as_sc_hs__dfxtp_2 _51947_ (.CLK(clknet_leaf_131_wb_clk_i),
    .Q(\tholin_riscv.regs[16][0] ),
    .D(net713));
 sky130_as_sc_hs__dfxtp_2 _51948_ (.CLK(clknet_leaf_127_wb_clk_i),
    .Q(\tholin_riscv.regs[16][1] ),
    .D(_00054_));
 sky130_as_sc_hs__dfxtp_2 _51949_ (.CLK(clknet_leaf_8_wb_clk_i),
    .Q(\tholin_riscv.regs[16][2] ),
    .D(_00055_));
 sky130_as_sc_hs__dfxtp_2 _51950_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[16][3] ),
    .D(_00056_));
 sky130_as_sc_hs__dfxtp_2 _51951_ (.CLK(clknet_leaf_69_wb_clk_i),
    .Q(\tholin_riscv.regs[16][4] ),
    .D(_00057_));
 sky130_as_sc_hs__dfxtp_2 _51952_ (.CLK(clknet_leaf_57_wb_clk_i),
    .Q(\tholin_riscv.regs[16][5] ),
    .D(_00058_));
 sky130_as_sc_hs__dfxtp_2 _51953_ (.CLK(clknet_leaf_62_wb_clk_i),
    .Q(\tholin_riscv.regs[16][6] ),
    .D(_00059_));
 sky130_as_sc_hs__dfxtp_2 _51954_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[16][7] ),
    .D(_00060_));
 sky130_as_sc_hs__dfxtp_2 _51955_ (.CLK(clknet_leaf_80_wb_clk_i),
    .Q(\tholin_riscv.regs[16][8] ),
    .D(_00061_));
 sky130_as_sc_hs__dfxtp_2 _51956_ (.CLK(clknet_leaf_38_wb_clk_i),
    .Q(\tholin_riscv.regs[16][9] ),
    .D(_00062_));
 sky130_as_sc_hs__dfxtp_2 _51957_ (.CLK(clknet_leaf_31_wb_clk_i),
    .Q(\tholin_riscv.regs[16][10] ),
    .D(_00063_));
 sky130_as_sc_hs__dfxtp_2 _51958_ (.CLK(clknet_leaf_29_wb_clk_i),
    .Q(\tholin_riscv.regs[16][11] ),
    .D(_00064_));
 sky130_as_sc_hs__dfxtp_2 _51959_ (.CLK(clknet_leaf_27_wb_clk_i),
    .Q(\tholin_riscv.regs[16][12] ),
    .D(_00065_));
 sky130_as_sc_hs__dfxtp_2 _51960_ (.CLK(clknet_leaf_22_wb_clk_i),
    .Q(\tholin_riscv.regs[16][13] ),
    .D(_00066_));
 sky130_as_sc_hs__dfxtp_2 _51961_ (.CLK(clknet_leaf_18_wb_clk_i),
    .Q(\tholin_riscv.regs[16][14] ),
    .D(_00067_));
 sky130_as_sc_hs__dfxtp_2 _51962_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[16][15] ),
    .D(_00068_));
 sky130_as_sc_hs__dfxtp_2 _51963_ (.CLK(clknet_leaf_78_wb_clk_i),
    .Q(\tholin_riscv.regs[16][16] ),
    .D(_00069_));
 sky130_as_sc_hs__dfxtp_2 _51964_ (.CLK(clknet_leaf_78_wb_clk_i),
    .Q(\tholin_riscv.regs[16][17] ),
    .D(_00070_));
 sky130_as_sc_hs__dfxtp_2 _51965_ (.CLK(clknet_leaf_73_wb_clk_i),
    .Q(\tholin_riscv.regs[16][18] ),
    .D(_00071_));
 sky130_as_sc_hs__dfxtp_2 _51966_ (.CLK(clknet_leaf_74_wb_clk_i),
    .Q(\tholin_riscv.regs[16][19] ),
    .D(_00072_));
 sky130_as_sc_hs__dfxtp_2 _51967_ (.CLK(clknet_leaf_73_wb_clk_i),
    .Q(\tholin_riscv.regs[16][20] ),
    .D(_00073_));
 sky130_as_sc_hs__dfxtp_2 _51968_ (.CLK(clknet_leaf_81_wb_clk_i),
    .Q(\tholin_riscv.regs[16][21] ),
    .D(_00074_));
 sky130_as_sc_hs__dfxtp_2 _51969_ (.CLK(clknet_leaf_123_wb_clk_i),
    .Q(\tholin_riscv.regs[16][22] ),
    .D(_00075_));
 sky130_as_sc_hs__dfxtp_2 _51970_ (.CLK(clknet_leaf_66_wb_clk_i),
    .Q(\tholin_riscv.regs[16][23] ),
    .D(_00076_));
 sky130_as_sc_hs__dfxtp_2 _51971_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[16][24] ),
    .D(_00077_));
 sky130_as_sc_hs__dfxtp_2 _51972_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[16][25] ),
    .D(_00078_));
 sky130_as_sc_hs__dfxtp_2 _51973_ (.CLK(clknet_leaf_89_wb_clk_i),
    .Q(\tholin_riscv.regs[16][26] ),
    .D(_00079_));
 sky130_as_sc_hs__dfxtp_2 _51974_ (.CLK(clknet_leaf_90_wb_clk_i),
    .Q(\tholin_riscv.regs[16][27] ),
    .D(_00080_));
 sky130_as_sc_hs__dfxtp_2 _51975_ (.CLK(clknet_leaf_89_wb_clk_i),
    .Q(\tholin_riscv.regs[16][28] ),
    .D(_00081_));
 sky130_as_sc_hs__dfxtp_2 _51976_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[16][29] ),
    .D(_00082_));
 sky130_as_sc_hs__dfxtp_2 _51977_ (.CLK(clknet_leaf_116_wb_clk_i),
    .Q(\tholin_riscv.regs[16][30] ),
    .D(_00083_));
 sky130_as_sc_hs__dfxtp_2 _51978_ (.CLK(clknet_leaf_121_wb_clk_i),
    .Q(\tholin_riscv.regs[16][31] ),
    .D(_00084_));
 sky130_as_sc_hs__dfxtp_2 _51979_ (.CLK(clknet_leaf_133_wb_clk_i),
    .Q(\tholin_riscv.regs[14][0] ),
    .D(net740));
 sky130_as_sc_hs__dfxtp_2 _51980_ (.CLK(clknet_leaf_128_wb_clk_i),
    .Q(\tholin_riscv.regs[14][1] ),
    .D(_00086_));
 sky130_as_sc_hs__dfxtp_2 _51981_ (.CLK(clknet_leaf_64_wb_clk_i),
    .Q(\tholin_riscv.regs[14][2] ),
    .D(_00087_));
 sky130_as_sc_hs__dfxtp_2 _51982_ (.CLK(clknet_leaf_62_wb_clk_i),
    .Q(\tholin_riscv.regs[14][3] ),
    .D(_00088_));
 sky130_as_sc_hs__dfxtp_2 _51983_ (.CLK(clknet_leaf_71_wb_clk_i),
    .Q(\tholin_riscv.regs[14][4] ),
    .D(_00089_));
 sky130_as_sc_hs__dfxtp_2 _51984_ (.CLK(clknet_leaf_59_wb_clk_i),
    .Q(\tholin_riscv.regs[14][5] ),
    .D(_00090_));
 sky130_as_sc_hs__dfxtp_2 _51985_ (.CLK(clknet_leaf_61_wb_clk_i),
    .Q(\tholin_riscv.regs[14][6] ),
    .D(_00091_));
 sky130_as_sc_hs__dfxtp_2 _51986_ (.CLK(clknet_leaf_47_wb_clk_i),
    .Q(\tholin_riscv.regs[14][7] ),
    .D(_00092_));
 sky130_as_sc_hs__dfxtp_2 _51987_ (.CLK(clknet_leaf_84_wb_clk_i),
    .Q(\tholin_riscv.regs[14][8] ),
    .D(_00093_));
 sky130_as_sc_hs__dfxtp_2 _51988_ (.CLK(clknet_leaf_83_wb_clk_i),
    .Q(\tholin_riscv.regs[14][9] ),
    .D(_00094_));
 sky130_as_sc_hs__dfxtp_2 _51989_ (.CLK(clknet_leaf_48_wb_clk_i),
    .Q(\tholin_riscv.regs[14][10] ),
    .D(_00095_));
 sky130_as_sc_hs__dfxtp_2 _51990_ (.CLK(clknet_leaf_49_wb_clk_i),
    .Q(\tholin_riscv.regs[14][11] ),
    .D(_00096_));
 sky130_as_sc_hs__dfxtp_2 _51991_ (.CLK(clknet_leaf_32_wb_clk_i),
    .Q(\tholin_riscv.regs[14][12] ),
    .D(_00097_));
 sky130_as_sc_hs__dfxtp_2 _51992_ (.CLK(clknet_leaf_25_wb_clk_i),
    .Q(\tholin_riscv.regs[14][13] ),
    .D(_00098_));
 sky130_as_sc_hs__dfxtp_2 _51993_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[14][14] ),
    .D(_00099_));
 sky130_as_sc_hs__dfxtp_2 _51994_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[14][15] ),
    .D(_00100_));
 sky130_as_sc_hs__dfxtp_2 _51995_ (.CLK(clknet_leaf_89_wb_clk_i),
    .Q(\tholin_riscv.regs[14][16] ),
    .D(_00101_));
 sky130_as_sc_hs__dfxtp_2 _51996_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[14][17] ),
    .D(_00102_));
 sky130_as_sc_hs__dfxtp_2 _51997_ (.CLK(clknet_leaf_82_wb_clk_i),
    .Q(\tholin_riscv.regs[14][18] ),
    .D(_00103_));
 sky130_as_sc_hs__dfxtp_2 _51998_ (.CLK(clknet_leaf_60_wb_clk_i),
    .Q(\tholin_riscv.regs[14][19] ),
    .D(_00104_));
 sky130_as_sc_hs__dfxtp_2 _51999_ (.CLK(clknet_leaf_73_wb_clk_i),
    .Q(\tholin_riscv.regs[14][20] ),
    .D(_00105_));
 sky130_as_sc_hs__dfxtp_2 _52000_ (.CLK(clknet_leaf_86_wb_clk_i),
    .Q(\tholin_riscv.regs[14][21] ),
    .D(_00106_));
 sky130_as_sc_hs__dfxtp_2 _52001_ (.CLK(clknet_leaf_71_wb_clk_i),
    .Q(\tholin_riscv.regs[14][22] ),
    .D(_00107_));
 sky130_as_sc_hs__dfxtp_2 _52002_ (.CLK(clknet_leaf_68_wb_clk_i),
    .Q(\tholin_riscv.regs[14][23] ),
    .D(_00108_));
 sky130_as_sc_hs__dfxtp_2 _52003_ (.CLK(clknet_leaf_35_wb_clk_i),
    .Q(\tholin_riscv.regs[14][24] ),
    .D(_00109_));
 sky130_as_sc_hs__dfxtp_2 _52004_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[14][25] ),
    .D(_00110_));
 sky130_as_sc_hs__dfxtp_2 _52005_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[14][26] ),
    .D(_00111_));
 sky130_as_sc_hs__dfxtp_2 _52006_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[14][27] ),
    .D(_00112_));
 sky130_as_sc_hs__dfxtp_2 _52007_ (.CLK(clknet_leaf_23_wb_clk_i),
    .Q(\tholin_riscv.regs[14][28] ),
    .D(_00113_));
 sky130_as_sc_hs__dfxtp_2 _52008_ (.CLK(clknet_leaf_38_wb_clk_i),
    .Q(\tholin_riscv.regs[14][29] ),
    .D(_00114_));
 sky130_as_sc_hs__dfxtp_2 _52009_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.regs[14][30] ),
    .D(_00115_));
 sky130_as_sc_hs__dfxtp_2 _52010_ (.CLK(clknet_leaf_113_wb_clk_i),
    .Q(\tholin_riscv.regs[14][31] ),
    .D(_00116_));
 sky130_as_sc_hs__dfxtp_2 _52011_ (.CLK(clknet_leaf_130_wb_clk_i),
    .Q(\tholin_riscv.regs[11][0] ),
    .D(net692));
 sky130_as_sc_hs__dfxtp_2 _52012_ (.CLK(clknet_leaf_68_wb_clk_i),
    .Q(\tholin_riscv.regs[11][1] ),
    .D(_00118_));
 sky130_as_sc_hs__dfxtp_2 _52013_ (.CLK(clknet_leaf_66_wb_clk_i),
    .Q(\tholin_riscv.regs[11][2] ),
    .D(_00119_));
 sky130_as_sc_hs__dfxtp_2 _52014_ (.CLK(clknet_leaf_55_wb_clk_i),
    .Q(\tholin_riscv.regs[11][3] ),
    .D(_00120_));
 sky130_as_sc_hs__dfxtp_2 _52015_ (.CLK(clknet_leaf_103_wb_clk_i),
    .Q(\tholin_riscv.regs[11][4] ),
    .D(_00121_));
 sky130_as_sc_hs__dfxtp_2 _52016_ (.CLK(clknet_leaf_59_wb_clk_i),
    .Q(\tholin_riscv.regs[11][5] ),
    .D(_00122_));
 sky130_as_sc_hs__dfxtp_2 _52017_ (.CLK(clknet_leaf_64_wb_clk_i),
    .Q(\tholin_riscv.regs[11][6] ),
    .D(_00123_));
 sky130_as_sc_hs__dfxtp_2 _52018_ (.CLK(clknet_leaf_58_wb_clk_i),
    .Q(\tholin_riscv.regs[11][7] ),
    .D(_00124_));
 sky130_as_sc_hs__dfxtp_2 _52019_ (.CLK(clknet_leaf_83_wb_clk_i),
    .Q(\tholin_riscv.regs[11][8] ),
    .D(_00125_));
 sky130_as_sc_hs__dfxtp_2 _52020_ (.CLK(clknet_leaf_44_wb_clk_i),
    .Q(\tholin_riscv.regs[11][9] ),
    .D(_00126_));
 sky130_as_sc_hs__dfxtp_2 _52021_ (.CLK(clknet_leaf_50_wb_clk_i),
    .Q(\tholin_riscv.regs[11][10] ),
    .D(_00127_));
 sky130_as_sc_hs__dfxtp_2 _52022_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[11][11] ),
    .D(_00128_));
 sky130_as_sc_hs__dfxtp_2 _52023_ (.CLK(clknet_leaf_31_wb_clk_i),
    .Q(\tholin_riscv.regs[11][12] ),
    .D(_00129_));
 sky130_as_sc_hs__dfxtp_2 _52024_ (.CLK(clknet_leaf_28_wb_clk_i),
    .Q(\tholin_riscv.regs[11][13] ),
    .D(_00130_));
 sky130_as_sc_hs__dfxtp_2 _52025_ (.CLK(clknet_leaf_14_wb_clk_i),
    .Q(\tholin_riscv.regs[11][14] ),
    .D(_00131_));
 sky130_as_sc_hs__dfxtp_2 _52026_ (.CLK(clknet_leaf_15_wb_clk_i),
    .Q(\tholin_riscv.regs[11][15] ),
    .D(_00132_));
 sky130_as_sc_hs__dfxtp_2 _52027_ (.CLK(clknet_leaf_118_wb_clk_i),
    .Q(\tholin_riscv.regs[11][16] ),
    .D(_00133_));
 sky130_as_sc_hs__dfxtp_2 _52028_ (.CLK(clknet_leaf_101_wb_clk_i),
    .Q(\tholin_riscv.regs[11][17] ),
    .D(_00134_));
 sky130_as_sc_hs__dfxtp_2 _52029_ (.CLK(clknet_leaf_104_wb_clk_i),
    .Q(\tholin_riscv.regs[11][18] ),
    .D(_00135_));
 sky130_as_sc_hs__dfxtp_2 _52030_ (.CLK(clknet_leaf_108_wb_clk_i),
    .Q(\tholin_riscv.regs[11][19] ),
    .D(_00136_));
 sky130_as_sc_hs__dfxtp_2 _52031_ (.CLK(clknet_leaf_109_wb_clk_i),
    .Q(\tholin_riscv.regs[11][20] ),
    .D(_00137_));
 sky130_as_sc_hs__dfxtp_2 _52032_ (.CLK(clknet_leaf_100_wb_clk_i),
    .Q(\tholin_riscv.regs[11][21] ),
    .D(_00138_));
 sky130_as_sc_hs__dfxtp_2 _52033_ (.CLK(clknet_leaf_77_wb_clk_i),
    .Q(\tholin_riscv.regs[11][22] ),
    .D(_00139_));
 sky130_as_sc_hs__dfxtp_2 _52034_ (.CLK(clknet_leaf_102_wb_clk_i),
    .Q(\tholin_riscv.regs[11][23] ),
    .D(_00140_));
 sky130_as_sc_hs__dfxtp_2 _52035_ (.CLK(clknet_leaf_32_wb_clk_i),
    .Q(\tholin_riscv.regs[11][24] ),
    .D(_00141_));
 sky130_as_sc_hs__dfxtp_2 _52036_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[11][25] ),
    .D(_00142_));
 sky130_as_sc_hs__dfxtp_2 _52037_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[11][26] ),
    .D(_00143_));
 sky130_as_sc_hs__dfxtp_2 _52038_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[11][27] ),
    .D(_00144_));
 sky130_as_sc_hs__dfxtp_2 _52039_ (.CLK(clknet_leaf_23_wb_clk_i),
    .Q(\tholin_riscv.regs[11][28] ),
    .D(_00145_));
 sky130_as_sc_hs__dfxtp_2 _52040_ (.CLK(clknet_leaf_36_wb_clk_i),
    .Q(\tholin_riscv.regs[11][29] ),
    .D(_00146_));
 sky130_as_sc_hs__dfxtp_2 _52041_ (.CLK(clknet_leaf_120_wb_clk_i),
    .Q(\tholin_riscv.regs[11][30] ),
    .D(_00147_));
 sky130_as_sc_hs__dfxtp_2 _52042_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.regs[11][31] ),
    .D(_00148_));
 sky130_as_sc_hs__dfxtp_2 _52043_ (.CLK(clknet_leaf_130_wb_clk_i),
    .Q(\tholin_riscv.regs[8][0] ),
    .D(net704));
 sky130_as_sc_hs__dfxtp_2 _52044_ (.CLK(clknet_leaf_128_wb_clk_i),
    .Q(\tholin_riscv.regs[8][1] ),
    .D(_00150_));
 sky130_as_sc_hs__dfxtp_2 _52045_ (.CLK(clknet_leaf_64_wb_clk_i),
    .Q(\tholin_riscv.regs[8][2] ),
    .D(_00151_));
 sky130_as_sc_hs__dfxtp_2 _52046_ (.CLK(clknet_leaf_55_wb_clk_i),
    .Q(\tholin_riscv.regs[8][3] ),
    .D(_00152_));
 sky130_as_sc_hs__dfxtp_2 _52047_ (.CLK(clknet_leaf_69_wb_clk_i),
    .Q(\tholin_riscv.regs[8][4] ),
    .D(_00153_));
 sky130_as_sc_hs__dfxtp_2 _52048_ (.CLK(clknet_leaf_59_wb_clk_i),
    .Q(\tholin_riscv.regs[8][5] ),
    .D(_00154_));
 sky130_as_sc_hs__dfxtp_2 _52049_ (.CLK(clknet_leaf_61_wb_clk_i),
    .Q(\tholin_riscv.regs[8][6] ),
    .D(_00155_));
 sky130_as_sc_hs__dfxtp_2 _52050_ (.CLK(clknet_leaf_54_wb_clk_i),
    .Q(\tholin_riscv.regs[8][7] ),
    .D(_00156_));
 sky130_as_sc_hs__dfxtp_2 _52051_ (.CLK(clknet_leaf_83_wb_clk_i),
    .Q(\tholin_riscv.regs[8][8] ),
    .D(_00157_));
 sky130_as_sc_hs__dfxtp_2 _52052_ (.CLK(clknet_leaf_44_wb_clk_i),
    .Q(\tholin_riscv.regs[8][9] ),
    .D(_00158_));
 sky130_as_sc_hs__dfxtp_2 _52053_ (.CLK(clknet_leaf_47_wb_clk_i),
    .Q(\tholin_riscv.regs[8][10] ),
    .D(_00159_));
 sky130_as_sc_hs__dfxtp_2 _52054_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[8][11] ),
    .D(_00160_));
 sky130_as_sc_hs__dfxtp_2 _52055_ (.CLK(clknet_leaf_32_wb_clk_i),
    .Q(\tholin_riscv.regs[8][12] ),
    .D(_00161_));
 sky130_as_sc_hs__dfxtp_2 _52056_ (.CLK(clknet_leaf_25_wb_clk_i),
    .Q(\tholin_riscv.regs[8][13] ),
    .D(_00162_));
 sky130_as_sc_hs__dfxtp_2 _52057_ (.CLK(clknet_leaf_14_wb_clk_i),
    .Q(\tholin_riscv.regs[8][14] ),
    .D(_00163_));
 sky130_as_sc_hs__dfxtp_2 _52058_ (.CLK(clknet_leaf_16_wb_clk_i),
    .Q(\tholin_riscv.regs[8][15] ),
    .D(_00164_));
 sky130_as_sc_hs__dfxtp_2 _52059_ (.CLK(clknet_leaf_89_wb_clk_i),
    .Q(\tholin_riscv.regs[8][16] ),
    .D(_00165_));
 sky130_as_sc_hs__dfxtp_2 _52060_ (.CLK(clknet_leaf_41_wb_clk_i),
    .Q(\tholin_riscv.regs[8][17] ),
    .D(_00166_));
 sky130_as_sc_hs__dfxtp_2 _52061_ (.CLK(clknet_leaf_82_wb_clk_i),
    .Q(\tholin_riscv.regs[8][18] ),
    .D(_00167_));
 sky130_as_sc_hs__dfxtp_2 _52062_ (.CLK(clknet_leaf_46_wb_clk_i),
    .Q(\tholin_riscv.regs[8][19] ),
    .D(_00168_));
 sky130_as_sc_hs__dfxtp_2 _52063_ (.CLK(clknet_leaf_68_wb_clk_i),
    .Q(\tholin_riscv.regs[8][20] ),
    .D(_00169_));
 sky130_as_sc_hs__dfxtp_2 _52064_ (.CLK(clknet_leaf_86_wb_clk_i),
    .Q(\tholin_riscv.regs[8][21] ),
    .D(_00170_));
 sky130_as_sc_hs__dfxtp_2 _52065_ (.CLK(clknet_leaf_71_wb_clk_i),
    .Q(\tholin_riscv.regs[8][22] ),
    .D(_00171_));
 sky130_as_sc_hs__dfxtp_2 _52066_ (.CLK(clknet_leaf_68_wb_clk_i),
    .Q(\tholin_riscv.regs[8][23] ),
    .D(_00172_));
 sky130_as_sc_hs__dfxtp_2 _52067_ (.CLK(clknet_leaf_35_wb_clk_i),
    .Q(\tholin_riscv.regs[8][24] ),
    .D(_00173_));
 sky130_as_sc_hs__dfxtp_2 _52068_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[8][25] ),
    .D(_00174_));
 sky130_as_sc_hs__dfxtp_2 _52069_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[8][26] ),
    .D(_00175_));
 sky130_as_sc_hs__dfxtp_2 _52070_ (.CLK(clknet_leaf_23_wb_clk_i),
    .Q(\tholin_riscv.regs[8][27] ),
    .D(_00176_));
 sky130_as_sc_hs__dfxtp_2 _52071_ (.CLK(clknet_leaf_23_wb_clk_i),
    .Q(\tholin_riscv.regs[8][28] ),
    .D(_00177_));
 sky130_as_sc_hs__dfxtp_2 _52072_ (.CLK(clknet_leaf_36_wb_clk_i),
    .Q(\tholin_riscv.regs[8][29] ),
    .D(_00178_));
 sky130_as_sc_hs__dfxtp_2 _52073_ (.CLK(clknet_leaf_115_wb_clk_i),
    .Q(\tholin_riscv.regs[8][30] ),
    .D(_00179_));
 sky130_as_sc_hs__dfxtp_2 _52074_ (.CLK(clknet_leaf_114_wb_clk_i),
    .Q(\tholin_riscv.regs[8][31] ),
    .D(_00180_));
 sky130_as_sc_hs__dfxtp_2 _52075_ (.CLK(clknet_leaf_131_wb_clk_i),
    .Q(\tholin_riscv.regs[20][0] ),
    .D(net656));
 sky130_as_sc_hs__dfxtp_2 _52076_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.regs[20][1] ),
    .D(_00182_));
 sky130_as_sc_hs__dfxtp_2 _52077_ (.CLK(clknet_leaf_65_wb_clk_i),
    .Q(\tholin_riscv.regs[20][2] ),
    .D(_00183_));
 sky130_as_sc_hs__dfxtp_2 _52078_ (.CLK(clknet_leaf_9_wb_clk_i),
    .Q(\tholin_riscv.regs[20][3] ),
    .D(_00184_));
 sky130_as_sc_hs__dfxtp_2 _52079_ (.CLK(clknet_leaf_67_wb_clk_i),
    .Q(\tholin_riscv.regs[20][4] ),
    .D(_00185_));
 sky130_as_sc_hs__dfxtp_2 _52080_ (.CLK(clknet_leaf_56_wb_clk_i),
    .Q(\tholin_riscv.regs[20][5] ),
    .D(_00186_));
 sky130_as_sc_hs__dfxtp_2 _52081_ (.CLK(clknet_leaf_60_wb_clk_i),
    .Q(\tholin_riscv.regs[20][6] ),
    .D(_00187_));
 sky130_as_sc_hs__dfxtp_2 _52082_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[20][7] ),
    .D(_00188_));
 sky130_as_sc_hs__dfxtp_2 _52083_ (.CLK(clknet_leaf_80_wb_clk_i),
    .Q(\tholin_riscv.regs[20][8] ),
    .D(_00189_));
 sky130_as_sc_hs__dfxtp_2 _52084_ (.CLK(clknet_leaf_42_wb_clk_i),
    .Q(\tholin_riscv.regs[20][9] ),
    .D(_00190_));
 sky130_as_sc_hs__dfxtp_2 _52085_ (.CLK(clknet_leaf_49_wb_clk_i),
    .Q(\tholin_riscv.regs[20][10] ),
    .D(_00191_));
 sky130_as_sc_hs__dfxtp_2 _52086_ (.CLK(clknet_leaf_29_wb_clk_i),
    .Q(\tholin_riscv.regs[20][11] ),
    .D(_00192_));
 sky130_as_sc_hs__dfxtp_2 _52087_ (.CLK(clknet_leaf_27_wb_clk_i),
    .Q(\tholin_riscv.regs[20][12] ),
    .D(_00193_));
 sky130_as_sc_hs__dfxtp_2 _52088_ (.CLK(clknet_leaf_29_wb_clk_i),
    .Q(\tholin_riscv.regs[20][13] ),
    .D(_00194_));
 sky130_as_sc_hs__dfxtp_2 _52089_ (.CLK(clknet_leaf_18_wb_clk_i),
    .Q(\tholin_riscv.regs[20][14] ),
    .D(_00195_));
 sky130_as_sc_hs__dfxtp_2 _52090_ (.CLK(clknet_leaf_16_wb_clk_i),
    .Q(\tholin_riscv.regs[20][15] ),
    .D(_00196_));
 sky130_as_sc_hs__dfxtp_2 _52091_ (.CLK(clknet_leaf_74_wb_clk_i),
    .Q(\tholin_riscv.regs[20][16] ),
    .D(_00197_));
 sky130_as_sc_hs__dfxtp_2 _52092_ (.CLK(clknet_leaf_78_wb_clk_i),
    .Q(\tholin_riscv.regs[20][17] ),
    .D(_00198_));
 sky130_as_sc_hs__dfxtp_2 _52093_ (.CLK(clknet_leaf_123_wb_clk_i),
    .Q(\tholin_riscv.regs[20][18] ),
    .D(_00199_));
 sky130_as_sc_hs__dfxtp_2 _52094_ (.CLK(clknet_leaf_75_wb_clk_i),
    .Q(\tholin_riscv.regs[20][19] ),
    .D(_00200_));
 sky130_as_sc_hs__dfxtp_2 _52095_ (.CLK(clknet_leaf_72_wb_clk_i),
    .Q(\tholin_riscv.regs[20][20] ),
    .D(_00201_));
 sky130_as_sc_hs__dfxtp_2 _52096_ (.CLK(clknet_leaf_80_wb_clk_i),
    .Q(\tholin_riscv.regs[20][21] ),
    .D(_00202_));
 sky130_as_sc_hs__dfxtp_2 _52097_ (.CLK(clknet_leaf_127_wb_clk_i),
    .Q(\tholin_riscv.regs[20][22] ),
    .D(_00203_));
 sky130_as_sc_hs__dfxtp_2 _52098_ (.CLK(clknet_leaf_65_wb_clk_i),
    .Q(\tholin_riscv.regs[20][23] ),
    .D(_00204_));
 sky130_as_sc_hs__dfxtp_2 _52099_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[20][24] ),
    .D(_00205_));
 sky130_as_sc_hs__dfxtp_2 _52100_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[20][25] ),
    .D(_00206_));
 sky130_as_sc_hs__dfxtp_2 _52101_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[20][26] ),
    .D(_00207_));
 sky130_as_sc_hs__dfxtp_2 _52102_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[20][27] ),
    .D(_00208_));
 sky130_as_sc_hs__dfxtp_2 _52103_ (.CLK(clknet_leaf_90_wb_clk_i),
    .Q(\tholin_riscv.regs[20][28] ),
    .D(_00209_));
 sky130_as_sc_hs__dfxtp_2 _52104_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[20][29] ),
    .D(_00210_));
 sky130_as_sc_hs__dfxtp_2 _52105_ (.CLK(clknet_leaf_153_wb_clk_i),
    .Q(\tholin_riscv.regs[20][30] ),
    .D(_00211_));
 sky130_as_sc_hs__dfxtp_2 _52106_ (.CLK(clknet_leaf_102_wb_clk_i),
    .Q(\tholin_riscv.regs[20][31] ),
    .D(_00212_));
 sky130_as_sc_hs__dfxtp_2 _52107_ (.CLK(clknet_leaf_198_wb_clk_i),
    .Q(\tholin_riscv.PC[1] ),
    .D(_00213_));
 sky130_as_sc_hs__dfxtp_2 _52108_ (.CLK(clknet_leaf_65_wb_clk_i),
    .Q(\tholin_riscv.regs[18][0] ),
    .D(net731));
 sky130_as_sc_hs__dfxtp_2 _52109_ (.CLK(clknet_leaf_127_wb_clk_i),
    .Q(\tholin_riscv.regs[18][1] ),
    .D(_00215_));
 sky130_as_sc_hs__dfxtp_2 _52110_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[18][2] ),
    .D(_00216_));
 sky130_as_sc_hs__dfxtp_2 _52111_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[18][3] ),
    .D(_00217_));
 sky130_as_sc_hs__dfxtp_2 _52112_ (.CLK(clknet_leaf_69_wb_clk_i),
    .Q(\tholin_riscv.regs[18][4] ),
    .D(_00218_));
 sky130_as_sc_hs__dfxtp_2 _52113_ (.CLK(clknet_leaf_57_wb_clk_i),
    .Q(\tholin_riscv.regs[18][5] ),
    .D(_00219_));
 sky130_as_sc_hs__dfxtp_2 _52114_ (.CLK(clknet_leaf_56_wb_clk_i),
    .Q(\tholin_riscv.regs[18][6] ),
    .D(_00220_));
 sky130_as_sc_hs__dfxtp_2 _52115_ (.CLK(clknet_leaf_53_wb_clk_i),
    .Q(\tholin_riscv.regs[18][7] ),
    .D(_00221_));
 sky130_as_sc_hs__dfxtp_2 _52116_ (.CLK(clknet_leaf_84_wb_clk_i),
    .Q(\tholin_riscv.regs[18][8] ),
    .D(_00222_));
 sky130_as_sc_hs__dfxtp_2 _52117_ (.CLK(clknet_leaf_38_wb_clk_i),
    .Q(\tholin_riscv.regs[18][9] ),
    .D(_00223_));
 sky130_as_sc_hs__dfxtp_2 _52118_ (.CLK(clknet_leaf_31_wb_clk_i),
    .Q(\tholin_riscv.regs[18][10] ),
    .D(_00224_));
 sky130_as_sc_hs__dfxtp_2 _52119_ (.CLK(clknet_leaf_29_wb_clk_i),
    .Q(\tholin_riscv.regs[18][11] ),
    .D(_00225_));
 sky130_as_sc_hs__dfxtp_2 _52120_ (.CLK(clknet_leaf_27_wb_clk_i),
    .Q(\tholin_riscv.regs[18][12] ),
    .D(_00226_));
 sky130_as_sc_hs__dfxtp_2 _52121_ (.CLK(clknet_leaf_22_wb_clk_i),
    .Q(\tholin_riscv.regs[18][13] ),
    .D(_00227_));
 sky130_as_sc_hs__dfxtp_2 _52122_ (.CLK(clknet_leaf_19_wb_clk_i),
    .Q(\tholin_riscv.regs[18][14] ),
    .D(_00228_));
 sky130_as_sc_hs__dfxtp_2 _52123_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[18][15] ),
    .D(_00229_));
 sky130_as_sc_hs__dfxtp_2 _52124_ (.CLK(clknet_leaf_78_wb_clk_i),
    .Q(\tholin_riscv.regs[18][16] ),
    .D(_00230_));
 sky130_as_sc_hs__dfxtp_2 _52125_ (.CLK(clknet_leaf_78_wb_clk_i),
    .Q(\tholin_riscv.regs[18][17] ),
    .D(_00231_));
 sky130_as_sc_hs__dfxtp_2 _52126_ (.CLK(clknet_leaf_73_wb_clk_i),
    .Q(\tholin_riscv.regs[18][18] ),
    .D(_00232_));
 sky130_as_sc_hs__dfxtp_2 _52127_ (.CLK(clknet_leaf_74_wb_clk_i),
    .Q(\tholin_riscv.regs[18][19] ),
    .D(_00233_));
 sky130_as_sc_hs__dfxtp_2 _52128_ (.CLK(clknet_leaf_73_wb_clk_i),
    .Q(\tholin_riscv.regs[18][20] ),
    .D(_00234_));
 sky130_as_sc_hs__dfxtp_2 _52129_ (.CLK(clknet_leaf_81_wb_clk_i),
    .Q(\tholin_riscv.regs[18][21] ),
    .D(_00235_));
 sky130_as_sc_hs__dfxtp_2 _52130_ (.CLK(clknet_leaf_123_wb_clk_i),
    .Q(\tholin_riscv.regs[18][22] ),
    .D(_00236_));
 sky130_as_sc_hs__dfxtp_2 _52131_ (.CLK(clknet_leaf_66_wb_clk_i),
    .Q(\tholin_riscv.regs[18][23] ),
    .D(_00237_));
 sky130_as_sc_hs__dfxtp_2 _52132_ (.CLK(clknet_leaf_38_wb_clk_i),
    .Q(\tholin_riscv.regs[18][24] ),
    .D(_00238_));
 sky130_as_sc_hs__dfxtp_2 _52133_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[18][25] ),
    .D(_00239_));
 sky130_as_sc_hs__dfxtp_2 _52134_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[18][26] ),
    .D(_00240_));
 sky130_as_sc_hs__dfxtp_2 _52135_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[18][27] ),
    .D(_00241_));
 sky130_as_sc_hs__dfxtp_2 _52136_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[18][28] ),
    .D(_00242_));
 sky130_as_sc_hs__dfxtp_2 _52137_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[18][29] ),
    .D(_00243_));
 sky130_as_sc_hs__dfxtp_2 _52138_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.regs[18][30] ),
    .D(_00244_));
 sky130_as_sc_hs__dfxtp_2 _52139_ (.CLK(clknet_leaf_109_wb_clk_i),
    .Q(\tholin_riscv.regs[18][31] ),
    .D(_00245_));
 sky130_as_sc_hs__dfxtp_2 _52140_ (.CLK(clknet_leaf_65_wb_clk_i),
    .Q(\tholin_riscv.regs[17][0] ),
    .D(net668));
 sky130_as_sc_hs__dfxtp_2 _52141_ (.CLK(clknet_leaf_127_wb_clk_i),
    .Q(\tholin_riscv.regs[17][1] ),
    .D(_00247_));
 sky130_as_sc_hs__dfxtp_2 _52142_ (.CLK(clknet_leaf_8_wb_clk_i),
    .Q(\tholin_riscv.regs[17][2] ),
    .D(_00248_));
 sky130_as_sc_hs__dfxtp_2 _52143_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[17][3] ),
    .D(_00249_));
 sky130_as_sc_hs__dfxtp_2 _52144_ (.CLK(clknet_leaf_147_wb_clk_i),
    .Q(\tholin_riscv.regs[17][4] ),
    .D(_00250_));
 sky130_as_sc_hs__dfxtp_2 _52145_ (.CLK(clknet_leaf_57_wb_clk_i),
    .Q(\tholin_riscv.regs[17][5] ),
    .D(_00251_));
 sky130_as_sc_hs__dfxtp_2 _52146_ (.CLK(clknet_leaf_62_wb_clk_i),
    .Q(\tholin_riscv.regs[17][6] ),
    .D(_00252_));
 sky130_as_sc_hs__dfxtp_2 _52147_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[17][7] ),
    .D(_00253_));
 sky130_as_sc_hs__dfxtp_2 _52148_ (.CLK(clknet_leaf_84_wb_clk_i),
    .Q(\tholin_riscv.regs[17][8] ),
    .D(_00254_));
 sky130_as_sc_hs__dfxtp_2 _52149_ (.CLK(clknet_leaf_42_wb_clk_i),
    .Q(\tholin_riscv.regs[17][9] ),
    .D(_00255_));
 sky130_as_sc_hs__dfxtp_2 _52150_ (.CLK(clknet_leaf_31_wb_clk_i),
    .Q(\tholin_riscv.regs[17][10] ),
    .D(_00256_));
 sky130_as_sc_hs__dfxtp_2 _52151_ (.CLK(clknet_leaf_29_wb_clk_i),
    .Q(\tholin_riscv.regs[17][11] ),
    .D(_00257_));
 sky130_as_sc_hs__dfxtp_2 _52152_ (.CLK(clknet_leaf_27_wb_clk_i),
    .Q(\tholin_riscv.regs[17][12] ),
    .D(_00258_));
 sky130_as_sc_hs__dfxtp_2 _52153_ (.CLK(clknet_leaf_22_wb_clk_i),
    .Q(\tholin_riscv.regs[17][13] ),
    .D(_00259_));
 sky130_as_sc_hs__dfxtp_2 _52154_ (.CLK(clknet_leaf_19_wb_clk_i),
    .Q(\tholin_riscv.regs[17][14] ),
    .D(_00260_));
 sky130_as_sc_hs__dfxtp_2 _52155_ (.CLK(clknet_leaf_16_wb_clk_i),
    .Q(\tholin_riscv.regs[17][15] ),
    .D(_00261_));
 sky130_as_sc_hs__dfxtp_2 _52156_ (.CLK(clknet_leaf_104_wb_clk_i),
    .Q(\tholin_riscv.regs[17][16] ),
    .D(_00262_));
 sky130_as_sc_hs__dfxtp_2 _52157_ (.CLK(clknet_leaf_106_wb_clk_i),
    .Q(\tholin_riscv.regs[17][17] ),
    .D(_00263_));
 sky130_as_sc_hs__dfxtp_2 _52158_ (.CLK(clknet_leaf_115_wb_clk_i),
    .Q(\tholin_riscv.regs[17][18] ),
    .D(_00264_));
 sky130_as_sc_hs__dfxtp_2 _52159_ (.CLK(clknet_leaf_118_wb_clk_i),
    .Q(\tholin_riscv.regs[17][19] ),
    .D(_00265_));
 sky130_as_sc_hs__dfxtp_2 _52160_ (.CLK(clknet_leaf_118_wb_clk_i),
    .Q(\tholin_riscv.regs[17][20] ),
    .D(_00266_));
 sky130_as_sc_hs__dfxtp_2 _52161_ (.CLK(clknet_leaf_115_wb_clk_i),
    .Q(\tholin_riscv.regs[17][21] ),
    .D(_00267_));
 sky130_as_sc_hs__dfxtp_2 _52162_ (.CLK(clknet_leaf_149_wb_clk_i),
    .Q(\tholin_riscv.regs[17][22] ),
    .D(_00268_));
 sky130_as_sc_hs__dfxtp_2 _52163_ (.CLK(clknet_leaf_115_wb_clk_i),
    .Q(\tholin_riscv.regs[17][23] ),
    .D(_00269_));
 sky130_as_sc_hs__dfxtp_2 _52164_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[17][24] ),
    .D(_00270_));
 sky130_as_sc_hs__dfxtp_2 _52165_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[17][25] ),
    .D(_00271_));
 sky130_as_sc_hs__dfxtp_2 _52166_ (.CLK(clknet_leaf_89_wb_clk_i),
    .Q(\tholin_riscv.regs[17][26] ),
    .D(_00272_));
 sky130_as_sc_hs__dfxtp_2 _52167_ (.CLK(clknet_leaf_90_wb_clk_i),
    .Q(\tholin_riscv.regs[17][27] ),
    .D(_00273_));
 sky130_as_sc_hs__dfxtp_2 _52168_ (.CLK(clknet_leaf_89_wb_clk_i),
    .Q(\tholin_riscv.regs[17][28] ),
    .D(_00274_));
 sky130_as_sc_hs__dfxtp_2 _52169_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[17][29] ),
    .D(_00275_));
 sky130_as_sc_hs__dfxtp_2 _52170_ (.CLK(clknet_leaf_94_wb_clk_i),
    .Q(\tholin_riscv.regs[17][30] ),
    .D(_00276_));
 sky130_as_sc_hs__dfxtp_2 _52171_ (.CLK(clknet_leaf_150_wb_clk_i),
    .Q(\tholin_riscv.regs[17][31] ),
    .D(_00277_));
 sky130_as_sc_hs__dfxtp_2 _52172_ (.CLK(clknet_leaf_133_wb_clk_i),
    .Q(\tholin_riscv.regs[15][0] ),
    .D(net689));
 sky130_as_sc_hs__dfxtp_2 _52173_ (.CLK(clknet_leaf_129_wb_clk_i),
    .Q(\tholin_riscv.regs[15][1] ),
    .D(_00279_));
 sky130_as_sc_hs__dfxtp_2 _52174_ (.CLK(clknet_leaf_64_wb_clk_i),
    .Q(\tholin_riscv.regs[15][2] ),
    .D(_00280_));
 sky130_as_sc_hs__dfxtp_2 _52175_ (.CLK(clknet_leaf_56_wb_clk_i),
    .Q(\tholin_riscv.regs[15][3] ),
    .D(_00281_));
 sky130_as_sc_hs__dfxtp_2 _52176_ (.CLK(clknet_leaf_103_wb_clk_i),
    .Q(\tholin_riscv.regs[15][4] ),
    .D(_00282_));
 sky130_as_sc_hs__dfxtp_2 _52177_ (.CLK(clknet_leaf_47_wb_clk_i),
    .Q(\tholin_riscv.regs[15][5] ),
    .D(_00283_));
 sky130_as_sc_hs__dfxtp_2 _52178_ (.CLK(clknet_leaf_61_wb_clk_i),
    .Q(\tholin_riscv.regs[15][6] ),
    .D(_00284_));
 sky130_as_sc_hs__dfxtp_2 _52179_ (.CLK(clknet_leaf_47_wb_clk_i),
    .Q(\tholin_riscv.regs[15][7] ),
    .D(_00285_));
 sky130_as_sc_hs__dfxtp_2 _52180_ (.CLK(clknet_leaf_84_wb_clk_i),
    .Q(\tholin_riscv.regs[15][8] ),
    .D(_00286_));
 sky130_as_sc_hs__dfxtp_2 _52181_ (.CLK(clknet_leaf_45_wb_clk_i),
    .Q(\tholin_riscv.regs[15][9] ),
    .D(_00287_));
 sky130_as_sc_hs__dfxtp_2 _52182_ (.CLK(clknet_leaf_48_wb_clk_i),
    .Q(\tholin_riscv.regs[15][10] ),
    .D(_00288_));
 sky130_as_sc_hs__dfxtp_2 _52183_ (.CLK(clknet_leaf_49_wb_clk_i),
    .Q(\tholin_riscv.regs[15][11] ),
    .D(_00289_));
 sky130_as_sc_hs__dfxtp_2 _52184_ (.CLK(clknet_leaf_32_wb_clk_i),
    .Q(\tholin_riscv.regs[15][12] ),
    .D(_00290_));
 sky130_as_sc_hs__dfxtp_2 _52185_ (.CLK(clknet_leaf_25_wb_clk_i),
    .Q(\tholin_riscv.regs[15][13] ),
    .D(_00291_));
 sky130_as_sc_hs__dfxtp_2 _52186_ (.CLK(clknet_leaf_14_wb_clk_i),
    .Q(\tholin_riscv.regs[15][14] ),
    .D(_00292_));
 sky130_as_sc_hs__dfxtp_2 _52187_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[15][15] ),
    .D(_00293_));
 sky130_as_sc_hs__dfxtp_2 _52188_ (.CLK(clknet_leaf_119_wb_clk_i),
    .Q(\tholin_riscv.regs[15][16] ),
    .D(_00294_));
 sky130_as_sc_hs__dfxtp_2 _52189_ (.CLK(clknet_leaf_109_wb_clk_i),
    .Q(\tholin_riscv.regs[15][17] ),
    .D(_00295_));
 sky130_as_sc_hs__dfxtp_2 _52190_ (.CLK(clknet_leaf_113_wb_clk_i),
    .Q(\tholin_riscv.regs[15][18] ),
    .D(_00296_));
 sky130_as_sc_hs__dfxtp_2 _52191_ (.CLK(clknet_leaf_107_wb_clk_i),
    .Q(\tholin_riscv.regs[15][19] ),
    .D(_00297_));
 sky130_as_sc_hs__dfxtp_2 _52192_ (.CLK(clknet_leaf_149_wb_clk_i),
    .Q(\tholin_riscv.regs[15][20] ),
    .D(_00298_));
 sky130_as_sc_hs__dfxtp_2 _52193_ (.CLK(clknet_leaf_145_wb_clk_i),
    .Q(\tholin_riscv.regs[15][21] ),
    .D(_00299_));
 sky130_as_sc_hs__dfxtp_2 _52194_ (.CLK(clknet_leaf_149_wb_clk_i),
    .Q(\tholin_riscv.regs[15][22] ),
    .D(_00300_));
 sky130_as_sc_hs__dfxtp_2 _52195_ (.CLK(clknet_leaf_103_wb_clk_i),
    .Q(\tholin_riscv.regs[15][23] ),
    .D(_00301_));
 sky130_as_sc_hs__dfxtp_2 _52196_ (.CLK(clknet_leaf_35_wb_clk_i),
    .Q(\tholin_riscv.regs[15][24] ),
    .D(_00302_));
 sky130_as_sc_hs__dfxtp_2 _52197_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[15][25] ),
    .D(_00303_));
 sky130_as_sc_hs__dfxtp_2 _52198_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[15][26] ),
    .D(_00304_));
 sky130_as_sc_hs__dfxtp_2 _52199_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[15][27] ),
    .D(_00305_));
 sky130_as_sc_hs__dfxtp_2 _52200_ (.CLK(clknet_leaf_23_wb_clk_i),
    .Q(\tholin_riscv.regs[15][28] ),
    .D(_00306_));
 sky130_as_sc_hs__dfxtp_2 _52201_ (.CLK(clknet_leaf_38_wb_clk_i),
    .Q(\tholin_riscv.regs[15][29] ),
    .D(_00307_));
 sky130_as_sc_hs__dfxtp_2 _52202_ (.CLK(clknet_leaf_120_wb_clk_i),
    .Q(\tholin_riscv.regs[15][30] ),
    .D(_00308_));
 sky130_as_sc_hs__dfxtp_2 _52203_ (.CLK(clknet_leaf_158_wb_clk_i),
    .Q(\tholin_riscv.regs[15][31] ),
    .D(_00309_));
 sky130_as_sc_hs__dfxtp_2 _52204_ (.CLK(clknet_leaf_132_wb_clk_i),
    .Q(\tholin_riscv.regs[13][0] ),
    .D(net653));
 sky130_as_sc_hs__dfxtp_2 _52205_ (.CLK(clknet_leaf_128_wb_clk_i),
    .Q(\tholin_riscv.regs[13][1] ),
    .D(_00311_));
 sky130_as_sc_hs__dfxtp_2 _52206_ (.CLK(clknet_leaf_64_wb_clk_i),
    .Q(\tholin_riscv.regs[13][2] ),
    .D(_00312_));
 sky130_as_sc_hs__dfxtp_2 _52207_ (.CLK(clknet_leaf_56_wb_clk_i),
    .Q(\tholin_riscv.regs[13][3] ),
    .D(_00313_));
 sky130_as_sc_hs__dfxtp_2 _52208_ (.CLK(clknet_leaf_101_wb_clk_i),
    .Q(\tholin_riscv.regs[13][4] ),
    .D(_00314_));
 sky130_as_sc_hs__dfxtp_2 _52209_ (.CLK(clknet_leaf_47_wb_clk_i),
    .Q(\tholin_riscv.regs[13][5] ),
    .D(_00315_));
 sky130_as_sc_hs__dfxtp_2 _52210_ (.CLK(clknet_leaf_61_wb_clk_i),
    .Q(\tholin_riscv.regs[13][6] ),
    .D(_00316_));
 sky130_as_sc_hs__dfxtp_2 _52211_ (.CLK(clknet_leaf_50_wb_clk_i),
    .Q(\tholin_riscv.regs[13][7] ),
    .D(_00317_));
 sky130_as_sc_hs__dfxtp_2 _52212_ (.CLK(clknet_leaf_82_wb_clk_i),
    .Q(\tholin_riscv.regs[13][8] ),
    .D(_00318_));
 sky130_as_sc_hs__dfxtp_2 _52213_ (.CLK(clknet_leaf_83_wb_clk_i),
    .Q(\tholin_riscv.regs[13][9] ),
    .D(_00319_));
 sky130_as_sc_hs__dfxtp_2 _52214_ (.CLK(clknet_leaf_48_wb_clk_i),
    .Q(\tholin_riscv.regs[13][10] ),
    .D(_00320_));
 sky130_as_sc_hs__dfxtp_2 _52215_ (.CLK(clknet_leaf_50_wb_clk_i),
    .Q(\tholin_riscv.regs[13][11] ),
    .D(_00321_));
 sky130_as_sc_hs__dfxtp_2 _52216_ (.CLK(clknet_leaf_32_wb_clk_i),
    .Q(\tholin_riscv.regs[13][12] ),
    .D(_00322_));
 sky130_as_sc_hs__dfxtp_2 _52217_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[13][13] ),
    .D(_00323_));
 sky130_as_sc_hs__dfxtp_2 _52218_ (.CLK(clknet_leaf_15_wb_clk_i),
    .Q(\tholin_riscv.regs[13][14] ),
    .D(_00324_));
 sky130_as_sc_hs__dfxtp_2 _52219_ (.CLK(clknet_leaf_16_wb_clk_i),
    .Q(\tholin_riscv.regs[13][15] ),
    .D(_00325_));
 sky130_as_sc_hs__dfxtp_2 _52220_ (.CLK(clknet_leaf_115_wb_clk_i),
    .Q(\tholin_riscv.regs[13][16] ),
    .D(_00326_));
 sky130_as_sc_hs__dfxtp_2 _52221_ (.CLK(clknet_leaf_147_wb_clk_i),
    .Q(\tholin_riscv.regs[13][17] ),
    .D(_00327_));
 sky130_as_sc_hs__dfxtp_2 _52222_ (.CLK(clknet_leaf_150_wb_clk_i),
    .Q(\tholin_riscv.regs[13][18] ),
    .D(_00328_));
 sky130_as_sc_hs__dfxtp_2 _52223_ (.CLK(clknet_leaf_105_wb_clk_i),
    .Q(\tholin_riscv.regs[13][19] ),
    .D(_00329_));
 sky130_as_sc_hs__dfxtp_2 _52224_ (.CLK(clknet_leaf_108_wb_clk_i),
    .Q(\tholin_riscv.regs[13][20] ),
    .D(_00330_));
 sky130_as_sc_hs__dfxtp_2 _52225_ (.CLK(clknet_leaf_102_wb_clk_i),
    .Q(\tholin_riscv.regs[13][21] ),
    .D(_00331_));
 sky130_as_sc_hs__dfxtp_2 _52226_ (.CLK(clknet_leaf_142_wb_clk_i),
    .Q(\tholin_riscv.regs[13][22] ),
    .D(_00332_));
 sky130_as_sc_hs__dfxtp_2 _52227_ (.CLK(clknet_leaf_147_wb_clk_i),
    .Q(\tholin_riscv.regs[13][23] ),
    .D(_00333_));
 sky130_as_sc_hs__dfxtp_2 _52228_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[13][24] ),
    .D(_00334_));
 sky130_as_sc_hs__dfxtp_2 _52229_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[13][25] ),
    .D(_00335_));
 sky130_as_sc_hs__dfxtp_2 _52230_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[13][26] ),
    .D(_00336_));
 sky130_as_sc_hs__dfxtp_2 _52231_ (.CLK(clknet_leaf_23_wb_clk_i),
    .Q(\tholin_riscv.regs[13][27] ),
    .D(_00337_));
 sky130_as_sc_hs__dfxtp_2 _52232_ (.CLK(clknet_leaf_23_wb_clk_i),
    .Q(\tholin_riscv.regs[13][28] ),
    .D(_00338_));
 sky130_as_sc_hs__dfxtp_2 _52233_ (.CLK(clknet_leaf_38_wb_clk_i),
    .Q(\tholin_riscv.regs[13][29] ),
    .D(_00339_));
 sky130_as_sc_hs__dfxtp_2 _52234_ (.CLK(clknet_leaf_115_wb_clk_i),
    .Q(\tholin_riscv.regs[13][30] ),
    .D(_00340_));
 sky130_as_sc_hs__dfxtp_2 _52235_ (.CLK(clknet_leaf_158_wb_clk_i),
    .Q(\tholin_riscv.regs[13][31] ),
    .D(_00341_));
 sky130_as_sc_hs__dfxtp_2 _52236_ (.CLK(clknet_leaf_132_wb_clk_i),
    .Q(\tholin_riscv.regs[12][0] ),
    .D(net698));
 sky130_as_sc_hs__dfxtp_2 _52237_ (.CLK(clknet_leaf_128_wb_clk_i),
    .Q(\tholin_riscv.regs[12][1] ),
    .D(_00343_));
 sky130_as_sc_hs__dfxtp_2 _52238_ (.CLK(clknet_leaf_64_wb_clk_i),
    .Q(\tholin_riscv.regs[12][2] ),
    .D(_00344_));
 sky130_as_sc_hs__dfxtp_2 _52239_ (.CLK(clknet_leaf_56_wb_clk_i),
    .Q(\tholin_riscv.regs[12][3] ),
    .D(_00345_));
 sky130_as_sc_hs__dfxtp_2 _52240_ (.CLK(clknet_leaf_70_wb_clk_i),
    .Q(\tholin_riscv.regs[12][4] ),
    .D(_00346_));
 sky130_as_sc_hs__dfxtp_2 _52241_ (.CLK(clknet_leaf_47_wb_clk_i),
    .Q(\tholin_riscv.regs[12][5] ),
    .D(_00347_));
 sky130_as_sc_hs__dfxtp_2 _52242_ (.CLK(clknet_leaf_61_wb_clk_i),
    .Q(\tholin_riscv.regs[12][6] ),
    .D(_00348_));
 sky130_as_sc_hs__dfxtp_2 _52243_ (.CLK(clknet_leaf_47_wb_clk_i),
    .Q(\tholin_riscv.regs[12][7] ),
    .D(_00349_));
 sky130_as_sc_hs__dfxtp_2 _52244_ (.CLK(clknet_leaf_84_wb_clk_i),
    .Q(\tholin_riscv.regs[12][8] ),
    .D(_00350_));
 sky130_as_sc_hs__dfxtp_2 _52245_ (.CLK(clknet_leaf_45_wb_clk_i),
    .Q(\tholin_riscv.regs[12][9] ),
    .D(_00351_));
 sky130_as_sc_hs__dfxtp_2 _52246_ (.CLK(clknet_leaf_48_wb_clk_i),
    .Q(\tholin_riscv.regs[12][10] ),
    .D(_00352_));
 sky130_as_sc_hs__dfxtp_2 _52247_ (.CLK(clknet_leaf_50_wb_clk_i),
    .Q(\tholin_riscv.regs[12][11] ),
    .D(_00353_));
 sky130_as_sc_hs__dfxtp_2 _52248_ (.CLK(clknet_leaf_32_wb_clk_i),
    .Q(\tholin_riscv.regs[12][12] ),
    .D(_00354_));
 sky130_as_sc_hs__dfxtp_2 _52249_ (.CLK(clknet_leaf_28_wb_clk_i),
    .Q(\tholin_riscv.regs[12][13] ),
    .D(_00355_));
 sky130_as_sc_hs__dfxtp_2 _52250_ (.CLK(clknet_leaf_14_wb_clk_i),
    .Q(\tholin_riscv.regs[12][14] ),
    .D(_00356_));
 sky130_as_sc_hs__dfxtp_2 _52251_ (.CLK(clknet_leaf_16_wb_clk_i),
    .Q(\tholin_riscv.regs[12][15] ),
    .D(_00357_));
 sky130_as_sc_hs__dfxtp_2 _52252_ (.CLK(clknet_leaf_89_wb_clk_i),
    .Q(\tholin_riscv.regs[12][16] ),
    .D(_00358_));
 sky130_as_sc_hs__dfxtp_2 _52253_ (.CLK(clknet_leaf_41_wb_clk_i),
    .Q(\tholin_riscv.regs[12][17] ),
    .D(_00359_));
 sky130_as_sc_hs__dfxtp_2 _52254_ (.CLK(clknet_leaf_82_wb_clk_i),
    .Q(\tholin_riscv.regs[12][18] ),
    .D(_00360_));
 sky130_as_sc_hs__dfxtp_2 _52255_ (.CLK(clknet_leaf_46_wb_clk_i),
    .Q(\tholin_riscv.regs[12][19] ),
    .D(_00361_));
 sky130_as_sc_hs__dfxtp_2 _52256_ (.CLK(clknet_leaf_73_wb_clk_i),
    .Q(\tholin_riscv.regs[12][20] ),
    .D(_00362_));
 sky130_as_sc_hs__dfxtp_2 _52257_ (.CLK(clknet_leaf_86_wb_clk_i),
    .Q(\tholin_riscv.regs[12][21] ),
    .D(_00363_));
 sky130_as_sc_hs__dfxtp_2 _52258_ (.CLK(clknet_leaf_71_wb_clk_i),
    .Q(\tholin_riscv.regs[12][22] ),
    .D(_00364_));
 sky130_as_sc_hs__dfxtp_2 _52259_ (.CLK(clknet_leaf_68_wb_clk_i),
    .Q(\tholin_riscv.regs[12][23] ),
    .D(_00365_));
 sky130_as_sc_hs__dfxtp_2 _52260_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[12][24] ),
    .D(_00366_));
 sky130_as_sc_hs__dfxtp_2 _52261_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[12][25] ),
    .D(_00367_));
 sky130_as_sc_hs__dfxtp_2 _52262_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[12][26] ),
    .D(_00368_));
 sky130_as_sc_hs__dfxtp_2 _52263_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[12][27] ),
    .D(_00369_));
 sky130_as_sc_hs__dfxtp_2 _52264_ (.CLK(clknet_leaf_23_wb_clk_i),
    .Q(\tholin_riscv.regs[12][28] ),
    .D(_00370_));
 sky130_as_sc_hs__dfxtp_2 _52265_ (.CLK(clknet_leaf_38_wb_clk_i),
    .Q(\tholin_riscv.regs[12][29] ),
    .D(_00371_));
 sky130_as_sc_hs__dfxtp_2 _52266_ (.CLK(clknet_leaf_112_wb_clk_i),
    .Q(\tholin_riscv.regs[12][30] ),
    .D(_00372_));
 sky130_as_sc_hs__dfxtp_2 _52267_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.regs[12][31] ),
    .D(_00373_));
 sky130_as_sc_hs__dfxtp_2 _52268_ (.CLK(clknet_leaf_130_wb_clk_i),
    .Q(\tholin_riscv.regs[10][0] ),
    .D(net707));
 sky130_as_sc_hs__dfxtp_2 _52269_ (.CLK(clknet_leaf_128_wb_clk_i),
    .Q(\tholin_riscv.regs[10][1] ),
    .D(_00375_));
 sky130_as_sc_hs__dfxtp_2 _52270_ (.CLK(clknet_leaf_66_wb_clk_i),
    .Q(\tholin_riscv.regs[10][2] ),
    .D(_00376_));
 sky130_as_sc_hs__dfxtp_2 _52271_ (.CLK(clknet_leaf_55_wb_clk_i),
    .Q(\tholin_riscv.regs[10][3] ),
    .D(_00377_));
 sky130_as_sc_hs__dfxtp_2 _52272_ (.CLK(clknet_leaf_69_wb_clk_i),
    .Q(\tholin_riscv.regs[10][4] ),
    .D(_00378_));
 sky130_as_sc_hs__dfxtp_2 _52273_ (.CLK(clknet_leaf_59_wb_clk_i),
    .Q(\tholin_riscv.regs[10][5] ),
    .D(_00379_));
 sky130_as_sc_hs__dfxtp_2 _52274_ (.CLK(clknet_leaf_64_wb_clk_i),
    .Q(\tholin_riscv.regs[10][6] ),
    .D(_00380_));
 sky130_as_sc_hs__dfxtp_2 _52275_ (.CLK(clknet_leaf_58_wb_clk_i),
    .Q(\tholin_riscv.regs[10][7] ),
    .D(_00381_));
 sky130_as_sc_hs__dfxtp_2 _52276_ (.CLK(clknet_leaf_83_wb_clk_i),
    .Q(\tholin_riscv.regs[10][8] ),
    .D(_00382_));
 sky130_as_sc_hs__dfxtp_2 _52277_ (.CLK(clknet_leaf_44_wb_clk_i),
    .Q(\tholin_riscv.regs[10][9] ),
    .D(_00383_));
 sky130_as_sc_hs__dfxtp_2 _52278_ (.CLK(clknet_leaf_49_wb_clk_i),
    .Q(\tholin_riscv.regs[10][10] ),
    .D(_00384_));
 sky130_as_sc_hs__dfxtp_2 _52279_ (.CLK(clknet_leaf_31_wb_clk_i),
    .Q(\tholin_riscv.regs[10][11] ),
    .D(_00385_));
 sky130_as_sc_hs__dfxtp_2 _52280_ (.CLK(clknet_leaf_31_wb_clk_i),
    .Q(\tholin_riscv.regs[10][12] ),
    .D(_00386_));
 sky130_as_sc_hs__dfxtp_2 _52281_ (.CLK(clknet_leaf_27_wb_clk_i),
    .Q(\tholin_riscv.regs[10][13] ),
    .D(_00387_));
 sky130_as_sc_hs__dfxtp_2 _52282_ (.CLK(clknet_leaf_14_wb_clk_i),
    .Q(\tholin_riscv.regs[10][14] ),
    .D(_00388_));
 sky130_as_sc_hs__dfxtp_2 _52283_ (.CLK(clknet_leaf_15_wb_clk_i),
    .Q(\tholin_riscv.regs[10][15] ),
    .D(_00389_));
 sky130_as_sc_hs__dfxtp_2 _52284_ (.CLK(clknet_leaf_89_wb_clk_i),
    .Q(\tholin_riscv.regs[10][16] ),
    .D(_00390_));
 sky130_as_sc_hs__dfxtp_2 _52285_ (.CLK(clknet_leaf_41_wb_clk_i),
    .Q(\tholin_riscv.regs[10][17] ),
    .D(_00391_));
 sky130_as_sc_hs__dfxtp_2 _52286_ (.CLK(clknet_leaf_82_wb_clk_i),
    .Q(\tholin_riscv.regs[10][18] ),
    .D(_00392_));
 sky130_as_sc_hs__dfxtp_2 _52287_ (.CLK(clknet_leaf_46_wb_clk_i),
    .Q(\tholin_riscv.regs[10][19] ),
    .D(_00393_));
 sky130_as_sc_hs__dfxtp_2 _52288_ (.CLK(clknet_leaf_68_wb_clk_i),
    .Q(\tholin_riscv.regs[10][20] ),
    .D(_00394_));
 sky130_as_sc_hs__dfxtp_2 _52289_ (.CLK(clknet_leaf_86_wb_clk_i),
    .Q(\tholin_riscv.regs[10][21] ),
    .D(_00395_));
 sky130_as_sc_hs__dfxtp_2 _52290_ (.CLK(clknet_leaf_71_wb_clk_i),
    .Q(\tholin_riscv.regs[10][22] ),
    .D(_00396_));
 sky130_as_sc_hs__dfxtp_2 _52291_ (.CLK(clknet_leaf_69_wb_clk_i),
    .Q(\tholin_riscv.regs[10][23] ),
    .D(_00397_));
 sky130_as_sc_hs__dfxtp_2 _52292_ (.CLK(clknet_leaf_33_wb_clk_i),
    .Q(\tholin_riscv.regs[10][24] ),
    .D(_00398_));
 sky130_as_sc_hs__dfxtp_2 _52293_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[10][25] ),
    .D(_00399_));
 sky130_as_sc_hs__dfxtp_2 _52294_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[10][26] ),
    .D(_00400_));
 sky130_as_sc_hs__dfxtp_2 _52295_ (.CLK(clknet_leaf_25_wb_clk_i),
    .Q(\tholin_riscv.regs[10][27] ),
    .D(_00401_));
 sky130_as_sc_hs__dfxtp_2 _52296_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[10][28] ),
    .D(_00402_));
 sky130_as_sc_hs__dfxtp_2 _52297_ (.CLK(clknet_leaf_39_wb_clk_i),
    .Q(\tholin_riscv.regs[10][29] ),
    .D(_00403_));
 sky130_as_sc_hs__dfxtp_2 _52298_ (.CLK(clknet_leaf_117_wb_clk_i),
    .Q(\tholin_riscv.regs[10][30] ),
    .D(_00404_));
 sky130_as_sc_hs__dfxtp_2 _52299_ (.CLK(clknet_leaf_157_wb_clk_i),
    .Q(\tholin_riscv.regs[10][31] ),
    .D(_00405_));
 sky130_as_sc_hs__dfxtp_2 _52300_ (.CLK(clknet_leaf_130_wb_clk_i),
    .Q(\tholin_riscv.regs[0][0] ),
    .D(_00406_));
 sky130_as_sc_hs__dfxtp_2 _52301_ (.CLK(clknet_leaf_129_wb_clk_i),
    .Q(\tholin_riscv.regs[0][1] ),
    .D(_00407_));
 sky130_as_sc_hs__dfxtp_2 _52302_ (.CLK(clknet_leaf_66_wb_clk_i),
    .Q(\tholin_riscv.regs[0][2] ),
    .D(_00408_));
 sky130_as_sc_hs__dfxtp_2 _52303_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[0][3] ),
    .D(_00409_));
 sky130_as_sc_hs__dfxtp_2 _52304_ (.CLK(clknet_leaf_60_wb_clk_i),
    .Q(\tholin_riscv.regs[0][4] ),
    .D(_00410_));
 sky130_as_sc_hs__dfxtp_2 _52305_ (.CLK(clknet_leaf_58_wb_clk_i),
    .Q(\tholin_riscv.regs[0][5] ),
    .D(_00411_));
 sky130_as_sc_hs__dfxtp_2 _52306_ (.CLK(clknet_leaf_60_wb_clk_i),
    .Q(\tholin_riscv.regs[0][6] ),
    .D(_00412_));
 sky130_as_sc_hs__dfxtp_2 _52307_ (.CLK(clknet_leaf_51_wb_clk_i),
    .Q(\tholin_riscv.regs[0][7] ),
    .D(_00413_));
 sky130_as_sc_hs__dfxtp_2 _52308_ (.CLK(clknet_leaf_83_wb_clk_i),
    .Q(\tholin_riscv.regs[0][8] ),
    .D(_00414_));
 sky130_as_sc_hs__dfxtp_2 _52309_ (.CLK(clknet_leaf_45_wb_clk_i),
    .Q(\tholin_riscv.regs[0][9] ),
    .D(_00415_));
 sky130_as_sc_hs__dfxtp_2 _52310_ (.CLK(clknet_leaf_48_wb_clk_i),
    .Q(\tholin_riscv.regs[0][10] ),
    .D(_00416_));
 sky130_as_sc_hs__dfxtp_2 _52311_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[0][11] ),
    .D(_00417_));
 sky130_as_sc_hs__dfxtp_2 _52312_ (.CLK(clknet_leaf_37_wb_clk_i),
    .Q(\tholin_riscv.regs[0][12] ),
    .D(_00418_));
 sky130_as_sc_hs__dfxtp_2 _52313_ (.CLK(clknet_leaf_33_wb_clk_i),
    .Q(\tholin_riscv.regs[0][13] ),
    .D(_00419_));
 sky130_as_sc_hs__dfxtp_2 _52314_ (.CLK(clknet_leaf_12_wb_clk_i),
    .Q(\tholin_riscv.regs[0][14] ),
    .D(_00420_));
 sky130_as_sc_hs__dfxtp_2 _52315_ (.CLK(clknet_leaf_14_wb_clk_i),
    .Q(\tholin_riscv.regs[0][15] ),
    .D(_00421_));
 sky130_as_sc_hs__dfxtp_2 _52316_ (.CLK(clknet_leaf_85_wb_clk_i),
    .Q(\tholin_riscv.regs[0][16] ),
    .D(_00422_));
 sky130_as_sc_hs__dfxtp_2 _52317_ (.CLK(clknet_leaf_41_wb_clk_i),
    .Q(\tholin_riscv.regs[0][17] ),
    .D(_00423_));
 sky130_as_sc_hs__dfxtp_2 _52318_ (.CLK(clknet_leaf_83_wb_clk_i),
    .Q(\tholin_riscv.regs[0][18] ),
    .D(_00424_));
 sky130_as_sc_hs__dfxtp_2 _52319_ (.CLK(clknet_leaf_46_wb_clk_i),
    .Q(\tholin_riscv.regs[0][19] ),
    .D(_00425_));
 sky130_as_sc_hs__dfxtp_2 _52320_ (.CLK(clknet_leaf_69_wb_clk_i),
    .Q(\tholin_riscv.regs[0][20] ),
    .D(_00426_));
 sky130_as_sc_hs__dfxtp_2 _52321_ (.CLK(clknet_leaf_86_wb_clk_i),
    .Q(\tholin_riscv.regs[0][21] ),
    .D(_00427_));
 sky130_as_sc_hs__dfxtp_2 _52322_ (.CLK(clknet_leaf_82_wb_clk_i),
    .Q(\tholin_riscv.regs[0][22] ),
    .D(_00428_));
 sky130_as_sc_hs__dfxtp_2 _52323_ (.CLK(clknet_leaf_67_wb_clk_i),
    .Q(\tholin_riscv.regs[0][23] ),
    .D(_00429_));
 sky130_as_sc_hs__dfxtp_2 _52324_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[0][24] ),
    .D(_00430_));
 sky130_as_sc_hs__dfxtp_2 _52325_ (.CLK(clknet_leaf_16_wb_clk_i),
    .Q(\tholin_riscv.regs[0][25] ),
    .D(_00431_));
 sky130_as_sc_hs__dfxtp_2 _52326_ (.CLK(clknet_leaf_25_wb_clk_i),
    .Q(\tholin_riscv.regs[0][26] ),
    .D(_00432_));
 sky130_as_sc_hs__dfxtp_2 _52327_ (.CLK(clknet_leaf_25_wb_clk_i),
    .Q(\tholin_riscv.regs[0][27] ),
    .D(_00433_));
 sky130_as_sc_hs__dfxtp_2 _52328_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[0][28] ),
    .D(_00434_));
 sky130_as_sc_hs__dfxtp_2 _52329_ (.CLK(clknet_leaf_36_wb_clk_i),
    .Q(\tholin_riscv.regs[0][29] ),
    .D(_00435_));
 sky130_as_sc_hs__dfxtp_2 _52330_ (.CLK(clknet_leaf_72_wb_clk_i),
    .Q(\tholin_riscv.regs[0][30] ),
    .D(_00436_));
 sky130_as_sc_hs__dfxtp_2 _52331_ (.CLK(clknet_leaf_72_wb_clk_i),
    .Q(\tholin_riscv.regs[0][31] ),
    .D(_00437_));
 sky130_as_sc_hs__dfxtp_2 _52332_ (.CLK(clknet_leaf_133_wb_clk_i),
    .Q(\tholin_riscv.regs[7][0] ),
    .D(net683));
 sky130_as_sc_hs__dfxtp_2 _52333_ (.CLK(clknet_leaf_68_wb_clk_i),
    .Q(\tholin_riscv.regs[7][1] ),
    .D(_00439_));
 sky130_as_sc_hs__dfxtp_2 _52334_ (.CLK(clknet_leaf_65_wb_clk_i),
    .Q(\tholin_riscv.regs[7][2] ),
    .D(_00440_));
 sky130_as_sc_hs__dfxtp_2 _52335_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[7][3] ),
    .D(_00441_));
 sky130_as_sc_hs__dfxtp_2 _52336_ (.CLK(clknet_leaf_115_wb_clk_i),
    .Q(\tholin_riscv.regs[7][4] ),
    .D(_00442_));
 sky130_as_sc_hs__dfxtp_2 _52337_ (.CLK(clknet_leaf_58_wb_clk_i),
    .Q(\tholin_riscv.regs[7][5] ),
    .D(_00443_));
 sky130_as_sc_hs__dfxtp_2 _52338_ (.CLK(clknet_leaf_60_wb_clk_i),
    .Q(\tholin_riscv.regs[7][6] ),
    .D(_00444_));
 sky130_as_sc_hs__dfxtp_2 _52339_ (.CLK(clknet_leaf_50_wb_clk_i),
    .Q(\tholin_riscv.regs[7][7] ),
    .D(_00445_));
 sky130_as_sc_hs__dfxtp_2 _52340_ (.CLK(clknet_leaf_84_wb_clk_i),
    .Q(\tholin_riscv.regs[7][8] ),
    .D(_00446_));
 sky130_as_sc_hs__dfxtp_2 _52341_ (.CLK(clknet_leaf_45_wb_clk_i),
    .Q(\tholin_riscv.regs[7][9] ),
    .D(_00447_));
 sky130_as_sc_hs__dfxtp_2 _52342_ (.CLK(clknet_leaf_48_wb_clk_i),
    .Q(\tholin_riscv.regs[7][10] ),
    .D(_00448_));
 sky130_as_sc_hs__dfxtp_2 _52343_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[7][11] ),
    .D(_00449_));
 sky130_as_sc_hs__dfxtp_2 _52344_ (.CLK(clknet_leaf_31_wb_clk_i),
    .Q(\tholin_riscv.regs[7][12] ),
    .D(_00450_));
 sky130_as_sc_hs__dfxtp_2 _52345_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[7][13] ),
    .D(_00451_));
 sky130_as_sc_hs__dfxtp_2 _52346_ (.CLK(clknet_leaf_14_wb_clk_i),
    .Q(\tholin_riscv.regs[7][14] ),
    .D(_00452_));
 sky130_as_sc_hs__dfxtp_2 _52347_ (.CLK(clknet_leaf_14_wb_clk_i),
    .Q(\tholin_riscv.regs[7][15] ),
    .D(_00453_));
 sky130_as_sc_hs__dfxtp_2 _52348_ (.CLK(clknet_leaf_119_wb_clk_i),
    .Q(\tholin_riscv.regs[7][16] ),
    .D(_00454_));
 sky130_as_sc_hs__dfxtp_2 _52349_ (.CLK(clknet_leaf_102_wb_clk_i),
    .Q(\tholin_riscv.regs[7][17] ),
    .D(_00455_));
 sky130_as_sc_hs__dfxtp_2 _52350_ (.CLK(clknet_leaf_101_wb_clk_i),
    .Q(\tholin_riscv.regs[7][18] ),
    .D(_00456_));
 sky130_as_sc_hs__dfxtp_2 _52351_ (.CLK(clknet_leaf_148_wb_clk_i),
    .Q(\tholin_riscv.regs[7][19] ),
    .D(_00457_));
 sky130_as_sc_hs__dfxtp_2 _52352_ (.CLK(clknet_leaf_135_wb_clk_i),
    .Q(\tholin_riscv.regs[7][20] ),
    .D(_00458_));
 sky130_as_sc_hs__dfxtp_2 _52353_ (.CLK(clknet_leaf_108_wb_clk_i),
    .Q(\tholin_riscv.regs[7][21] ),
    .D(_00459_));
 sky130_as_sc_hs__dfxtp_2 _52354_ (.CLK(clknet_leaf_105_wb_clk_i),
    .Q(\tholin_riscv.regs[7][22] ),
    .D(_00460_));
 sky130_as_sc_hs__dfxtp_2 _52355_ (.CLK(clknet_leaf_77_wb_clk_i),
    .Q(\tholin_riscv.regs[7][23] ),
    .D(_00461_));
 sky130_as_sc_hs__dfxtp_2 _52356_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[7][24] ),
    .D(_00462_));
 sky130_as_sc_hs__dfxtp_2 _52357_ (.CLK(clknet_leaf_22_wb_clk_i),
    .Q(\tholin_riscv.regs[7][25] ),
    .D(_00463_));
 sky130_as_sc_hs__dfxtp_2 _52358_ (.CLK(clknet_leaf_33_wb_clk_i),
    .Q(\tholin_riscv.regs[7][26] ),
    .D(_00464_));
 sky130_as_sc_hs__dfxtp_2 _52359_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[7][27] ),
    .D(_00465_));
 sky130_as_sc_hs__dfxtp_2 _52360_ (.CLK(clknet_leaf_23_wb_clk_i),
    .Q(\tholin_riscv.regs[7][28] ),
    .D(_00466_));
 sky130_as_sc_hs__dfxtp_2 _52361_ (.CLK(clknet_leaf_37_wb_clk_i),
    .Q(\tholin_riscv.regs[7][29] ),
    .D(_00467_));
 sky130_as_sc_hs__dfxtp_2 _52362_ (.CLK(clknet_leaf_148_wb_clk_i),
    .Q(\tholin_riscv.regs[7][30] ),
    .D(_00468_));
 sky130_as_sc_hs__dfxtp_2 _52363_ (.CLK(clknet_leaf_98_wb_clk_i),
    .Q(\tholin_riscv.regs[7][31] ),
    .D(_00469_));
 sky130_as_sc_hs__dfxtp_2 _52364_ (.CLK(clknet_leaf_202_wb_clk_i),
    .Q(\tholin_riscv.PC[0] ),
    .D(_00470_));
 sky130_as_sc_hs__dfxtp_2 _52365_ (.CLK(clknet_leaf_133_wb_clk_i),
    .Q(\tholin_riscv.regs[6][0] ),
    .D(net695));
 sky130_as_sc_hs__dfxtp_2 _52366_ (.CLK(clknet_leaf_68_wb_clk_i),
    .Q(\tholin_riscv.regs[6][1] ),
    .D(_00472_));
 sky130_as_sc_hs__dfxtp_2 _52367_ (.CLK(clknet_leaf_65_wb_clk_i),
    .Q(\tholin_riscv.regs[6][2] ),
    .D(_00473_));
 sky130_as_sc_hs__dfxtp_2 _52368_ (.CLK(clknet_leaf_14_wb_clk_i),
    .Q(\tholin_riscv.regs[6][3] ),
    .D(_00474_));
 sky130_as_sc_hs__dfxtp_2 _52369_ (.CLK(clknet_leaf_60_wb_clk_i),
    .Q(\tholin_riscv.regs[6][4] ),
    .D(_00475_));
 sky130_as_sc_hs__dfxtp_2 _52370_ (.CLK(clknet_leaf_58_wb_clk_i),
    .Q(\tholin_riscv.regs[6][5] ),
    .D(_00476_));
 sky130_as_sc_hs__dfxtp_2 _52371_ (.CLK(clknet_leaf_60_wb_clk_i),
    .Q(\tholin_riscv.regs[6][6] ),
    .D(_00477_));
 sky130_as_sc_hs__dfxtp_2 _52372_ (.CLK(clknet_leaf_50_wb_clk_i),
    .Q(\tholin_riscv.regs[6][7] ),
    .D(_00478_));
 sky130_as_sc_hs__dfxtp_2 _52373_ (.CLK(clknet_leaf_84_wb_clk_i),
    .Q(\tholin_riscv.regs[6][8] ),
    .D(_00479_));
 sky130_as_sc_hs__dfxtp_2 _52374_ (.CLK(clknet_leaf_45_wb_clk_i),
    .Q(\tholin_riscv.regs[6][9] ),
    .D(_00480_));
 sky130_as_sc_hs__dfxtp_2 _52375_ (.CLK(clknet_leaf_48_wb_clk_i),
    .Q(\tholin_riscv.regs[6][10] ),
    .D(_00481_));
 sky130_as_sc_hs__dfxtp_2 _52376_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[6][11] ),
    .D(_00482_));
 sky130_as_sc_hs__dfxtp_2 _52377_ (.CLK(clknet_leaf_31_wb_clk_i),
    .Q(\tholin_riscv.regs[6][12] ),
    .D(_00483_));
 sky130_as_sc_hs__dfxtp_2 _52378_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[6][13] ),
    .D(_00484_));
 sky130_as_sc_hs__dfxtp_2 _52379_ (.CLK(clknet_leaf_12_wb_clk_i),
    .Q(\tholin_riscv.regs[6][14] ),
    .D(_00485_));
 sky130_as_sc_hs__dfxtp_2 _52380_ (.CLK(clknet_leaf_15_wb_clk_i),
    .Q(\tholin_riscv.regs[6][15] ),
    .D(_00486_));
 sky130_as_sc_hs__dfxtp_2 _52381_ (.CLK(clknet_leaf_85_wb_clk_i),
    .Q(\tholin_riscv.regs[6][16] ),
    .D(_00487_));
 sky130_as_sc_hs__dfxtp_2 _52382_ (.CLK(clknet_leaf_41_wb_clk_i),
    .Q(\tholin_riscv.regs[6][17] ),
    .D(_00488_));
 sky130_as_sc_hs__dfxtp_2 _52383_ (.CLK(clknet_leaf_82_wb_clk_i),
    .Q(\tholin_riscv.regs[6][18] ),
    .D(_00489_));
 sky130_as_sc_hs__dfxtp_2 _52384_ (.CLK(clknet_leaf_46_wb_clk_i),
    .Q(\tholin_riscv.regs[6][19] ),
    .D(_00490_));
 sky130_as_sc_hs__dfxtp_2 _52385_ (.CLK(clknet_leaf_73_wb_clk_i),
    .Q(\tholin_riscv.regs[6][20] ),
    .D(_00491_));
 sky130_as_sc_hs__dfxtp_2 _52386_ (.CLK(clknet_leaf_86_wb_clk_i),
    .Q(\tholin_riscv.regs[6][21] ),
    .D(_00492_));
 sky130_as_sc_hs__dfxtp_2 _52387_ (.CLK(clknet_leaf_81_wb_clk_i),
    .Q(\tholin_riscv.regs[6][22] ),
    .D(_00493_));
 sky130_as_sc_hs__dfxtp_2 _52388_ (.CLK(clknet_leaf_67_wb_clk_i),
    .Q(\tholin_riscv.regs[6][23] ),
    .D(_00494_));
 sky130_as_sc_hs__dfxtp_2 _52389_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[6][24] ),
    .D(_00495_));
 sky130_as_sc_hs__dfxtp_2 _52390_ (.CLK(clknet_leaf_22_wb_clk_i),
    .Q(\tholin_riscv.regs[6][25] ),
    .D(_00496_));
 sky130_as_sc_hs__dfxtp_2 _52391_ (.CLK(clknet_leaf_33_wb_clk_i),
    .Q(\tholin_riscv.regs[6][26] ),
    .D(_00497_));
 sky130_as_sc_hs__dfxtp_2 _52392_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[6][27] ),
    .D(_00498_));
 sky130_as_sc_hs__dfxtp_2 _52393_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[6][28] ),
    .D(_00499_));
 sky130_as_sc_hs__dfxtp_2 _52394_ (.CLK(clknet_leaf_37_wb_clk_i),
    .Q(\tholin_riscv.regs[6][29] ),
    .D(_00500_));
 sky130_as_sc_hs__dfxtp_2 _52395_ (.CLK(clknet_leaf_136_wb_clk_i),
    .Q(\tholin_riscv.regs[6][30] ),
    .D(_00501_));
 sky130_as_sc_hs__dfxtp_2 _52396_ (.CLK(clknet_leaf_153_wb_clk_i),
    .Q(\tholin_riscv.regs[6][31] ),
    .D(_00502_));
 sky130_as_sc_hs__dfxtp_2 _52397_ (.CLK(clknet_leaf_132_wb_clk_i),
    .Q(\tholin_riscv.regs[30][0] ),
    .D(net686));
 sky130_as_sc_hs__dfxtp_2 _52398_ (.CLK(clknet_leaf_126_wb_clk_i),
    .Q(\tholin_riscv.regs[30][1] ),
    .D(_00504_));
 sky130_as_sc_hs__dfxtp_2 _52399_ (.CLK(clknet_leaf_64_wb_clk_i),
    .Q(\tholin_riscv.regs[30][2] ),
    .D(_00505_));
 sky130_as_sc_hs__dfxtp_2 _52400_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[30][3] ),
    .D(_00506_));
 sky130_as_sc_hs__dfxtp_2 _52401_ (.CLK(clknet_leaf_69_wb_clk_i),
    .Q(\tholin_riscv.regs[30][4] ),
    .D(_00507_));
 sky130_as_sc_hs__dfxtp_2 _52402_ (.CLK(clknet_leaf_55_wb_clk_i),
    .Q(\tholin_riscv.regs[30][5] ),
    .D(_00508_));
 sky130_as_sc_hs__dfxtp_2 _52403_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[30][6] ),
    .D(_00509_));
 sky130_as_sc_hs__dfxtp_2 _52404_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[30][7] ),
    .D(_00510_));
 sky130_as_sc_hs__dfxtp_2 _52405_ (.CLK(clknet_leaf_79_wb_clk_i),
    .Q(\tholin_riscv.regs[30][8] ),
    .D(_00511_));
 sky130_as_sc_hs__dfxtp_2 _52406_ (.CLK(clknet_leaf_41_wb_clk_i),
    .Q(\tholin_riscv.regs[30][9] ),
    .D(_00512_));
 sky130_as_sc_hs__dfxtp_2 _52407_ (.CLK(clknet_leaf_43_wb_clk_i),
    .Q(\tholin_riscv.regs[30][10] ),
    .D(_00513_));
 sky130_as_sc_hs__dfxtp_2 _52408_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[30][11] ),
    .D(_00514_));
 sky130_as_sc_hs__dfxtp_2 _52409_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[30][12] ),
    .D(_00515_));
 sky130_as_sc_hs__dfxtp_2 _52410_ (.CLK(clknet_leaf_29_wb_clk_i),
    .Q(\tholin_riscv.regs[30][13] ),
    .D(_00516_));
 sky130_as_sc_hs__dfxtp_2 _52411_ (.CLK(clknet_leaf_19_wb_clk_i),
    .Q(\tholin_riscv.regs[30][14] ),
    .D(_00517_));
 sky130_as_sc_hs__dfxtp_2 _52412_ (.CLK(clknet_leaf_18_wb_clk_i),
    .Q(\tholin_riscv.regs[30][15] ),
    .D(_00518_));
 sky130_as_sc_hs__dfxtp_2 _52413_ (.CLK(clknet_leaf_75_wb_clk_i),
    .Q(\tholin_riscv.regs[30][16] ),
    .D(_00519_));
 sky130_as_sc_hs__dfxtp_2 _52414_ (.CLK(clknet_leaf_79_wb_clk_i),
    .Q(\tholin_riscv.regs[30][17] ),
    .D(_00520_));
 sky130_as_sc_hs__dfxtp_2 _52415_ (.CLK(clknet_leaf_122_wb_clk_i),
    .Q(\tholin_riscv.regs[30][18] ),
    .D(_00521_));
 sky130_as_sc_hs__dfxtp_2 _52416_ (.CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\tholin_riscv.regs[30][19] ),
    .D(_00522_));
 sky130_as_sc_hs__dfxtp_2 _52417_ (.CLK(clknet_leaf_72_wb_clk_i),
    .Q(\tholin_riscv.regs[30][20] ),
    .D(_00523_));
 sky130_as_sc_hs__dfxtp_2 _52418_ (.CLK(clknet_leaf_78_wb_clk_i),
    .Q(\tholin_riscv.regs[30][21] ),
    .D(_00524_));
 sky130_as_sc_hs__dfxtp_2 _52419_ (.CLK(clknet_leaf_124_wb_clk_i),
    .Q(\tholin_riscv.regs[30][22] ),
    .D(_00525_));
 sky130_as_sc_hs__dfxtp_2 _52420_ (.CLK(clknet_leaf_131_wb_clk_i),
    .Q(\tholin_riscv.regs[30][23] ),
    .D(_00526_));
 sky130_as_sc_hs__dfxtp_2 _52421_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[30][24] ),
    .D(_00527_));
 sky130_as_sc_hs__dfxtp_2 _52422_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[30][25] ),
    .D(_00528_));
 sky130_as_sc_hs__dfxtp_2 _52423_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[30][26] ),
    .D(_00529_));
 sky130_as_sc_hs__dfxtp_2 _52424_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[30][27] ),
    .D(_00530_));
 sky130_as_sc_hs__dfxtp_2 _52425_ (.CLK(clknet_leaf_91_wb_clk_i),
    .Q(\tholin_riscv.regs[30][28] ),
    .D(_00531_));
 sky130_as_sc_hs__dfxtp_2 _52426_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[30][29] ),
    .D(_00532_));
 sky130_as_sc_hs__dfxtp_2 _52427_ (.CLK(clknet_leaf_154_wb_clk_i),
    .Q(\tholin_riscv.regs[30][30] ),
    .D(_00533_));
 sky130_as_sc_hs__dfxtp_2 _52428_ (.CLK(clknet_leaf_147_wb_clk_i),
    .Q(\tholin_riscv.regs[30][31] ),
    .D(_00534_));
 sky130_as_sc_hs__dfxtp_2 _52429_ (.CLK(clknet_leaf_129_wb_clk_i),
    .Q(\tholin_riscv.regs[2][0] ),
    .D(net710));
 sky130_as_sc_hs__dfxtp_2 _52430_ (.CLK(clknet_leaf_68_wb_clk_i),
    .Q(\tholin_riscv.regs[2][1] ),
    .D(_00536_));
 sky130_as_sc_hs__dfxtp_2 _52431_ (.CLK(clknet_leaf_65_wb_clk_i),
    .Q(\tholin_riscv.regs[2][2] ),
    .D(_00537_));
 sky130_as_sc_hs__dfxtp_2 _52432_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[2][3] ),
    .D(_00538_));
 sky130_as_sc_hs__dfxtp_2 _52433_ (.CLK(clknet_leaf_70_wb_clk_i),
    .Q(\tholin_riscv.regs[2][4] ),
    .D(_00539_));
 sky130_as_sc_hs__dfxtp_2 _52434_ (.CLK(clknet_leaf_58_wb_clk_i),
    .Q(\tholin_riscv.regs[2][5] ),
    .D(_00540_));
 sky130_as_sc_hs__dfxtp_2 _52435_ (.CLK(clknet_leaf_61_wb_clk_i),
    .Q(\tholin_riscv.regs[2][6] ),
    .D(_00541_));
 sky130_as_sc_hs__dfxtp_2 _52436_ (.CLK(clknet_leaf_51_wb_clk_i),
    .Q(\tholin_riscv.regs[2][7] ),
    .D(_00542_));
 sky130_as_sc_hs__dfxtp_2 _52437_ (.CLK(clknet_leaf_83_wb_clk_i),
    .Q(\tholin_riscv.regs[2][8] ),
    .D(_00543_));
 sky130_as_sc_hs__dfxtp_2 _52438_ (.CLK(clknet_leaf_44_wb_clk_i),
    .Q(\tholin_riscv.regs[2][9] ),
    .D(_00544_));
 sky130_as_sc_hs__dfxtp_2 _52439_ (.CLK(clknet_leaf_48_wb_clk_i),
    .Q(\tholin_riscv.regs[2][10] ),
    .D(_00545_));
 sky130_as_sc_hs__dfxtp_2 _52440_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[2][11] ),
    .D(_00546_));
 sky130_as_sc_hs__dfxtp_2 _52441_ (.CLK(clknet_leaf_31_wb_clk_i),
    .Q(\tholin_riscv.regs[2][12] ),
    .D(_00547_));
 sky130_as_sc_hs__dfxtp_2 _52442_ (.CLK(clknet_leaf_32_wb_clk_i),
    .Q(\tholin_riscv.regs[2][13] ),
    .D(_00548_));
 sky130_as_sc_hs__dfxtp_2 _52443_ (.CLK(clknet_leaf_11_wb_clk_i),
    .Q(\tholin_riscv.regs[2][14] ),
    .D(_00549_));
 sky130_as_sc_hs__dfxtp_2 _52444_ (.CLK(clknet_leaf_15_wb_clk_i),
    .Q(\tholin_riscv.regs[2][15] ),
    .D(_00550_));
 sky130_as_sc_hs__dfxtp_2 _52445_ (.CLK(clknet_leaf_85_wb_clk_i),
    .Q(\tholin_riscv.regs[2][16] ),
    .D(_00551_));
 sky130_as_sc_hs__dfxtp_2 _52446_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[2][17] ),
    .D(_00552_));
 sky130_as_sc_hs__dfxtp_2 _52447_ (.CLK(clknet_leaf_83_wb_clk_i),
    .Q(\tholin_riscv.regs[2][18] ),
    .D(_00553_));
 sky130_as_sc_hs__dfxtp_2 _52448_ (.CLK(clknet_leaf_46_wb_clk_i),
    .Q(\tholin_riscv.regs[2][19] ),
    .D(_00554_));
 sky130_as_sc_hs__dfxtp_2 _52449_ (.CLK(clknet_leaf_68_wb_clk_i),
    .Q(\tholin_riscv.regs[2][20] ),
    .D(_00555_));
 sky130_as_sc_hs__dfxtp_2 _52450_ (.CLK(clknet_leaf_86_wb_clk_i),
    .Q(\tholin_riscv.regs[2][21] ),
    .D(_00556_));
 sky130_as_sc_hs__dfxtp_2 _52451_ (.CLK(clknet_leaf_82_wb_clk_i),
    .Q(\tholin_riscv.regs[2][22] ),
    .D(_00557_));
 sky130_as_sc_hs__dfxtp_2 _52452_ (.CLK(clknet_leaf_67_wb_clk_i),
    .Q(\tholin_riscv.regs[2][23] ),
    .D(_00558_));
 sky130_as_sc_hs__dfxtp_2 _52453_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[2][24] ),
    .D(_00559_));
 sky130_as_sc_hs__dfxtp_2 _52454_ (.CLK(clknet_leaf_21_wb_clk_i),
    .Q(\tholin_riscv.regs[2][25] ),
    .D(_00560_));
 sky130_as_sc_hs__dfxtp_2 _52455_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[2][26] ),
    .D(_00561_));
 sky130_as_sc_hs__dfxtp_2 _52456_ (.CLK(clknet_leaf_25_wb_clk_i),
    .Q(\tholin_riscv.regs[2][27] ),
    .D(_00562_));
 sky130_as_sc_hs__dfxtp_2 _52457_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[2][28] ),
    .D(_00563_));
 sky130_as_sc_hs__dfxtp_2 _52458_ (.CLK(clknet_leaf_36_wb_clk_i),
    .Q(\tholin_riscv.regs[2][29] ),
    .D(_00564_));
 sky130_as_sc_hs__dfxtp_2 _52459_ (.CLK(clknet_leaf_136_wb_clk_i),
    .Q(\tholin_riscv.regs[2][30] ),
    .D(_00565_));
 sky130_as_sc_hs__dfxtp_2 _52460_ (.CLK(clknet_leaf_97_wb_clk_i),
    .Q(\tholin_riscv.regs[2][31] ),
    .D(_00566_));
 sky130_as_sc_hs__dfxtp_2 _52461_ (.CLK(clknet_leaf_131_wb_clk_i),
    .Q(\tholin_riscv.regs[28][0] ),
    .D(net662));
 sky130_as_sc_hs__dfxtp_2 _52462_ (.CLK(clknet_leaf_126_wb_clk_i),
    .Q(\tholin_riscv.regs[28][1] ),
    .D(_00568_));
 sky130_as_sc_hs__dfxtp_2 _52463_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[28][2] ),
    .D(_00569_));
 sky130_as_sc_hs__dfxtp_2 _52464_ (.CLK(clknet_leaf_55_wb_clk_i),
    .Q(\tholin_riscv.regs[28][3] ),
    .D(_00570_));
 sky130_as_sc_hs__dfxtp_2 _52465_ (.CLK(clknet_leaf_69_wb_clk_i),
    .Q(\tholin_riscv.regs[28][4] ),
    .D(_00571_));
 sky130_as_sc_hs__dfxtp_2 _52466_ (.CLK(clknet_leaf_54_wb_clk_i),
    .Q(\tholin_riscv.regs[28][5] ),
    .D(_00572_));
 sky130_as_sc_hs__dfxtp_2 _52467_ (.CLK(clknet_leaf_62_wb_clk_i),
    .Q(\tholin_riscv.regs[28][6] ),
    .D(_00573_));
 sky130_as_sc_hs__dfxtp_2 _52468_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[28][7] ),
    .D(_00574_));
 sky130_as_sc_hs__dfxtp_2 _52469_ (.CLK(clknet_leaf_80_wb_clk_i),
    .Q(\tholin_riscv.regs[28][8] ),
    .D(_00575_));
 sky130_as_sc_hs__dfxtp_2 _52470_ (.CLK(clknet_leaf_44_wb_clk_i),
    .Q(\tholin_riscv.regs[28][9] ),
    .D(_00576_));
 sky130_as_sc_hs__dfxtp_2 _52471_ (.CLK(clknet_leaf_49_wb_clk_i),
    .Q(\tholin_riscv.regs[28][10] ),
    .D(_00577_));
 sky130_as_sc_hs__dfxtp_2 _52472_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[28][11] ),
    .D(_00578_));
 sky130_as_sc_hs__dfxtp_2 _52473_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[28][12] ),
    .D(_00579_));
 sky130_as_sc_hs__dfxtp_2 _52474_ (.CLK(clknet_leaf_28_wb_clk_i),
    .Q(\tholin_riscv.regs[28][13] ),
    .D(_00580_));
 sky130_as_sc_hs__dfxtp_2 _52475_ (.CLK(clknet_leaf_19_wb_clk_i),
    .Q(\tholin_riscv.regs[28][14] ),
    .D(_00581_));
 sky130_as_sc_hs__dfxtp_2 _52476_ (.CLK(clknet_leaf_18_wb_clk_i),
    .Q(\tholin_riscv.regs[28][15] ),
    .D(_00582_));
 sky130_as_sc_hs__dfxtp_2 _52477_ (.CLK(clknet_leaf_75_wb_clk_i),
    .Q(\tholin_riscv.regs[28][16] ),
    .D(_00583_));
 sky130_as_sc_hs__dfxtp_2 _52478_ (.CLK(clknet_leaf_79_wb_clk_i),
    .Q(\tholin_riscv.regs[28][17] ),
    .D(_00584_));
 sky130_as_sc_hs__dfxtp_2 _52479_ (.CLK(clknet_leaf_74_wb_clk_i),
    .Q(\tholin_riscv.regs[28][18] ),
    .D(_00585_));
 sky130_as_sc_hs__dfxtp_2 _52480_ (.CLK(clknet_leaf_74_wb_clk_i),
    .Q(\tholin_riscv.regs[28][19] ),
    .D(_00586_));
 sky130_as_sc_hs__dfxtp_2 _52481_ (.CLK(clknet_leaf_71_wb_clk_i),
    .Q(\tholin_riscv.regs[28][20] ),
    .D(_00587_));
 sky130_as_sc_hs__dfxtp_2 _52482_ (.CLK(clknet_leaf_78_wb_clk_i),
    .Q(\tholin_riscv.regs[28][21] ),
    .D(_00588_));
 sky130_as_sc_hs__dfxtp_2 _52483_ (.CLK(clknet_leaf_123_wb_clk_i),
    .Q(\tholin_riscv.regs[28][22] ),
    .D(_00589_));
 sky130_as_sc_hs__dfxtp_2 _52484_ (.CLK(clknet_leaf_131_wb_clk_i),
    .Q(\tholin_riscv.regs[28][23] ),
    .D(_00590_));
 sky130_as_sc_hs__dfxtp_2 _52485_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[28][24] ),
    .D(_00591_));
 sky130_as_sc_hs__dfxtp_2 _52486_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[28][25] ),
    .D(_00592_));
 sky130_as_sc_hs__dfxtp_2 _52487_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[28][26] ),
    .D(_00593_));
 sky130_as_sc_hs__dfxtp_2 _52488_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[28][27] ),
    .D(_00594_));
 sky130_as_sc_hs__dfxtp_2 _52489_ (.CLK(clknet_leaf_90_wb_clk_i),
    .Q(\tholin_riscv.regs[28][28] ),
    .D(_00595_));
 sky130_as_sc_hs__dfxtp_2 _52490_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[28][29] ),
    .D(_00596_));
 sky130_as_sc_hs__dfxtp_2 _52491_ (.CLK(clknet_leaf_151_wb_clk_i),
    .Q(\tholin_riscv.regs[28][30] ),
    .D(_00597_));
 sky130_as_sc_hs__dfxtp_2 _52492_ (.CLK(clknet_leaf_121_wb_clk_i),
    .Q(\tholin_riscv.regs[28][31] ),
    .D(_00598_));
 sky130_as_sc_hs__dfxtp_2 _52493_ (.CLK(clknet_leaf_131_wb_clk_i),
    .Q(\tholin_riscv.regs[27][0] ),
    .D(net743));
 sky130_as_sc_hs__dfxtp_2 _52494_ (.CLK(clknet_leaf_126_wb_clk_i),
    .Q(\tholin_riscv.regs[27][1] ),
    .D(_00600_));
 sky130_as_sc_hs__dfxtp_2 _52495_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[27][2] ),
    .D(_00601_));
 sky130_as_sc_hs__dfxtp_2 _52496_ (.CLK(clknet_leaf_9_wb_clk_i),
    .Q(\tholin_riscv.regs[27][3] ),
    .D(_00602_));
 sky130_as_sc_hs__dfxtp_2 _52497_ (.CLK(clknet_leaf_111_wb_clk_i),
    .Q(\tholin_riscv.regs[27][4] ),
    .D(_00603_));
 sky130_as_sc_hs__dfxtp_2 _52498_ (.CLK(clknet_leaf_53_wb_clk_i),
    .Q(\tholin_riscv.regs[27][5] ),
    .D(_00604_));
 sky130_as_sc_hs__dfxtp_2 _52499_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[27][6] ),
    .D(_00605_));
 sky130_as_sc_hs__dfxtp_2 _52500_ (.CLK(clknet_leaf_53_wb_clk_i),
    .Q(\tholin_riscv.regs[27][7] ),
    .D(_00606_));
 sky130_as_sc_hs__dfxtp_2 _52501_ (.CLK(clknet_leaf_80_wb_clk_i),
    .Q(\tholin_riscv.regs[27][8] ),
    .D(_00607_));
 sky130_as_sc_hs__dfxtp_2 _52502_ (.CLK(clknet_leaf_43_wb_clk_i),
    .Q(\tholin_riscv.regs[27][9] ),
    .D(_00608_));
 sky130_as_sc_hs__dfxtp_2 _52503_ (.CLK(clknet_leaf_37_wb_clk_i),
    .Q(\tholin_riscv.regs[27][10] ),
    .D(_00609_));
 sky130_as_sc_hs__dfxtp_2 _52504_ (.CLK(clknet_leaf_28_wb_clk_i),
    .Q(\tholin_riscv.regs[27][11] ),
    .D(_00610_));
 sky130_as_sc_hs__dfxtp_2 _52505_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[27][12] ),
    .D(_00611_));
 sky130_as_sc_hs__dfxtp_2 _52506_ (.CLK(clknet_leaf_22_wb_clk_i),
    .Q(\tholin_riscv.regs[27][13] ),
    .D(_00612_));
 sky130_as_sc_hs__dfxtp_2 _52507_ (.CLK(clknet_leaf_17_wb_clk_i),
    .Q(\tholin_riscv.regs[27][14] ),
    .D(_00613_));
 sky130_as_sc_hs__dfxtp_2 _52508_ (.CLK(clknet_leaf_17_wb_clk_i),
    .Q(\tholin_riscv.regs[27][15] ),
    .D(_00614_));
 sky130_as_sc_hs__dfxtp_2 _52509_ (.CLK(clknet_leaf_106_wb_clk_i),
    .Q(\tholin_riscv.regs[27][16] ),
    .D(_00615_));
 sky130_as_sc_hs__dfxtp_2 _52510_ (.CLK(clknet_leaf_103_wb_clk_i),
    .Q(\tholin_riscv.regs[27][17] ),
    .D(_00616_));
 sky130_as_sc_hs__dfxtp_2 _52511_ (.CLK(clknet_leaf_115_wb_clk_i),
    .Q(\tholin_riscv.regs[27][18] ),
    .D(_00617_));
 sky130_as_sc_hs__dfxtp_2 _52512_ (.CLK(clknet_leaf_115_wb_clk_i),
    .Q(\tholin_riscv.regs[27][19] ),
    .D(_00618_));
 sky130_as_sc_hs__dfxtp_2 _52513_ (.CLK(clknet_leaf_107_wb_clk_i),
    .Q(\tholin_riscv.regs[27][20] ),
    .D(_00619_));
 sky130_as_sc_hs__dfxtp_2 _52514_ (.CLK(clknet_leaf_115_wb_clk_i),
    .Q(\tholin_riscv.regs[27][21] ),
    .D(_00620_));
 sky130_as_sc_hs__dfxtp_2 _52515_ (.CLK(clknet_leaf_116_wb_clk_i),
    .Q(\tholin_riscv.regs[27][22] ),
    .D(_00621_));
 sky130_as_sc_hs__dfxtp_2 _52516_ (.CLK(clknet_leaf_101_wb_clk_i),
    .Q(\tholin_riscv.regs[27][23] ),
    .D(_00622_));
 sky130_as_sc_hs__dfxtp_2 _52517_ (.CLK(clknet_leaf_39_wb_clk_i),
    .Q(\tholin_riscv.regs[27][24] ),
    .D(_00623_));
 sky130_as_sc_hs__dfxtp_2 _52518_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[27][25] ),
    .D(_00624_));
 sky130_as_sc_hs__dfxtp_2 _52519_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[27][26] ),
    .D(_00625_));
 sky130_as_sc_hs__dfxtp_2 _52520_ (.CLK(clknet_leaf_91_wb_clk_i),
    .Q(\tholin_riscv.regs[27][27] ),
    .D(_00626_));
 sky130_as_sc_hs__dfxtp_2 _52521_ (.CLK(clknet_leaf_91_wb_clk_i),
    .Q(\tholin_riscv.regs[27][28] ),
    .D(_00627_));
 sky130_as_sc_hs__dfxtp_2 _52522_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[27][29] ),
    .D(_00628_));
 sky130_as_sc_hs__dfxtp_2 _52523_ (.CLK(clknet_leaf_99_wb_clk_i),
    .Q(\tholin_riscv.regs[27][30] ),
    .D(_00629_));
 sky130_as_sc_hs__dfxtp_2 _52524_ (.CLK(clknet_leaf_135_wb_clk_i),
    .Q(\tholin_riscv.regs[27][31] ),
    .D(_00630_));
 sky130_as_sc_hs__dfxtp_2 _52525_ (.CLK(clknet_leaf_131_wb_clk_i),
    .Q(\tholin_riscv.regs[26][0] ),
    .D(net734));
 sky130_as_sc_hs__dfxtp_2 _52526_ (.CLK(clknet_leaf_126_wb_clk_i),
    .Q(\tholin_riscv.regs[26][1] ),
    .D(_00632_));
 sky130_as_sc_hs__dfxtp_2 _52527_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[26][2] ),
    .D(_00633_));
 sky130_as_sc_hs__dfxtp_2 _52528_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[26][3] ),
    .D(_00634_));
 sky130_as_sc_hs__dfxtp_2 _52529_ (.CLK(clknet_leaf_69_wb_clk_i),
    .Q(\tholin_riscv.regs[26][4] ),
    .D(_00635_));
 sky130_as_sc_hs__dfxtp_2 _52530_ (.CLK(clknet_leaf_54_wb_clk_i),
    .Q(\tholin_riscv.regs[26][5] ),
    .D(_00636_));
 sky130_as_sc_hs__dfxtp_2 _52531_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[26][6] ),
    .D(_00637_));
 sky130_as_sc_hs__dfxtp_2 _52532_ (.CLK(clknet_leaf_53_wb_clk_i),
    .Q(\tholin_riscv.regs[26][7] ),
    .D(_00638_));
 sky130_as_sc_hs__dfxtp_2 _52533_ (.CLK(clknet_leaf_80_wb_clk_i),
    .Q(\tholin_riscv.regs[26][8] ),
    .D(_00639_));
 sky130_as_sc_hs__dfxtp_2 _52534_ (.CLK(clknet_leaf_43_wb_clk_i),
    .Q(\tholin_riscv.regs[26][9] ),
    .D(_00640_));
 sky130_as_sc_hs__dfxtp_2 _52535_ (.CLK(clknet_leaf_37_wb_clk_i),
    .Q(\tholin_riscv.regs[26][10] ),
    .D(_00641_));
 sky130_as_sc_hs__dfxtp_2 _52536_ (.CLK(clknet_leaf_28_wb_clk_i),
    .Q(\tholin_riscv.regs[26][11] ),
    .D(_00642_));
 sky130_as_sc_hs__dfxtp_2 _52537_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[26][12] ),
    .D(_00643_));
 sky130_as_sc_hs__dfxtp_2 _52538_ (.CLK(clknet_leaf_27_wb_clk_i),
    .Q(\tholin_riscv.regs[26][13] ),
    .D(_00644_));
 sky130_as_sc_hs__dfxtp_2 _52539_ (.CLK(clknet_leaf_17_wb_clk_i),
    .Q(\tholin_riscv.regs[26][14] ),
    .D(_00645_));
 sky130_as_sc_hs__dfxtp_2 _52540_ (.CLK(clknet_leaf_17_wb_clk_i),
    .Q(\tholin_riscv.regs[26][15] ),
    .D(_00646_));
 sky130_as_sc_hs__dfxtp_2 _52541_ (.CLK(clknet_leaf_78_wb_clk_i),
    .Q(\tholin_riscv.regs[26][16] ),
    .D(_00647_));
 sky130_as_sc_hs__dfxtp_2 _52542_ (.CLK(clknet_leaf_78_wb_clk_i),
    .Q(\tholin_riscv.regs[26][17] ),
    .D(_00648_));
 sky130_as_sc_hs__dfxtp_2 _52543_ (.CLK(clknet_leaf_122_wb_clk_i),
    .Q(\tholin_riscv.regs[26][18] ),
    .D(_00649_));
 sky130_as_sc_hs__dfxtp_2 _52544_ (.CLK(clknet_leaf_73_wb_clk_i),
    .Q(\tholin_riscv.regs[26][19] ),
    .D(_00650_));
 sky130_as_sc_hs__dfxtp_2 _52545_ (.CLK(clknet_leaf_71_wb_clk_i),
    .Q(\tholin_riscv.regs[26][20] ),
    .D(_00651_));
 sky130_as_sc_hs__dfxtp_2 _52546_ (.CLK(clknet_leaf_81_wb_clk_i),
    .Q(\tholin_riscv.regs[26][21] ),
    .D(_00652_));
 sky130_as_sc_hs__dfxtp_2 _52547_ (.CLK(clknet_leaf_124_wb_clk_i),
    .Q(\tholin_riscv.regs[26][22] ),
    .D(_00653_));
 sky130_as_sc_hs__dfxtp_2 _52548_ (.CLK(clknet_leaf_129_wb_clk_i),
    .Q(\tholin_riscv.regs[26][23] ),
    .D(_00654_));
 sky130_as_sc_hs__dfxtp_2 _52549_ (.CLK(clknet_leaf_39_wb_clk_i),
    .Q(\tholin_riscv.regs[26][24] ),
    .D(_00655_));
 sky130_as_sc_hs__dfxtp_2 _52550_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[26][25] ),
    .D(_00656_));
 sky130_as_sc_hs__dfxtp_2 _52551_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[26][26] ),
    .D(_00657_));
 sky130_as_sc_hs__dfxtp_2 _52552_ (.CLK(clknet_leaf_91_wb_clk_i),
    .Q(\tholin_riscv.regs[26][27] ),
    .D(_00658_));
 sky130_as_sc_hs__dfxtp_2 _52553_ (.CLK(clknet_leaf_91_wb_clk_i),
    .Q(\tholin_riscv.regs[26][28] ),
    .D(_00659_));
 sky130_as_sc_hs__dfxtp_2 _52554_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[26][29] ),
    .D(_00660_));
 sky130_as_sc_hs__dfxtp_2 _52555_ (.CLK(clknet_leaf_117_wb_clk_i),
    .Q(\tholin_riscv.regs[26][30] ),
    .D(_00661_));
 sky130_as_sc_hs__dfxtp_2 _52556_ (.CLK(clknet_leaf_146_wb_clk_i),
    .Q(\tholin_riscv.regs[26][31] ),
    .D(_00662_));
 sky130_as_sc_hs__dfxtp_2 _52557_ (.CLK(clknet_leaf_66_wb_clk_i),
    .Q(\tholin_riscv.regs[25][0] ),
    .D(net659));
 sky130_as_sc_hs__dfxtp_2 _52558_ (.CLK(clknet_leaf_126_wb_clk_i),
    .Q(\tholin_riscv.regs[25][1] ),
    .D(_00664_));
 sky130_as_sc_hs__dfxtp_2 _52559_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[25][2] ),
    .D(_00665_));
 sky130_as_sc_hs__dfxtp_2 _52560_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[25][3] ),
    .D(_00666_));
 sky130_as_sc_hs__dfxtp_2 _52561_ (.CLK(clknet_leaf_102_wb_clk_i),
    .Q(\tholin_riscv.regs[25][4] ),
    .D(_00667_));
 sky130_as_sc_hs__dfxtp_2 _52562_ (.CLK(clknet_leaf_54_wb_clk_i),
    .Q(\tholin_riscv.regs[25][5] ),
    .D(_00668_));
 sky130_as_sc_hs__dfxtp_2 _52563_ (.CLK(clknet_leaf_62_wb_clk_i),
    .Q(\tholin_riscv.regs[25][6] ),
    .D(_00669_));
 sky130_as_sc_hs__dfxtp_2 _52564_ (.CLK(clknet_leaf_53_wb_clk_i),
    .Q(\tholin_riscv.regs[25][7] ),
    .D(_00670_));
 sky130_as_sc_hs__dfxtp_2 _52565_ (.CLK(clknet_leaf_80_wb_clk_i),
    .Q(\tholin_riscv.regs[25][8] ),
    .D(_00671_));
 sky130_as_sc_hs__dfxtp_2 _52566_ (.CLK(clknet_leaf_43_wb_clk_i),
    .Q(\tholin_riscv.regs[25][9] ),
    .D(_00672_));
 sky130_as_sc_hs__dfxtp_2 _52567_ (.CLK(clknet_leaf_37_wb_clk_i),
    .Q(\tholin_riscv.regs[25][10] ),
    .D(_00673_));
 sky130_as_sc_hs__dfxtp_2 _52568_ (.CLK(clknet_leaf_29_wb_clk_i),
    .Q(\tholin_riscv.regs[25][11] ),
    .D(_00674_));
 sky130_as_sc_hs__dfxtp_2 _52569_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[25][12] ),
    .D(_00675_));
 sky130_as_sc_hs__dfxtp_2 _52570_ (.CLK(clknet_leaf_22_wb_clk_i),
    .Q(\tholin_riscv.regs[25][13] ),
    .D(_00676_));
 sky130_as_sc_hs__dfxtp_2 _52571_ (.CLK(clknet_leaf_17_wb_clk_i),
    .Q(\tholin_riscv.regs[25][14] ),
    .D(_00677_));
 sky130_as_sc_hs__dfxtp_2 _52572_ (.CLK(clknet_leaf_17_wb_clk_i),
    .Q(\tholin_riscv.regs[25][15] ),
    .D(_00678_));
 sky130_as_sc_hs__dfxtp_2 _52573_ (.CLK(clknet_leaf_116_wb_clk_i),
    .Q(\tholin_riscv.regs[25][16] ),
    .D(_00679_));
 sky130_as_sc_hs__dfxtp_2 _52574_ (.CLK(clknet_leaf_94_wb_clk_i),
    .Q(\tholin_riscv.regs[25][17] ),
    .D(_00680_));
 sky130_as_sc_hs__dfxtp_2 _52575_ (.CLK(clknet_leaf_105_wb_clk_i),
    .Q(\tholin_riscv.regs[25][18] ),
    .D(_00681_));
 sky130_as_sc_hs__dfxtp_2 _52576_ (.CLK(clknet_leaf_118_wb_clk_i),
    .Q(\tholin_riscv.regs[25][19] ),
    .D(_00682_));
 sky130_as_sc_hs__dfxtp_2 _52577_ (.CLK(clknet_leaf_101_wb_clk_i),
    .Q(\tholin_riscv.regs[25][20] ),
    .D(_00683_));
 sky130_as_sc_hs__dfxtp_2 _52578_ (.CLK(clknet_leaf_148_wb_clk_i),
    .Q(\tholin_riscv.regs[25][21] ),
    .D(_00684_));
 sky130_as_sc_hs__dfxtp_2 _52579_ (.CLK(clknet_leaf_103_wb_clk_i),
    .Q(\tholin_riscv.regs[25][22] ),
    .D(_00685_));
 sky130_as_sc_hs__dfxtp_2 _52580_ (.CLK(clknet_leaf_154_wb_clk_i),
    .Q(\tholin_riscv.regs[25][23] ),
    .D(_00686_));
 sky130_as_sc_hs__dfxtp_2 _52581_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[25][24] ),
    .D(_00687_));
 sky130_as_sc_hs__dfxtp_2 _52582_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[25][25] ),
    .D(_00688_));
 sky130_as_sc_hs__dfxtp_2 _52583_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[25][26] ),
    .D(_00689_));
 sky130_as_sc_hs__dfxtp_2 _52584_ (.CLK(clknet_leaf_90_wb_clk_i),
    .Q(\tholin_riscv.regs[25][27] ),
    .D(_00690_));
 sky130_as_sc_hs__dfxtp_2 _52585_ (.CLK(clknet_leaf_90_wb_clk_i),
    .Q(\tholin_riscv.regs[25][28] ),
    .D(_00691_));
 sky130_as_sc_hs__dfxtp_2 _52586_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[25][29] ),
    .D(_00692_));
 sky130_as_sc_hs__dfxtp_2 _52587_ (.CLK(clknet_leaf_126_wb_clk_i),
    .Q(\tholin_riscv.regs[25][30] ),
    .D(_00693_));
 sky130_as_sc_hs__dfxtp_2 _52588_ (.CLK(clknet_leaf_149_wb_clk_i),
    .Q(\tholin_riscv.regs[25][31] ),
    .D(_00694_));
 sky130_as_sc_hs__dfxtp_2 _52589_ (.CLK(clknet_leaf_131_wb_clk_i),
    .Q(\tholin_riscv.regs[24][0] ),
    .D(net665));
 sky130_as_sc_hs__dfxtp_2 _52590_ (.CLK(clknet_leaf_126_wb_clk_i),
    .Q(\tholin_riscv.regs[24][1] ),
    .D(_00696_));
 sky130_as_sc_hs__dfxtp_2 _52591_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[24][2] ),
    .D(_00697_));
 sky130_as_sc_hs__dfxtp_2 _52592_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[24][3] ),
    .D(_00698_));
 sky130_as_sc_hs__dfxtp_2 _52593_ (.CLK(clknet_leaf_69_wb_clk_i),
    .Q(\tholin_riscv.regs[24][4] ),
    .D(_00699_));
 sky130_as_sc_hs__dfxtp_2 _52594_ (.CLK(clknet_leaf_54_wb_clk_i),
    .Q(\tholin_riscv.regs[24][5] ),
    .D(_00700_));
 sky130_as_sc_hs__dfxtp_2 _52595_ (.CLK(clknet_leaf_62_wb_clk_i),
    .Q(\tholin_riscv.regs[24][6] ),
    .D(_00701_));
 sky130_as_sc_hs__dfxtp_2 _52596_ (.CLK(clknet_leaf_53_wb_clk_i),
    .Q(\tholin_riscv.regs[24][7] ),
    .D(_00702_));
 sky130_as_sc_hs__dfxtp_2 _52597_ (.CLK(clknet_leaf_80_wb_clk_i),
    .Q(\tholin_riscv.regs[24][8] ),
    .D(_00703_));
 sky130_as_sc_hs__dfxtp_2 _52598_ (.CLK(clknet_leaf_43_wb_clk_i),
    .Q(\tholin_riscv.regs[24][9] ),
    .D(_00704_));
 sky130_as_sc_hs__dfxtp_2 _52599_ (.CLK(clknet_leaf_37_wb_clk_i),
    .Q(\tholin_riscv.regs[24][10] ),
    .D(_00705_));
 sky130_as_sc_hs__dfxtp_2 _52600_ (.CLK(clknet_leaf_29_wb_clk_i),
    .Q(\tholin_riscv.regs[24][11] ),
    .D(_00706_));
 sky130_as_sc_hs__dfxtp_2 _52601_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[24][12] ),
    .D(_00707_));
 sky130_as_sc_hs__dfxtp_2 _52602_ (.CLK(clknet_leaf_22_wb_clk_i),
    .Q(\tholin_riscv.regs[24][13] ),
    .D(_00708_));
 sky130_as_sc_hs__dfxtp_2 _52603_ (.CLK(clknet_leaf_16_wb_clk_i),
    .Q(\tholin_riscv.regs[24][14] ),
    .D(_00709_));
 sky130_as_sc_hs__dfxtp_2 _52604_ (.CLK(clknet_leaf_17_wb_clk_i),
    .Q(\tholin_riscv.regs[24][15] ),
    .D(_00710_));
 sky130_as_sc_hs__dfxtp_2 _52605_ (.CLK(clknet_leaf_78_wb_clk_i),
    .Q(\tholin_riscv.regs[24][16] ),
    .D(_00711_));
 sky130_as_sc_hs__dfxtp_2 _52606_ (.CLK(clknet_leaf_79_wb_clk_i),
    .Q(\tholin_riscv.regs[24][17] ),
    .D(_00712_));
 sky130_as_sc_hs__dfxtp_2 _52607_ (.CLK(clknet_leaf_122_wb_clk_i),
    .Q(\tholin_riscv.regs[24][18] ),
    .D(_00713_));
 sky130_as_sc_hs__dfxtp_2 _52608_ (.CLK(clknet_leaf_74_wb_clk_i),
    .Q(\tholin_riscv.regs[24][19] ),
    .D(_00714_));
 sky130_as_sc_hs__dfxtp_2 _52609_ (.CLK(clknet_leaf_72_wb_clk_i),
    .Q(\tholin_riscv.regs[24][20] ),
    .D(_00715_));
 sky130_as_sc_hs__dfxtp_2 _52610_ (.CLK(clknet_leaf_81_wb_clk_i),
    .Q(\tholin_riscv.regs[24][21] ),
    .D(_00716_));
 sky130_as_sc_hs__dfxtp_2 _52611_ (.CLK(clknet_leaf_123_wb_clk_i),
    .Q(\tholin_riscv.regs[24][22] ),
    .D(_00717_));
 sky130_as_sc_hs__dfxtp_2 _52612_ (.CLK(clknet_leaf_129_wb_clk_i),
    .Q(\tholin_riscv.regs[24][23] ),
    .D(_00718_));
 sky130_as_sc_hs__dfxtp_2 _52613_ (.CLK(clknet_leaf_39_wb_clk_i),
    .Q(\tholin_riscv.regs[24][24] ),
    .D(_00719_));
 sky130_as_sc_hs__dfxtp_2 _52614_ (.CLK(clknet_leaf_79_wb_clk_i),
    .Q(\tholin_riscv.regs[24][25] ),
    .D(_00720_));
 sky130_as_sc_hs__dfxtp_2 _52615_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[24][26] ),
    .D(_00721_));
 sky130_as_sc_hs__dfxtp_2 _52616_ (.CLK(clknet_leaf_90_wb_clk_i),
    .Q(\tholin_riscv.regs[24][27] ),
    .D(_00722_));
 sky130_as_sc_hs__dfxtp_2 _52617_ (.CLK(clknet_leaf_90_wb_clk_i),
    .Q(\tholin_riscv.regs[24][28] ),
    .D(_00723_));
 sky130_as_sc_hs__dfxtp_2 _52618_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[24][29] ),
    .D(_00724_));
 sky130_as_sc_hs__dfxtp_2 _52619_ (.CLK(clknet_leaf_97_wb_clk_i),
    .Q(\tholin_riscv.regs[24][30] ),
    .D(_00725_));
 sky130_as_sc_hs__dfxtp_2 _52620_ (.CLK(clknet_leaf_151_wb_clk_i),
    .Q(\tholin_riscv.regs[24][31] ),
    .D(_00726_));
 sky130_as_sc_hs__dfxtp_2 _52621_ (.CLK(clknet_leaf_196_wb_clk_i),
    .Q(\tholin_riscv.regs[23][0] ),
    .D(net716));
 sky130_as_sc_hs__dfxtp_2 _52622_ (.CLK(clknet_leaf_127_wb_clk_i),
    .Q(\tholin_riscv.regs[23][1] ),
    .D(_00728_));
 sky130_as_sc_hs__dfxtp_2 _52623_ (.CLK(clknet_leaf_7_wb_clk_i),
    .Q(\tholin_riscv.regs[23][2] ),
    .D(_00729_));
 sky130_as_sc_hs__dfxtp_2 _52624_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[23][3] ),
    .D(_00730_));
 sky130_as_sc_hs__dfxtp_2 _52625_ (.CLK(clknet_leaf_107_wb_clk_i),
    .Q(\tholin_riscv.regs[23][4] ),
    .D(_00731_));
 sky130_as_sc_hs__dfxtp_2 _52626_ (.CLK(clknet_leaf_57_wb_clk_i),
    .Q(\tholin_riscv.regs[23][5] ),
    .D(_00732_));
 sky130_as_sc_hs__dfxtp_2 _52627_ (.CLK(clknet_leaf_56_wb_clk_i),
    .Q(\tholin_riscv.regs[23][6] ),
    .D(_00733_));
 sky130_as_sc_hs__dfxtp_2 _52628_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[23][7] ),
    .D(_00734_));
 sky130_as_sc_hs__dfxtp_2 _52629_ (.CLK(clknet_leaf_85_wb_clk_i),
    .Q(\tholin_riscv.regs[23][8] ),
    .D(_00735_));
 sky130_as_sc_hs__dfxtp_2 _52630_ (.CLK(clknet_leaf_42_wb_clk_i),
    .Q(\tholin_riscv.regs[23][9] ),
    .D(_00736_));
 sky130_as_sc_hs__dfxtp_2 _52631_ (.CLK(clknet_leaf_31_wb_clk_i),
    .Q(\tholin_riscv.regs[23][10] ),
    .D(_00737_));
 sky130_as_sc_hs__dfxtp_2 _52632_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[23][11] ),
    .D(_00738_));
 sky130_as_sc_hs__dfxtp_2 _52633_ (.CLK(clknet_leaf_28_wb_clk_i),
    .Q(\tholin_riscv.regs[23][12] ),
    .D(_00739_));
 sky130_as_sc_hs__dfxtp_2 _52634_ (.CLK(clknet_leaf_21_wb_clk_i),
    .Q(\tholin_riscv.regs[23][13] ),
    .D(_00740_));
 sky130_as_sc_hs__dfxtp_2 _52635_ (.CLK(clknet_leaf_17_wb_clk_i),
    .Q(\tholin_riscv.regs[23][14] ),
    .D(_00741_));
 sky130_as_sc_hs__dfxtp_2 _52636_ (.CLK(clknet_leaf_16_wb_clk_i),
    .Q(\tholin_riscv.regs[23][15] ),
    .D(_00742_));
 sky130_as_sc_hs__dfxtp_2 _52637_ (.CLK(clknet_leaf_149_wb_clk_i),
    .Q(\tholin_riscv.regs[23][16] ),
    .D(_00743_));
 sky130_as_sc_hs__dfxtp_2 _52638_ (.CLK(clknet_leaf_107_wb_clk_i),
    .Q(\tholin_riscv.regs[23][17] ),
    .D(_00744_));
 sky130_as_sc_hs__dfxtp_2 _52639_ (.CLK(clknet_leaf_100_wb_clk_i),
    .Q(\tholin_riscv.regs[23][18] ),
    .D(_00745_));
 sky130_as_sc_hs__dfxtp_2 _52640_ (.CLK(clknet_leaf_149_wb_clk_i),
    .Q(\tholin_riscv.regs[23][19] ),
    .D(_00746_));
 sky130_as_sc_hs__dfxtp_2 _52641_ (.CLK(clknet_leaf_118_wb_clk_i),
    .Q(\tholin_riscv.regs[23][20] ),
    .D(_00747_));
 sky130_as_sc_hs__dfxtp_2 _52642_ (.CLK(clknet_leaf_94_wb_clk_i),
    .Q(\tholin_riscv.regs[23][21] ),
    .D(_00748_));
 sky130_as_sc_hs__dfxtp_2 _52643_ (.CLK(clknet_leaf_103_wb_clk_i),
    .Q(\tholin_riscv.regs[23][22] ),
    .D(_00749_));
 sky130_as_sc_hs__dfxtp_2 _52644_ (.CLK(clknet_leaf_111_wb_clk_i),
    .Q(\tholin_riscv.regs[23][23] ),
    .D(_00750_));
 sky130_as_sc_hs__dfxtp_2 _52645_ (.CLK(clknet_leaf_42_wb_clk_i),
    .Q(\tholin_riscv.regs[23][24] ),
    .D(_00751_));
 sky130_as_sc_hs__dfxtp_2 _52646_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[23][25] ),
    .D(_00752_));
 sky130_as_sc_hs__dfxtp_2 _52647_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[23][26] ),
    .D(_00753_));
 sky130_as_sc_hs__dfxtp_2 _52648_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[23][27] ),
    .D(_00754_));
 sky130_as_sc_hs__dfxtp_2 _52649_ (.CLK(clknet_leaf_89_wb_clk_i),
    .Q(\tholin_riscv.regs[23][28] ),
    .D(_00755_));
 sky130_as_sc_hs__dfxtp_2 _52650_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[23][29] ),
    .D(_00756_));
 sky130_as_sc_hs__dfxtp_2 _52651_ (.CLK(clknet_leaf_147_wb_clk_i),
    .Q(\tholin_riscv.regs[23][30] ),
    .D(_00757_));
 sky130_as_sc_hs__dfxtp_2 _52652_ (.CLK(clknet_leaf_147_wb_clk_i),
    .Q(\tholin_riscv.regs[23][31] ),
    .D(_00758_));
 sky130_as_sc_hs__dfxtp_2 _52653_ (.CLK(clknet_leaf_195_wb_clk_i),
    .Q(\tholin_riscv.regs[22][0] ),
    .D(net701));
 sky130_as_sc_hs__dfxtp_2 _52654_ (.CLK(clknet_leaf_127_wb_clk_i),
    .Q(\tholin_riscv.regs[22][1] ),
    .D(_00760_));
 sky130_as_sc_hs__dfxtp_2 _52655_ (.CLK(clknet_leaf_7_wb_clk_i),
    .Q(\tholin_riscv.regs[22][2] ),
    .D(_00761_));
 sky130_as_sc_hs__dfxtp_2 _52656_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[22][3] ),
    .D(_00762_));
 sky130_as_sc_hs__dfxtp_2 _52657_ (.CLK(clknet_leaf_67_wb_clk_i),
    .Q(\tholin_riscv.regs[22][4] ),
    .D(_00763_));
 sky130_as_sc_hs__dfxtp_2 _52658_ (.CLK(clknet_leaf_56_wb_clk_i),
    .Q(\tholin_riscv.regs[22][5] ),
    .D(_00764_));
 sky130_as_sc_hs__dfxtp_2 _52659_ (.CLK(clknet_leaf_57_wb_clk_i),
    .Q(\tholin_riscv.regs[22][6] ),
    .D(_00765_));
 sky130_as_sc_hs__dfxtp_2 _52660_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[22][7] ),
    .D(_00766_));
 sky130_as_sc_hs__dfxtp_2 _52661_ (.CLK(clknet_leaf_85_wb_clk_i),
    .Q(\tholin_riscv.regs[22][8] ),
    .D(_00767_));
 sky130_as_sc_hs__dfxtp_2 _52662_ (.CLK(clknet_leaf_42_wb_clk_i),
    .Q(\tholin_riscv.regs[22][9] ),
    .D(_00768_));
 sky130_as_sc_hs__dfxtp_2 _52663_ (.CLK(clknet_leaf_31_wb_clk_i),
    .Q(\tholin_riscv.regs[22][10] ),
    .D(_00769_));
 sky130_as_sc_hs__dfxtp_2 _52664_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[22][11] ),
    .D(_00770_));
 sky130_as_sc_hs__dfxtp_2 _52665_ (.CLK(clknet_leaf_28_wb_clk_i),
    .Q(\tholin_riscv.regs[22][12] ),
    .D(_00771_));
 sky130_as_sc_hs__dfxtp_2 _52666_ (.CLK(clknet_leaf_21_wb_clk_i),
    .Q(\tholin_riscv.regs[22][13] ),
    .D(_00772_));
 sky130_as_sc_hs__dfxtp_2 _52667_ (.CLK(clknet_leaf_17_wb_clk_i),
    .Q(\tholin_riscv.regs[22][14] ),
    .D(_00773_));
 sky130_as_sc_hs__dfxtp_2 _52668_ (.CLK(clknet_leaf_16_wb_clk_i),
    .Q(\tholin_riscv.regs[22][15] ),
    .D(_00774_));
 sky130_as_sc_hs__dfxtp_2 _52669_ (.CLK(clknet_leaf_75_wb_clk_i),
    .Q(\tholin_riscv.regs[22][16] ),
    .D(_00775_));
 sky130_as_sc_hs__dfxtp_2 _52670_ (.CLK(clknet_leaf_78_wb_clk_i),
    .Q(\tholin_riscv.regs[22][17] ),
    .D(_00776_));
 sky130_as_sc_hs__dfxtp_2 _52671_ (.CLK(clknet_leaf_123_wb_clk_i),
    .Q(\tholin_riscv.regs[22][18] ),
    .D(_00777_));
 sky130_as_sc_hs__dfxtp_2 _52672_ (.CLK(clknet_leaf_75_wb_clk_i),
    .Q(\tholin_riscv.regs[22][19] ),
    .D(_00778_));
 sky130_as_sc_hs__dfxtp_2 _52673_ (.CLK(clknet_leaf_72_wb_clk_i),
    .Q(\tholin_riscv.regs[22][20] ),
    .D(_00779_));
 sky130_as_sc_hs__dfxtp_2 _52674_ (.CLK(clknet_leaf_80_wb_clk_i),
    .Q(\tholin_riscv.regs[22][21] ),
    .D(_00780_));
 sky130_as_sc_hs__dfxtp_2 _52675_ (.CLK(clknet_leaf_127_wb_clk_i),
    .Q(\tholin_riscv.regs[22][22] ),
    .D(_00781_));
 sky130_as_sc_hs__dfxtp_2 _52676_ (.CLK(clknet_leaf_66_wb_clk_i),
    .Q(\tholin_riscv.regs[22][23] ),
    .D(_00782_));
 sky130_as_sc_hs__dfxtp_2 _52677_ (.CLK(clknet_leaf_42_wb_clk_i),
    .Q(\tholin_riscv.regs[22][24] ),
    .D(_00783_));
 sky130_as_sc_hs__dfxtp_2 _52678_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[22][25] ),
    .D(_00784_));
 sky130_as_sc_hs__dfxtp_2 _52679_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[22][26] ),
    .D(_00785_));
 sky130_as_sc_hs__dfxtp_2 _52680_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[22][27] ),
    .D(_00786_));
 sky130_as_sc_hs__dfxtp_2 _52681_ (.CLK(clknet_leaf_89_wb_clk_i),
    .Q(\tholin_riscv.regs[22][28] ),
    .D(_00787_));
 sky130_as_sc_hs__dfxtp_2 _52682_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[22][29] ),
    .D(_00788_));
 sky130_as_sc_hs__dfxtp_2 _52683_ (.CLK(clknet_leaf_152_wb_clk_i),
    .Q(\tholin_riscv.regs[22][30] ),
    .D(_00789_));
 sky130_as_sc_hs__dfxtp_2 _52684_ (.CLK(clknet_leaf_113_wb_clk_i),
    .Q(\tholin_riscv.regs[22][31] ),
    .D(_00790_));
 sky130_as_sc_hs__dfxtp_2 _52685_ (.CLK(clknet_leaf_196_wb_clk_i),
    .Q(\tholin_riscv.regs[21][0] ),
    .D(net674));
 sky130_as_sc_hs__dfxtp_2 _52686_ (.CLK(clknet_leaf_127_wb_clk_i),
    .Q(\tholin_riscv.regs[21][1] ),
    .D(_00792_));
 sky130_as_sc_hs__dfxtp_2 _52687_ (.CLK(clknet_leaf_6_wb_clk_i),
    .Q(\tholin_riscv.regs[21][2] ),
    .D(_00793_));
 sky130_as_sc_hs__dfxtp_2 _52688_ (.CLK(clknet_leaf_9_wb_clk_i),
    .Q(\tholin_riscv.regs[21][3] ),
    .D(_00794_));
 sky130_as_sc_hs__dfxtp_2 _52689_ (.CLK(clknet_leaf_149_wb_clk_i),
    .Q(\tholin_riscv.regs[21][4] ),
    .D(_00795_));
 sky130_as_sc_hs__dfxtp_2 _52690_ (.CLK(clknet_leaf_56_wb_clk_i),
    .Q(\tholin_riscv.regs[21][5] ),
    .D(_00796_));
 sky130_as_sc_hs__dfxtp_2 _52691_ (.CLK(clknet_leaf_59_wb_clk_i),
    .Q(\tholin_riscv.regs[21][6] ),
    .D(_00797_));
 sky130_as_sc_hs__dfxtp_2 _52692_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[21][7] ),
    .D(_00798_));
 sky130_as_sc_hs__dfxtp_2 _52693_ (.CLK(clknet_leaf_80_wb_clk_i),
    .Q(\tholin_riscv.regs[21][8] ),
    .D(_00799_));
 sky130_as_sc_hs__dfxtp_2 _52694_ (.CLK(clknet_leaf_41_wb_clk_i),
    .Q(\tholin_riscv.regs[21][9] ),
    .D(_00800_));
 sky130_as_sc_hs__dfxtp_2 _52695_ (.CLK(clknet_leaf_49_wb_clk_i),
    .Q(\tholin_riscv.regs[21][10] ),
    .D(_00801_));
 sky130_as_sc_hs__dfxtp_2 _52696_ (.CLK(clknet_leaf_29_wb_clk_i),
    .Q(\tholin_riscv.regs[21][11] ),
    .D(_00802_));
 sky130_as_sc_hs__dfxtp_2 _52697_ (.CLK(clknet_leaf_27_wb_clk_i),
    .Q(\tholin_riscv.regs[21][12] ),
    .D(_00803_));
 sky130_as_sc_hs__dfxtp_2 _52698_ (.CLK(clknet_leaf_21_wb_clk_i),
    .Q(\tholin_riscv.regs[21][13] ),
    .D(_00804_));
 sky130_as_sc_hs__dfxtp_2 _52699_ (.CLK(clknet_leaf_18_wb_clk_i),
    .Q(\tholin_riscv.regs[21][14] ),
    .D(_00805_));
 sky130_as_sc_hs__dfxtp_2 _52700_ (.CLK(clknet_leaf_16_wb_clk_i),
    .Q(\tholin_riscv.regs[21][15] ),
    .D(_00806_));
 sky130_as_sc_hs__dfxtp_2 _52701_ (.CLK(clknet_leaf_100_wb_clk_i),
    .Q(\tholin_riscv.regs[21][16] ),
    .D(_00807_));
 sky130_as_sc_hs__dfxtp_2 _52702_ (.CLK(clknet_leaf_118_wb_clk_i),
    .Q(\tholin_riscv.regs[21][17] ),
    .D(_00808_));
 sky130_as_sc_hs__dfxtp_2 _52703_ (.CLK(clknet_leaf_146_wb_clk_i),
    .Q(\tholin_riscv.regs[21][18] ),
    .D(_00809_));
 sky130_as_sc_hs__dfxtp_2 _52704_ (.CLK(clknet_leaf_111_wb_clk_i),
    .Q(\tholin_riscv.regs[21][19] ),
    .D(_00810_));
 sky130_as_sc_hs__dfxtp_2 _52705_ (.CLK(clknet_leaf_101_wb_clk_i),
    .Q(\tholin_riscv.regs[21][20] ),
    .D(_00811_));
 sky130_as_sc_hs__dfxtp_2 _52706_ (.CLK(clknet_leaf_111_wb_clk_i),
    .Q(\tholin_riscv.regs[21][21] ),
    .D(_00812_));
 sky130_as_sc_hs__dfxtp_2 _52707_ (.CLK(clknet_leaf_116_wb_clk_i),
    .Q(\tholin_riscv.regs[21][22] ),
    .D(_00813_));
 sky130_as_sc_hs__dfxtp_2 _52708_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.regs[21][23] ),
    .D(_00814_));
 sky130_as_sc_hs__dfxtp_2 _52709_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[21][24] ),
    .D(_00815_));
 sky130_as_sc_hs__dfxtp_2 _52710_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[21][25] ),
    .D(_00816_));
 sky130_as_sc_hs__dfxtp_2 _52711_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[21][26] ),
    .D(_00817_));
 sky130_as_sc_hs__dfxtp_2 _52712_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[21][27] ),
    .D(_00818_));
 sky130_as_sc_hs__dfxtp_2 _52713_ (.CLK(clknet_leaf_89_wb_clk_i),
    .Q(\tholin_riscv.regs[21][28] ),
    .D(_00819_));
 sky130_as_sc_hs__dfxtp_2 _52714_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[21][29] ),
    .D(_00820_));
 sky130_as_sc_hs__dfxtp_2 _52715_ (.CLK(clknet_leaf_150_wb_clk_i),
    .Q(\tholin_riscv.regs[21][30] ),
    .D(_00821_));
 sky130_as_sc_hs__dfxtp_2 _52716_ (.CLK(clknet_leaf_157_wb_clk_i),
    .Q(\tholin_riscv.regs[21][31] ),
    .D(_00822_));
 sky130_as_sc_hs__dfxtp_2 _52717_ (.CLK(clknet_leaf_135_wb_clk_i),
    .Q(\tholin_riscv.regs[5][0] ),
    .D(net722));
 sky130_as_sc_hs__dfxtp_2 _52718_ (.CLK(clknet_leaf_68_wb_clk_i),
    .Q(\tholin_riscv.regs[5][1] ),
    .D(_00824_));
 sky130_as_sc_hs__dfxtp_2 _52719_ (.CLK(clknet_leaf_65_wb_clk_i),
    .Q(\tholin_riscv.regs[5][2] ),
    .D(_00825_));
 sky130_as_sc_hs__dfxtp_2 _52720_ (.CLK(clknet_leaf_55_wb_clk_i),
    .Q(\tholin_riscv.regs[5][3] ),
    .D(_00826_));
 sky130_as_sc_hs__dfxtp_2 _52721_ (.CLK(clknet_leaf_107_wb_clk_i),
    .Q(\tholin_riscv.regs[5][4] ),
    .D(_00827_));
 sky130_as_sc_hs__dfxtp_2 _52722_ (.CLK(clknet_leaf_58_wb_clk_i),
    .Q(\tholin_riscv.regs[5][5] ),
    .D(_00828_));
 sky130_as_sc_hs__dfxtp_2 _52723_ (.CLK(clknet_leaf_59_wb_clk_i),
    .Q(\tholin_riscv.regs[5][6] ),
    .D(_00829_));
 sky130_as_sc_hs__dfxtp_2 _52724_ (.CLK(clknet_leaf_50_wb_clk_i),
    .Q(\tholin_riscv.regs[5][7] ),
    .D(_00830_));
 sky130_as_sc_hs__dfxtp_2 _52725_ (.CLK(clknet_leaf_84_wb_clk_i),
    .Q(\tholin_riscv.regs[5][8] ),
    .D(_00831_));
 sky130_as_sc_hs__dfxtp_2 _52726_ (.CLK(clknet_leaf_46_wb_clk_i),
    .Q(\tholin_riscv.regs[5][9] ),
    .D(_00832_));
 sky130_as_sc_hs__dfxtp_2 _52727_ (.CLK(clknet_leaf_46_wb_clk_i),
    .Q(\tholin_riscv.regs[5][10] ),
    .D(_00833_));
 sky130_as_sc_hs__dfxtp_2 _52728_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[5][11] ),
    .D(_00834_));
 sky130_as_sc_hs__dfxtp_2 _52729_ (.CLK(clknet_leaf_37_wb_clk_i),
    .Q(\tholin_riscv.regs[5][12] ),
    .D(_00835_));
 sky130_as_sc_hs__dfxtp_2 _52730_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[5][13] ),
    .D(_00836_));
 sky130_as_sc_hs__dfxtp_2 _52731_ (.CLK(clknet_leaf_12_wb_clk_i),
    .Q(\tholin_riscv.regs[5][14] ),
    .D(_00837_));
 sky130_as_sc_hs__dfxtp_2 _52732_ (.CLK(clknet_leaf_53_wb_clk_i),
    .Q(\tholin_riscv.regs[5][15] ),
    .D(_00838_));
 sky130_as_sc_hs__dfxtp_2 _52733_ (.CLK(clknet_leaf_103_wb_clk_i),
    .Q(\tholin_riscv.regs[5][16] ),
    .D(_00839_));
 sky130_as_sc_hs__dfxtp_2 _52734_ (.CLK(clknet_leaf_107_wb_clk_i),
    .Q(\tholin_riscv.regs[5][17] ),
    .D(_00840_));
 sky130_as_sc_hs__dfxtp_2 _52735_ (.CLK(clknet_leaf_94_wb_clk_i),
    .Q(\tholin_riscv.regs[5][18] ),
    .D(_00841_));
 sky130_as_sc_hs__dfxtp_2 _52736_ (.CLK(clknet_leaf_103_wb_clk_i),
    .Q(\tholin_riscv.regs[5][19] ),
    .D(_00842_));
 sky130_as_sc_hs__dfxtp_2 _52737_ (.CLK(clknet_leaf_103_wb_clk_i),
    .Q(\tholin_riscv.regs[5][20] ),
    .D(_00843_));
 sky130_as_sc_hs__dfxtp_2 _52738_ (.CLK(clknet_leaf_109_wb_clk_i),
    .Q(\tholin_riscv.regs[5][21] ),
    .D(_00844_));
 sky130_as_sc_hs__dfxtp_2 _52739_ (.CLK(clknet_leaf_113_wb_clk_i),
    .Q(\tholin_riscv.regs[5][22] ),
    .D(_00845_));
 sky130_as_sc_hs__dfxtp_2 _52740_ (.CLK(clknet_leaf_93_wb_clk_i),
    .Q(\tholin_riscv.regs[5][23] ),
    .D(_00846_));
 sky130_as_sc_hs__dfxtp_2 _52741_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[5][24] ),
    .D(_00847_));
 sky130_as_sc_hs__dfxtp_2 _52742_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[5][25] ),
    .D(_00848_));
 sky130_as_sc_hs__dfxtp_2 _52743_ (.CLK(clknet_leaf_33_wb_clk_i),
    .Q(\tholin_riscv.regs[5][26] ),
    .D(_00849_));
 sky130_as_sc_hs__dfxtp_2 _52744_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[5][27] ),
    .D(_00850_));
 sky130_as_sc_hs__dfxtp_2 _52745_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[5][28] ),
    .D(_00851_));
 sky130_as_sc_hs__dfxtp_2 _52746_ (.CLK(clknet_leaf_36_wb_clk_i),
    .Q(\tholin_riscv.regs[5][29] ),
    .D(_00852_));
 sky130_as_sc_hs__dfxtp_2 _52747_ (.CLK(clknet_leaf_135_wb_clk_i),
    .Q(\tholin_riscv.regs[5][30] ),
    .D(_00853_));
 sky130_as_sc_hs__dfxtp_2 _52748_ (.CLK(clknet_leaf_93_wb_clk_i),
    .Q(\tholin_riscv.regs[5][31] ),
    .D(_00854_));
 sky130_as_sc_hs__dfxtp_2 _52749_ (.CLK(clknet_leaf_65_wb_clk_i),
    .Q(\tholin_riscv.regs[19][0] ),
    .D(net728));
 sky130_as_sc_hs__dfxtp_2 _52750_ (.CLK(clknet_leaf_127_wb_clk_i),
    .Q(\tholin_riscv.regs[19][1] ),
    .D(_00856_));
 sky130_as_sc_hs__dfxtp_2 _52751_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[19][2] ),
    .D(_00857_));
 sky130_as_sc_hs__dfxtp_2 _52752_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[19][3] ),
    .D(_00858_));
 sky130_as_sc_hs__dfxtp_2 _52753_ (.CLK(clknet_leaf_149_wb_clk_i),
    .Q(\tholin_riscv.regs[19][4] ),
    .D(_00859_));
 sky130_as_sc_hs__dfxtp_2 _52754_ (.CLK(clknet_leaf_58_wb_clk_i),
    .Q(\tholin_riscv.regs[19][5] ),
    .D(_00860_));
 sky130_as_sc_hs__dfxtp_2 _52755_ (.CLK(clknet_leaf_56_wb_clk_i),
    .Q(\tholin_riscv.regs[19][6] ),
    .D(_00861_));
 sky130_as_sc_hs__dfxtp_2 _52756_ (.CLK(clknet_leaf_53_wb_clk_i),
    .Q(\tholin_riscv.regs[19][7] ),
    .D(_00862_));
 sky130_as_sc_hs__dfxtp_2 _52757_ (.CLK(clknet_leaf_85_wb_clk_i),
    .Q(\tholin_riscv.regs[19][8] ),
    .D(_00863_));
 sky130_as_sc_hs__dfxtp_2 _52758_ (.CLK(clknet_leaf_38_wb_clk_i),
    .Q(\tholin_riscv.regs[19][9] ),
    .D(_00864_));
 sky130_as_sc_hs__dfxtp_2 _52759_ (.CLK(clknet_leaf_31_wb_clk_i),
    .Q(\tholin_riscv.regs[19][10] ),
    .D(_00865_));
 sky130_as_sc_hs__dfxtp_2 _52760_ (.CLK(clknet_leaf_29_wb_clk_i),
    .Q(\tholin_riscv.regs[19][11] ),
    .D(_00866_));
 sky130_as_sc_hs__dfxtp_2 _52761_ (.CLK(clknet_leaf_27_wb_clk_i),
    .Q(\tholin_riscv.regs[19][12] ),
    .D(_00867_));
 sky130_as_sc_hs__dfxtp_2 _52762_ (.CLK(clknet_leaf_22_wb_clk_i),
    .Q(\tholin_riscv.regs[19][13] ),
    .D(_00868_));
 sky130_as_sc_hs__dfxtp_2 _52763_ (.CLK(clknet_leaf_19_wb_clk_i),
    .Q(\tholin_riscv.regs[19][14] ),
    .D(_00869_));
 sky130_as_sc_hs__dfxtp_2 _52764_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[19][15] ),
    .D(_00870_));
 sky130_as_sc_hs__dfxtp_2 _52765_ (.CLK(clknet_leaf_106_wb_clk_i),
    .Q(\tholin_riscv.regs[19][16] ),
    .D(_00871_));
 sky130_as_sc_hs__dfxtp_2 _52766_ (.CLK(clknet_leaf_110_wb_clk_i),
    .Q(\tholin_riscv.regs[19][17] ),
    .D(_00872_));
 sky130_as_sc_hs__dfxtp_2 _52767_ (.CLK(clknet_leaf_109_wb_clk_i),
    .Q(\tholin_riscv.regs[19][18] ),
    .D(_00873_));
 sky130_as_sc_hs__dfxtp_2 _52768_ (.CLK(clknet_leaf_151_wb_clk_i),
    .Q(\tholin_riscv.regs[19][19] ),
    .D(_00874_));
 sky130_as_sc_hs__dfxtp_2 _52769_ (.CLK(clknet_leaf_104_wb_clk_i),
    .Q(\tholin_riscv.regs[19][20] ),
    .D(_00875_));
 sky130_as_sc_hs__dfxtp_2 _52770_ (.CLK(clknet_leaf_105_wb_clk_i),
    .Q(\tholin_riscv.regs[19][21] ),
    .D(_00876_));
 sky130_as_sc_hs__dfxtp_2 _52771_ (.CLK(clknet_leaf_114_wb_clk_i),
    .Q(\tholin_riscv.regs[19][22] ),
    .D(_00877_));
 sky130_as_sc_hs__dfxtp_2 _52772_ (.CLK(clknet_leaf_106_wb_clk_i),
    .Q(\tholin_riscv.regs[19][23] ),
    .D(_00878_));
 sky130_as_sc_hs__dfxtp_2 _52773_ (.CLK(clknet_leaf_42_wb_clk_i),
    .Q(\tholin_riscv.regs[19][24] ),
    .D(_00879_));
 sky130_as_sc_hs__dfxtp_2 _52774_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[19][25] ),
    .D(_00880_));
 sky130_as_sc_hs__dfxtp_2 _52775_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[19][26] ),
    .D(_00881_));
 sky130_as_sc_hs__dfxtp_2 _52776_ (.CLK(clknet_leaf_90_wb_clk_i),
    .Q(\tholin_riscv.regs[19][27] ),
    .D(_00882_));
 sky130_as_sc_hs__dfxtp_2 _52777_ (.CLK(clknet_leaf_88_wb_clk_i),
    .Q(\tholin_riscv.regs[19][28] ),
    .D(_00883_));
 sky130_as_sc_hs__dfxtp_2 _52778_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[19][29] ),
    .D(_00884_));
 sky130_as_sc_hs__dfxtp_2 _52779_ (.CLK(clknet_leaf_104_wb_clk_i),
    .Q(\tholin_riscv.regs[19][30] ),
    .D(_00885_));
 sky130_as_sc_hs__dfxtp_2 _52780_ (.CLK(clknet_leaf_152_wb_clk_i),
    .Q(\tholin_riscv.regs[19][31] ),
    .D(_00886_));
 sky130_as_sc_hs__dfxtp_2 _52781_ (.CLK(clknet_leaf_133_wb_clk_i),
    .Q(\tholin_riscv.regs[4][0] ),
    .D(net746));
 sky130_as_sc_hs__dfxtp_2 _52782_ (.CLK(clknet_leaf_68_wb_clk_i),
    .Q(\tholin_riscv.regs[4][1] ),
    .D(_00888_));
 sky130_as_sc_hs__dfxtp_2 _52783_ (.CLK(clknet_leaf_65_wb_clk_i),
    .Q(\tholin_riscv.regs[4][2] ),
    .D(_00889_));
 sky130_as_sc_hs__dfxtp_2 _52784_ (.CLK(clknet_leaf_55_wb_clk_i),
    .Q(\tholin_riscv.regs[4][3] ),
    .D(_00890_));
 sky130_as_sc_hs__dfxtp_2 _52785_ (.CLK(clknet_leaf_70_wb_clk_i),
    .Q(\tholin_riscv.regs[4][4] ),
    .D(_00891_));
 sky130_as_sc_hs__dfxtp_2 _52786_ (.CLK(clknet_leaf_47_wb_clk_i),
    .Q(\tholin_riscv.regs[4][5] ),
    .D(_00892_));
 sky130_as_sc_hs__dfxtp_2 _52787_ (.CLK(clknet_leaf_59_wb_clk_i),
    .Q(\tholin_riscv.regs[4][6] ),
    .D(_00893_));
 sky130_as_sc_hs__dfxtp_2 _52788_ (.CLK(clknet_leaf_50_wb_clk_i),
    .Q(\tholin_riscv.regs[4][7] ),
    .D(_00894_));
 sky130_as_sc_hs__dfxtp_2 _52789_ (.CLK(clknet_leaf_84_wb_clk_i),
    .Q(\tholin_riscv.regs[4][8] ),
    .D(_00895_));
 sky130_as_sc_hs__dfxtp_2 _52790_ (.CLK(clknet_leaf_46_wb_clk_i),
    .Q(\tholin_riscv.regs[4][9] ),
    .D(_00896_));
 sky130_as_sc_hs__dfxtp_2 _52791_ (.CLK(clknet_leaf_48_wb_clk_i),
    .Q(\tholin_riscv.regs[4][10] ),
    .D(_00897_));
 sky130_as_sc_hs__dfxtp_2 _52792_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[4][11] ),
    .D(_00898_));
 sky130_as_sc_hs__dfxtp_2 _52793_ (.CLK(clknet_leaf_37_wb_clk_i),
    .Q(\tholin_riscv.regs[4][12] ),
    .D(_00899_));
 sky130_as_sc_hs__dfxtp_2 _52794_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[4][13] ),
    .D(_00900_));
 sky130_as_sc_hs__dfxtp_2 _52795_ (.CLK(clknet_leaf_12_wb_clk_i),
    .Q(\tholin_riscv.regs[4][14] ),
    .D(_00901_));
 sky130_as_sc_hs__dfxtp_2 _52796_ (.CLK(clknet_leaf_15_wb_clk_i),
    .Q(\tholin_riscv.regs[4][15] ),
    .D(_00902_));
 sky130_as_sc_hs__dfxtp_2 _52797_ (.CLK(clknet_leaf_85_wb_clk_i),
    .Q(\tholin_riscv.regs[4][16] ),
    .D(_00903_));
 sky130_as_sc_hs__dfxtp_2 _52798_ (.CLK(clknet_leaf_41_wb_clk_i),
    .Q(\tholin_riscv.regs[4][17] ),
    .D(_00904_));
 sky130_as_sc_hs__dfxtp_2 _52799_ (.CLK(clknet_leaf_82_wb_clk_i),
    .Q(\tholin_riscv.regs[4][18] ),
    .D(_00905_));
 sky130_as_sc_hs__dfxtp_2 _52800_ (.CLK(clknet_leaf_46_wb_clk_i),
    .Q(\tholin_riscv.regs[4][19] ),
    .D(_00906_));
 sky130_as_sc_hs__dfxtp_2 _52801_ (.CLK(clknet_leaf_73_wb_clk_i),
    .Q(\tholin_riscv.regs[4][20] ),
    .D(_00907_));
 sky130_as_sc_hs__dfxtp_2 _52802_ (.CLK(clknet_leaf_86_wb_clk_i),
    .Q(\tholin_riscv.regs[4][21] ),
    .D(_00908_));
 sky130_as_sc_hs__dfxtp_2 _52803_ (.CLK(clknet_leaf_81_wb_clk_i),
    .Q(\tholin_riscv.regs[4][22] ),
    .D(_00909_));
 sky130_as_sc_hs__dfxtp_2 _52804_ (.CLK(clknet_leaf_67_wb_clk_i),
    .Q(\tholin_riscv.regs[4][23] ),
    .D(_00910_));
 sky130_as_sc_hs__dfxtp_2 _52805_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[4][24] ),
    .D(_00911_));
 sky130_as_sc_hs__dfxtp_2 _52806_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[4][25] ),
    .D(_00912_));
 sky130_as_sc_hs__dfxtp_2 _52807_ (.CLK(clknet_leaf_33_wb_clk_i),
    .Q(\tholin_riscv.regs[4][26] ),
    .D(_00913_));
 sky130_as_sc_hs__dfxtp_2 _52808_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[4][27] ),
    .D(_00914_));
 sky130_as_sc_hs__dfxtp_2 _52809_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[4][28] ),
    .D(_00915_));
 sky130_as_sc_hs__dfxtp_2 _52810_ (.CLK(clknet_leaf_38_wb_clk_i),
    .Q(\tholin_riscv.regs[4][29] ),
    .D(_00916_));
 sky130_as_sc_hs__dfxtp_2 _52811_ (.CLK(clknet_leaf_153_wb_clk_i),
    .Q(\tholin_riscv.regs[4][30] ),
    .D(_00917_));
 sky130_as_sc_hs__dfxtp_2 _52812_ (.CLK(clknet_leaf_158_wb_clk_i),
    .Q(\tholin_riscv.regs[4][31] ),
    .D(_00918_));
 sky130_as_sc_hs__dfxtp_2 _52813_ (.CLK(clknet_leaf_129_wb_clk_i),
    .Q(\tholin_riscv.regs[3][0] ),
    .D(net677));
 sky130_as_sc_hs__dfxtp_2 _52814_ (.CLK(clknet_leaf_68_wb_clk_i),
    .Q(\tholin_riscv.regs[3][1] ),
    .D(_00920_));
 sky130_as_sc_hs__dfxtp_2 _52815_ (.CLK(clknet_leaf_65_wb_clk_i),
    .Q(\tholin_riscv.regs[3][2] ),
    .D(_00921_));
 sky130_as_sc_hs__dfxtp_2 _52816_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[3][3] ),
    .D(_00922_));
 sky130_as_sc_hs__dfxtp_2 _52817_ (.CLK(clknet_leaf_107_wb_clk_i),
    .Q(\tholin_riscv.regs[3][4] ),
    .D(_00923_));
 sky130_as_sc_hs__dfxtp_2 _52818_ (.CLK(clknet_leaf_57_wb_clk_i),
    .Q(\tholin_riscv.regs[3][5] ),
    .D(_00924_));
 sky130_as_sc_hs__dfxtp_2 _52819_ (.CLK(clknet_leaf_60_wb_clk_i),
    .Q(\tholin_riscv.regs[3][6] ),
    .D(_00925_));
 sky130_as_sc_hs__dfxtp_2 _52820_ (.CLK(clknet_leaf_51_wb_clk_i),
    .Q(\tholin_riscv.regs[3][7] ),
    .D(_00926_));
 sky130_as_sc_hs__dfxtp_2 _52821_ (.CLK(clknet_leaf_83_wb_clk_i),
    .Q(\tholin_riscv.regs[3][8] ),
    .D(_00927_));
 sky130_as_sc_hs__dfxtp_2 _52822_ (.CLK(clknet_leaf_44_wb_clk_i),
    .Q(\tholin_riscv.regs[3][9] ),
    .D(_00928_));
 sky130_as_sc_hs__dfxtp_2 _52823_ (.CLK(clknet_leaf_48_wb_clk_i),
    .Q(\tholin_riscv.regs[3][10] ),
    .D(_00929_));
 sky130_as_sc_hs__dfxtp_2 _52824_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[3][11] ),
    .D(_00930_));
 sky130_as_sc_hs__dfxtp_2 _52825_ (.CLK(clknet_leaf_32_wb_clk_i),
    .Q(\tholin_riscv.regs[3][12] ),
    .D(_00931_));
 sky130_as_sc_hs__dfxtp_2 _52826_ (.CLK(clknet_leaf_33_wb_clk_i),
    .Q(\tholin_riscv.regs[3][13] ),
    .D(_00932_));
 sky130_as_sc_hs__dfxtp_2 _52827_ (.CLK(clknet_leaf_12_wb_clk_i),
    .Q(\tholin_riscv.regs[3][14] ),
    .D(_00933_));
 sky130_as_sc_hs__dfxtp_2 _52828_ (.CLK(clknet_leaf_15_wb_clk_i),
    .Q(\tholin_riscv.regs[3][15] ),
    .D(_00934_));
 sky130_as_sc_hs__dfxtp_2 _52829_ (.CLK(clknet_leaf_114_wb_clk_i),
    .Q(\tholin_riscv.regs[3][16] ),
    .D(_00935_));
 sky130_as_sc_hs__dfxtp_2 _52830_ (.CLK(clknet_leaf_107_wb_clk_i),
    .Q(\tholin_riscv.regs[3][17] ),
    .D(_00936_));
 sky130_as_sc_hs__dfxtp_2 _52831_ (.CLK(clknet_leaf_100_wb_clk_i),
    .Q(\tholin_riscv.regs[3][18] ),
    .D(_00937_));
 sky130_as_sc_hs__dfxtp_2 _52832_ (.CLK(clknet_leaf_108_wb_clk_i),
    .Q(\tholin_riscv.regs[3][19] ),
    .D(_00938_));
 sky130_as_sc_hs__dfxtp_2 _52833_ (.CLK(clknet_leaf_102_wb_clk_i),
    .Q(\tholin_riscv.regs[3][20] ),
    .D(_00939_));
 sky130_as_sc_hs__dfxtp_2 _52834_ (.CLK(clknet_leaf_108_wb_clk_i),
    .Q(\tholin_riscv.regs[3][21] ),
    .D(_00940_));
 sky130_as_sc_hs__dfxtp_2 _52835_ (.CLK(clknet_leaf_104_wb_clk_i),
    .Q(\tholin_riscv.regs[3][22] ),
    .D(_00941_));
 sky130_as_sc_hs__dfxtp_2 _52836_ (.CLK(clknet_leaf_105_wb_clk_i),
    .Q(\tholin_riscv.regs[3][23] ),
    .D(_00942_));
 sky130_as_sc_hs__dfxtp_2 _52837_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[3][24] ),
    .D(_00943_));
 sky130_as_sc_hs__dfxtp_2 _52838_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[3][25] ),
    .D(_00944_));
 sky130_as_sc_hs__dfxtp_2 _52839_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[3][26] ),
    .D(_00945_));
 sky130_as_sc_hs__dfxtp_2 _52840_ (.CLK(clknet_leaf_25_wb_clk_i),
    .Q(\tholin_riscv.regs[3][27] ),
    .D(_00946_));
 sky130_as_sc_hs__dfxtp_2 _52841_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[3][28] ),
    .D(_00947_));
 sky130_as_sc_hs__dfxtp_2 _52842_ (.CLK(clknet_leaf_36_wb_clk_i),
    .Q(\tholin_riscv.regs[3][29] ),
    .D(_00948_));
 sky130_as_sc_hs__dfxtp_2 _52843_ (.CLK(clknet_leaf_104_wb_clk_i),
    .Q(\tholin_riscv.regs[3][30] ),
    .D(_00949_));
 sky130_as_sc_hs__dfxtp_2 _52844_ (.CLK(clknet_leaf_135_wb_clk_i),
    .Q(\tholin_riscv.regs[3][31] ),
    .D(_00950_));
 sky130_as_sc_hs__dfxtp_2 _52845_ (.CLK(clknet_leaf_137_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_counter[0] ),
    .D(_00951_));
 sky130_as_sc_hs__dfxtp_2 _52846_ (.CLK(clknet_leaf_137_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_counter[1] ),
    .D(_00952_));
 sky130_as_sc_hs__dfxtp_2 _52847_ (.CLK(clknet_leaf_116_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_counter[2] ),
    .D(_00953_));
 sky130_as_sc_hs__dfxtp_2 _52848_ (.CLK(clknet_leaf_116_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_counter[3] ),
    .D(_00954_));
 sky130_as_sc_hs__dfxtp_2 _52849_ (.CLK(clknet_leaf_141_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[0] ),
    .D(_00955_));
 sky130_as_sc_hs__dfxtp_2 _52850_ (.CLK(clknet_leaf_141_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[1] ),
    .D(_00956_));
 sky130_as_sc_hs__dfxtp_2 _52851_ (.CLK(clknet_leaf_138_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[2] ),
    .D(_00957_));
 sky130_as_sc_hs__dfxtp_2 _52852_ (.CLK(clknet_leaf_147_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[3] ),
    .D(_00958_));
 sky130_as_sc_hs__dfxtp_2 _52853_ (.CLK(clknet_leaf_138_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[4] ),
    .D(_00959_));
 sky130_as_sc_hs__dfxtp_2 _52854_ (.CLK(clknet_leaf_138_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[5] ),
    .D(_00960_));
 sky130_as_sc_hs__dfxtp_2 _52855_ (.CLK(clknet_leaf_138_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[6] ),
    .D(_00961_));
 sky130_as_sc_hs__dfxtp_2 _52856_ (.CLK(clknet_leaf_138_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[7] ),
    .D(_00962_));
 sky130_as_sc_hs__dfxtp_2 _52857_ (.CLK(clknet_leaf_138_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[8] ),
    .D(_00963_));
 sky130_as_sc_hs__dfxtp_2 _52858_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[9] ),
    .D(_00964_));
 sky130_as_sc_hs__dfxtp_2 _52859_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[10] ),
    .D(_00965_));
 sky130_as_sc_hs__dfxtp_2 _52860_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[11] ),
    .D(_00966_));
 sky130_as_sc_hs__dfxtp_2 _52861_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[12] ),
    .D(_00967_));
 sky130_as_sc_hs__dfxtp_2 _52862_ (.CLK(clknet_leaf_138_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[13] ),
    .D(_00968_));
 sky130_as_sc_hs__dfxtp_2 _52863_ (.CLK(clknet_leaf_138_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[14] ),
    .D(_00969_));
 sky130_as_sc_hs__dfxtp_2 _52864_ (.CLK(clknet_leaf_140_wb_clk_i),
    .Q(\tholin_riscv.uart.div_counter[15] ),
    .D(_00970_));
 sky130_as_sc_hs__dfxtp_2 _52865_ (.CLK(clknet_leaf_124_wb_clk_i),
    .Q(\tholin_riscv.uart.dout[0] ),
    .D(net607));
 sky130_as_sc_hs__dfxtp_2 _52866_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.uart.dout[1] ),
    .D(net595));
 sky130_as_sc_hs__dfxtp_2 _52867_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.uart.dout[2] ),
    .D(net589));
 sky130_as_sc_hs__dfxtp_2 _52868_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.uart.dout[3] ),
    .D(net577));
 sky130_as_sc_hs__dfxtp_2 _52869_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.uart.dout[4] ),
    .D(net1726));
 sky130_as_sc_hs__dfxtp_2 _52870_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.uart.dout[5] ),
    .D(net592));
 sky130_as_sc_hs__dfxtp_2 _52871_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.uart.dout[6] ),
    .D(net586));
 sky130_as_sc_hs__dfxtp_2 _52872_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.uart.dout[7] ),
    .D(net568));
 sky130_as_sc_hs__dfxtp_2 _52873_ (.CLK(clknet_leaf_113_wb_clk_i),
    .Q(\tholin_riscv.spi.data_in_buff[0] ),
    .D(_00979_));
 sky130_as_sc_hs__dfxtp_2 _52874_ (.CLK(clknet_leaf_193_wb_clk_i),
    .Q(\tholin_riscv.spi.data_in_buff[1] ),
    .D(_00980_));
 sky130_as_sc_hs__dfxtp_2 _52875_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.spi.data_in_buff[2] ),
    .D(_00981_));
 sky130_as_sc_hs__dfxtp_2 _52876_ (.CLK(clknet_leaf_193_wb_clk_i),
    .Q(\tholin_riscv.spi.data_in_buff[3] ),
    .D(_00982_));
 sky130_as_sc_hs__dfxtp_2 _52877_ (.CLK(clknet_leaf_186_wb_clk_i),
    .Q(\tholin_riscv.spi.data_in_buff[4] ),
    .D(_00983_));
 sky130_as_sc_hs__dfxtp_2 _52878_ (.CLK(clknet_leaf_192_wb_clk_i),
    .Q(\tholin_riscv.spi.data_in_buff[5] ),
    .D(_00984_));
 sky130_as_sc_hs__dfxtp_2 _52879_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.spi.data_in_buff[6] ),
    .D(_00985_));
 sky130_as_sc_hs__dfxtp_2 _52880_ (.CLK(clknet_leaf_193_wb_clk_i),
    .Q(\tholin_riscv.spi.data_in_buff[7] ),
    .D(_00986_));
 sky130_as_sc_hs__dfxtp_2 _52881_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(net59),
    .D(_00987_));
 sky130_as_sc_hs__dfxtp_2 _52882_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(\tholin_riscv.uart.busy ),
    .D(_00988_));
 sky130_as_sc_hs__dfxtp_2 _52883_ (.CLK(clknet_leaf_188_wb_clk_i),
    .Q(\tholin_riscv.uart.has_byte ),
    .D(_00989_));
 sky130_as_sc_hs__dfxtp_2 _52884_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.uart.data_buff[0] ),
    .D(_00990_));
 sky130_as_sc_hs__dfxtp_2 _52885_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.uart.data_buff[1] ),
    .D(_00991_));
 sky130_as_sc_hs__dfxtp_2 _52886_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.uart.data_buff[2] ),
    .D(_00992_));
 sky130_as_sc_hs__dfxtp_2 _52887_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.uart.data_buff[3] ),
    .D(_00993_));
 sky130_as_sc_hs__dfxtp_2 _52888_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.uart.data_buff[4] ),
    .D(_00994_));
 sky130_as_sc_hs__dfxtp_2 _52889_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.uart.data_buff[5] ),
    .D(_00995_));
 sky130_as_sc_hs__dfxtp_2 _52890_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.uart.data_buff[6] ),
    .D(_00996_));
 sky130_as_sc_hs__dfxtp_2 _52891_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.uart.data_buff[7] ),
    .D(_00997_));
 sky130_as_sc_hs__dfxtp_2 _52892_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.uart.data_buff[8] ),
    .D(_00998_));
 sky130_as_sc_hs__dfxtp_2 _52893_ (.CLK(clknet_leaf_140_wb_clk_i),
    .Q(\tholin_riscv.uart.data_buff[9] ),
    .D(net583));
 sky130_as_sc_hs__dfxtp_2 _52894_ (.CLK(clknet_leaf_141_wb_clk_i),
    .Q(\tholin_riscv.uart.counter[0] ),
    .D(_01000_));
 sky130_as_sc_hs__dfxtp_2 _52895_ (.CLK(clknet_leaf_140_wb_clk_i),
    .Q(\tholin_riscv.uart.counter[1] ),
    .D(net756));
 sky130_as_sc_hs__dfxtp_2 _52896_ (.CLK(clknet_leaf_140_wb_clk_i),
    .Q(\tholin_riscv.uart.counter[2] ),
    .D(_01002_));
 sky130_as_sc_hs__dfxtp_2 _52897_ (.CLK(clknet_leaf_140_wb_clk_i),
    .Q(\tholin_riscv.uart.counter[3] ),
    .D(net623));
 sky130_as_sc_hs__dfxtp_2 _52898_ (.CLK(clknet_leaf_126_wb_clk_i),
    .Q(\tholin_riscv.uart.receiving ),
    .D(_01004_));
 sky130_as_sc_hs__dfxtp_2 _52899_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_buff[0] ),
    .D(_01005_));
 sky130_as_sc_hs__dfxtp_2 _52900_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_buff[1] ),
    .D(_01006_));
 sky130_as_sc_hs__dfxtp_2 _52901_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_buff[2] ),
    .D(_01007_));
 sky130_as_sc_hs__dfxtp_2 _52902_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_buff[3] ),
    .D(_01008_));
 sky130_as_sc_hs__dfxtp_2 _52903_ (.CLK(clknet_leaf_124_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_buff[4] ),
    .D(_01009_));
 sky130_as_sc_hs__dfxtp_2 _52904_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_buff[5] ),
    .D(_01010_));
 sky130_as_sc_hs__dfxtp_2 _52905_ (.CLK(clknet_leaf_125_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_buff[6] ),
    .D(_01011_));
 sky130_as_sc_hs__dfxtp_2 _52906_ (.CLK(clknet_leaf_126_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_buff[7] ),
    .D(net617));
 sky130_as_sc_hs__dfxtp_2 _52907_ (.CLK(clknet_leaf_137_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[0] ),
    .D(_01013_));
 sky130_as_sc_hs__dfxtp_2 _52908_ (.CLK(clknet_leaf_136_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[1] ),
    .D(_01014_));
 sky130_as_sc_hs__dfxtp_2 _52909_ (.CLK(clknet_leaf_136_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[2] ),
    .D(_01015_));
 sky130_as_sc_hs__dfxtp_2 _52910_ (.CLK(clknet_leaf_137_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[3] ),
    .D(_01016_));
 sky130_as_sc_hs__dfxtp_2 _52911_ (.CLK(clknet_leaf_137_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[4] ),
    .D(_01017_));
 sky130_as_sc_hs__dfxtp_2 _52912_ (.CLK(clknet_leaf_137_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[5] ),
    .D(_01018_));
 sky130_as_sc_hs__dfxtp_2 _52913_ (.CLK(clknet_leaf_138_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[6] ),
    .D(_01019_));
 sky130_as_sc_hs__dfxtp_2 _52914_ (.CLK(clknet_leaf_138_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[7] ),
    .D(_01020_));
 sky130_as_sc_hs__dfxtp_2 _52915_ (.CLK(clknet_leaf_138_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[8] ),
    .D(_01021_));
 sky130_as_sc_hs__dfxtp_2 _52916_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[9] ),
    .D(_01022_));
 sky130_as_sc_hs__dfxtp_2 _52917_ (.CLK(clknet_leaf_135_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[10] ),
    .D(_01023_));
 sky130_as_sc_hs__dfxtp_2 _52918_ (.CLK(clknet_leaf_135_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[11] ),
    .D(_01024_));
 sky130_as_sc_hs__dfxtp_2 _52919_ (.CLK(clknet_leaf_136_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[12] ),
    .D(_01025_));
 sky130_as_sc_hs__dfxtp_2 _52920_ (.CLK(clknet_leaf_136_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[13] ),
    .D(_01026_));
 sky130_as_sc_hs__dfxtp_2 _52921_ (.CLK(clknet_leaf_136_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[14] ),
    .D(_01027_));
 sky130_as_sc_hs__dfxtp_2 _52922_ (.CLK(clknet_leaf_136_wb_clk_i),
    .Q(\tholin_riscv.uart.receive_div_counter[15] ),
    .D(_01028_));
 sky130_as_sc_hs__dfxtp_2 _52923_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.spi.div_counter[0] ),
    .D(_01029_));
 sky130_as_sc_hs__dfxtp_2 _52924_ (.CLK(clknet_leaf_187_wb_clk_i),
    .Q(\tholin_riscv.spi.div_counter[1] ),
    .D(_01030_));
 sky130_as_sc_hs__dfxtp_2 _52925_ (.CLK(clknet_leaf_181_wb_clk_i),
    .Q(\tholin_riscv.spi.div_counter[2] ),
    .D(_01031_));
 sky130_as_sc_hs__dfxtp_2 _52926_ (.CLK(clknet_leaf_181_wb_clk_i),
    .Q(\tholin_riscv.spi.div_counter[3] ),
    .D(_01032_));
 sky130_as_sc_hs__dfxtp_2 _52927_ (.CLK(clknet_leaf_188_wb_clk_i),
    .Q(\tholin_riscv.spi.div_counter[4] ),
    .D(_01033_));
 sky130_as_sc_hs__dfxtp_2 _52928_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.spi.div_counter[5] ),
    .D(_01034_));
 sky130_as_sc_hs__dfxtp_2 _52929_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.spi.div_counter[6] ),
    .D(_01035_));
 sky130_as_sc_hs__dfxtp_2 _52930_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.spi.div_counter[7] ),
    .D(_01036_));
 sky130_as_sc_hs__dfxtp_2 _52931_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.spi.dout[0] ),
    .D(_01037_));
 sky130_as_sc_hs__dfxtp_2 _52932_ (.CLK(clknet_leaf_193_wb_clk_i),
    .Q(\tholin_riscv.spi.dout[1] ),
    .D(net571));
 sky130_as_sc_hs__dfxtp_2 _52933_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.spi.dout[2] ),
    .D(net574));
 sky130_as_sc_hs__dfxtp_2 _52934_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.spi.dout[3] ),
    .D(net1734));
 sky130_as_sc_hs__dfxtp_2 _52935_ (.CLK(clknet_leaf_186_wb_clk_i),
    .Q(\tholin_riscv.spi.dout[4] ),
    .D(net580));
 sky130_as_sc_hs__dfxtp_2 _52936_ (.CLK(clknet_leaf_186_wb_clk_i),
    .Q(\tholin_riscv.spi.dout[5] ),
    .D(net1743));
 sky130_as_sc_hs__dfxtp_2 _52937_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.spi.dout[6] ),
    .D(net601));
 sky130_as_sc_hs__dfxtp_2 _52938_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.spi.dout[7] ),
    .D(net1730));
 sky130_as_sc_hs__dfxtp_2 _52939_ (.CLK(clknet_leaf_161_wb_clk_i),
    .Q(net58),
    .D(_01045_));
 sky130_as_sc_hs__dfxtp_2 _52940_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(net57),
    .D(_01046_));
 sky130_as_sc_hs__dfxtp_2 _52941_ (.CLK(clknet_leaf_186_wb_clk_i),
    .Q(\tholin_riscv.spi.busy ),
    .D(net610));
 sky130_as_sc_hs__dfxtp_2 _52942_ (.CLK(clknet_leaf_186_wb_clk_i),
    .Q(\tholin_riscv.spi.counter[0] ),
    .D(_01048_));
 sky130_as_sc_hs__dfxtp_2 _52943_ (.CLK(clknet_leaf_186_wb_clk_i),
    .Q(\tholin_riscv.spi.counter[1] ),
    .D(_01049_));
 sky130_as_sc_hs__dfxtp_2 _52944_ (.CLK(clknet_leaf_186_wb_clk_i),
    .Q(\tholin_riscv.spi.counter[2] ),
    .D(_01050_));
 sky130_as_sc_hs__dfxtp_2 _52945_ (.CLK(clknet_leaf_186_wb_clk_i),
    .Q(\tholin_riscv.spi.counter[3] ),
    .D(_01051_));
 sky130_as_sc_hs__dfxtp_2 _52946_ (.CLK(clknet_leaf_186_wb_clk_i),
    .Q(\tholin_riscv.spi.counter[4] ),
    .D(_01052_));
 sky130_as_sc_hs__dfxtp_2 _52947_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.spi.data_out_buff[0] ),
    .D(net1322));
 sky130_as_sc_hs__dfxtp_2 _52948_ (.CLK(clknet_leaf_187_wb_clk_i),
    .Q(\tholin_riscv.spi.data_out_buff[1] ),
    .D(_01054_));
 sky130_as_sc_hs__dfxtp_2 _52949_ (.CLK(clknet_leaf_187_wb_clk_i),
    .Q(\tholin_riscv.spi.data_out_buff[2] ),
    .D(_01055_));
 sky130_as_sc_hs__dfxtp_2 _52950_ (.CLK(clknet_leaf_187_wb_clk_i),
    .Q(\tholin_riscv.spi.data_out_buff[3] ),
    .D(_01056_));
 sky130_as_sc_hs__dfxtp_2 _52951_ (.CLK(clknet_leaf_187_wb_clk_i),
    .Q(\tholin_riscv.spi.data_out_buff[4] ),
    .D(_01057_));
 sky130_as_sc_hs__dfxtp_2 _52952_ (.CLK(clknet_leaf_186_wb_clk_i),
    .Q(\tholin_riscv.spi.data_out_buff[5] ),
    .D(_01058_));
 sky130_as_sc_hs__dfxtp_2 _52953_ (.CLK(clknet_leaf_187_wb_clk_i),
    .Q(\tholin_riscv.spi.data_out_buff[6] ),
    .D(_01059_));
 sky130_as_sc_hs__dfxtp_2 _52954_ (.CLK(clknet_leaf_187_wb_clk_i),
    .Q(\tholin_riscv.spi.data_out_buff[7] ),
    .D(_01060_));
 sky130_as_sc_hs__dfxtp_2 _52955_ (.CLK(clknet_leaf_140_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[0] ),
    .D(_01061_));
 sky130_as_sc_hs__dfxtp_2 _52956_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[1] ),
    .D(_01062_));
 sky130_as_sc_hs__dfxtp_2 _52957_ (.CLK(clknet_leaf_136_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[2] ),
    .D(_01063_));
 sky130_as_sc_hs__dfxtp_2 _52958_ (.CLK(clknet_leaf_137_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[3] ),
    .D(_01064_));
 sky130_as_sc_hs__dfxtp_2 _52959_ (.CLK(clknet_leaf_137_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[4] ),
    .D(_01065_));
 sky130_as_sc_hs__dfxtp_2 _52960_ (.CLK(clknet_leaf_136_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[5] ),
    .D(_01066_));
 sky130_as_sc_hs__dfxtp_2 _52961_ (.CLK(clknet_leaf_138_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[6] ),
    .D(_01067_));
 sky130_as_sc_hs__dfxtp_2 _52962_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[7] ),
    .D(_01068_));
 sky130_as_sc_hs__dfxtp_2 _52963_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[8] ),
    .D(_01069_));
 sky130_as_sc_hs__dfxtp_2 _52964_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[9] ),
    .D(_01070_));
 sky130_as_sc_hs__dfxtp_2 _52965_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[10] ),
    .D(_01071_));
 sky130_as_sc_hs__dfxtp_2 _52966_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[11] ),
    .D(net1345));
 sky130_as_sc_hs__dfxtp_2 _52967_ (.CLK(clknet_leaf_135_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[12] ),
    .D(_01073_));
 sky130_as_sc_hs__dfxtp_2 _52968_ (.CLK(clknet_leaf_135_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[13] ),
    .D(_01074_));
 sky130_as_sc_hs__dfxtp_2 _52969_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[14] ),
    .D(_01075_));
 sky130_as_sc_hs__dfxtp_2 _52970_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.uart.divisor[15] ),
    .D(_01076_));
 sky130_as_sc_hs__dfxtp_2 _52971_ (.CLK(clknet_leaf_187_wb_clk_i),
    .Q(\tholin_riscv.spi.divisor[0] ),
    .D(net629));
 sky130_as_sc_hs__dfxtp_2 _52972_ (.CLK(clknet_leaf_188_wb_clk_i),
    .Q(\tholin_riscv.spi.divisor[1] ),
    .D(net613));
 sky130_as_sc_hs__dfxtp_2 _52973_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.spi.divisor[2] ),
    .D(net620));
 sky130_as_sc_hs__dfxtp_2 _52974_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.spi.divisor[3] ),
    .D(net774));
 sky130_as_sc_hs__dfxtp_2 _52975_ (.CLK(clknet_leaf_181_wb_clk_i),
    .Q(\tholin_riscv.spi.divisor[4] ),
    .D(net650));
 sky130_as_sc_hs__dfxtp_2 _52976_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.spi.divisor[5] ),
    .D(net626));
 sky130_as_sc_hs__dfxtp_2 _52977_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.spi.divisor[6] ),
    .D(net753));
 sky130_as_sc_hs__dfxtp_2 _52978_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.spi.divisor[7] ),
    .D(_01084_));
 sky130_as_sc_hs__dfxtp_2 _52979_ (.CLK(clknet_leaf_192_wb_clk_i),
    .Q(\tholin_riscv.load_dest[0] ),
    .D(net647));
 sky130_as_sc_hs__dfxtp_2 _52980_ (.CLK(clknet_leaf_191_wb_clk_i),
    .Q(\tholin_riscv.load_dest[1] ),
    .D(net632));
 sky130_as_sc_hs__dfxtp_2 _52981_ (.CLK(clknet_leaf_192_wb_clk_i),
    .Q(\tholin_riscv.load_dest[2] ),
    .D(net644));
 sky130_as_sc_hs__dfxtp_2 _52982_ (.CLK(clknet_leaf_193_wb_clk_i),
    .Q(\tholin_riscv.load_dest[3] ),
    .D(net638));
 sky130_as_sc_hs__dfxtp_2 _52983_ (.CLK(clknet_leaf_194_wb_clk_i),
    .Q(\tholin_riscv.load_dest[4] ),
    .D(net635));
 sky130_as_sc_hs__dfxtp_2 _52984_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.div_counter[0] ),
    .D(_01090_));
 sky130_as_sc_hs__dfxtp_2 _52985_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.div_counter[1] ),
    .D(_01091_));
 sky130_as_sc_hs__dfxtp_2 _52986_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.div_counter[2] ),
    .D(_01092_));
 sky130_as_sc_hs__dfxtp_2 _52987_ (.CLK(clknet_leaf_180_wb_clk_i),
    .Q(\tholin_riscv.div_counter[3] ),
    .D(_01093_));
 sky130_as_sc_hs__dfxtp_2 _52988_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.div_counter[4] ),
    .D(_01094_));
 sky130_as_sc_hs__dfxtp_2 _52989_ (.CLK(clknet_leaf_200_wb_clk_i),
    .Q(\tholin_riscv.div_res[0] ),
    .D(_01095_));
 sky130_as_sc_hs__dfxtp_2 _52990_ (.CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(\tholin_riscv.div_res[1] ),
    .D(_01096_));
 sky130_as_sc_hs__dfxtp_2 _52991_ (.CLK(clknet_leaf_207_wb_clk_i),
    .Q(\tholin_riscv.div_res[2] ),
    .D(_01097_));
 sky130_as_sc_hs__dfxtp_2 _52992_ (.CLK(clknet_leaf_207_wb_clk_i),
    .Q(\tholin_riscv.div_res[3] ),
    .D(_01098_));
 sky130_as_sc_hs__dfxtp_2 _52993_ (.CLK(clknet_leaf_206_wb_clk_i),
    .Q(\tholin_riscv.div_res[4] ),
    .D(_01099_));
 sky130_as_sc_hs__dfxtp_2 _52994_ (.CLK(clknet_leaf_206_wb_clk_i),
    .Q(\tholin_riscv.div_res[5] ),
    .D(_01100_));
 sky130_as_sc_hs__dfxtp_2 _52995_ (.CLK(clknet_leaf_206_wb_clk_i),
    .Q(\tholin_riscv.div_res[6] ),
    .D(_01101_));
 sky130_as_sc_hs__dfxtp_2 _52996_ (.CLK(clknet_leaf_206_wb_clk_i),
    .Q(\tholin_riscv.div_res[7] ),
    .D(_01102_));
 sky130_as_sc_hs__dfxtp_2 _52997_ (.CLK(clknet_leaf_206_wb_clk_i),
    .Q(\tholin_riscv.div_res[8] ),
    .D(_01103_));
 sky130_as_sc_hs__dfxtp_2 _52998_ (.CLK(clknet_leaf_206_wb_clk_i),
    .Q(\tholin_riscv.div_res[9] ),
    .D(_01104_));
 sky130_as_sc_hs__dfxtp_2 _52999_ (.CLK(clknet_leaf_206_wb_clk_i),
    .Q(\tholin_riscv.div_res[10] ),
    .D(_01105_));
 sky130_as_sc_hs__dfxtp_2 _53000_ (.CLK(clknet_leaf_206_wb_clk_i),
    .Q(\tholin_riscv.div_res[11] ),
    .D(_01106_));
 sky130_as_sc_hs__dfxtp_2 _53001_ (.CLK(clknet_leaf_209_wb_clk_i),
    .Q(\tholin_riscv.div_res[12] ),
    .D(_01107_));
 sky130_as_sc_hs__dfxtp_2 _53002_ (.CLK(clknet_leaf_209_wb_clk_i),
    .Q(\tholin_riscv.div_res[13] ),
    .D(_01108_));
 sky130_as_sc_hs__dfxtp_2 _53003_ (.CLK(clknet_leaf_209_wb_clk_i),
    .Q(\tholin_riscv.div_res[14] ),
    .D(_01109_));
 sky130_as_sc_hs__dfxtp_2 _53004_ (.CLK(clknet_leaf_209_wb_clk_i),
    .Q(\tholin_riscv.div_res[15] ),
    .D(_01110_));
 sky130_as_sc_hs__dfxtp_2 _53005_ (.CLK(clknet_leaf_212_wb_clk_i),
    .Q(\tholin_riscv.div_res[16] ),
    .D(_01111_));
 sky130_as_sc_hs__dfxtp_2 _53006_ (.CLK(clknet_leaf_213_wb_clk_i),
    .Q(\tholin_riscv.div_res[17] ),
    .D(_01112_));
 sky130_as_sc_hs__dfxtp_2 _53007_ (.CLK(clknet_leaf_213_wb_clk_i),
    .Q(\tholin_riscv.div_res[18] ),
    .D(_01113_));
 sky130_as_sc_hs__dfxtp_2 _53008_ (.CLK(clknet_leaf_213_wb_clk_i),
    .Q(\tholin_riscv.div_res[19] ),
    .D(_01114_));
 sky130_as_sc_hs__dfxtp_2 _53009_ (.CLK(clknet_leaf_213_wb_clk_i),
    .Q(\tholin_riscv.div_res[20] ),
    .D(_01115_));
 sky130_as_sc_hs__dfxtp_2 _53010_ (.CLK(clknet_leaf_213_wb_clk_i),
    .Q(\tholin_riscv.div_res[21] ),
    .D(_01116_));
 sky130_as_sc_hs__dfxtp_2 _53011_ (.CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(\tholin_riscv.div_res[22] ),
    .D(_01117_));
 sky130_as_sc_hs__dfxtp_2 _53012_ (.CLK(clknet_leaf_216_wb_clk_i),
    .Q(\tholin_riscv.div_res[23] ),
    .D(_01118_));
 sky130_as_sc_hs__dfxtp_2 _53013_ (.CLK(clknet_leaf_215_wb_clk_i),
    .Q(\tholin_riscv.div_res[24] ),
    .D(_01119_));
 sky130_as_sc_hs__dfxtp_2 _53014_ (.CLK(clknet_leaf_215_wb_clk_i),
    .Q(\tholin_riscv.div_res[25] ),
    .D(_01120_));
 sky130_as_sc_hs__dfxtp_2 _53015_ (.CLK(clknet_leaf_215_wb_clk_i),
    .Q(\tholin_riscv.div_res[26] ),
    .D(_01121_));
 sky130_as_sc_hs__dfxtp_2 _53016_ (.CLK(clknet_leaf_216_wb_clk_i),
    .Q(\tholin_riscv.div_res[27] ),
    .D(_01122_));
 sky130_as_sc_hs__dfxtp_2 _53017_ (.CLK(clknet_leaf_216_wb_clk_i),
    .Q(\tholin_riscv.div_res[28] ),
    .D(_01123_));
 sky130_as_sc_hs__dfxtp_2 _53018_ (.CLK(clknet_leaf_216_wb_clk_i),
    .Q(\tholin_riscv.div_res[29] ),
    .D(_01124_));
 sky130_as_sc_hs__dfxtp_2 _53019_ (.CLK(clknet_leaf_205_wb_clk_i),
    .Q(\tholin_riscv.div_res[30] ),
    .D(_01125_));
 sky130_as_sc_hs__dfxtp_2 _53020_ (.CLK(clknet_leaf_205_wb_clk_i),
    .Q(\tholin_riscv.div_res[31] ),
    .D(_01126_));
 sky130_as_sc_hs__dfxtp_2 _53021_ (.CLK(clknet_leaf_112_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[0] ),
    .D(_01127_));
 sky130_as_sc_hs__dfxtp_2 _53022_ (.CLK(clknet_leaf_3_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[1] ),
    .D(_01128_));
 sky130_as_sc_hs__dfxtp_2 _53023_ (.CLK(clknet_leaf_8_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[2] ),
    .D(_01129_));
 sky130_as_sc_hs__dfxtp_2 _53024_ (.CLK(clknet_leaf_5_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[3] ),
    .D(_01130_));
 sky130_as_sc_hs__dfxtp_2 _53025_ (.CLK(clknet_leaf_3_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[4] ),
    .D(_01131_));
 sky130_as_sc_hs__dfxtp_2 _53026_ (.CLK(clknet_leaf_8_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[5] ),
    .D(_01132_));
 sky130_as_sc_hs__dfxtp_2 _53027_ (.CLK(clknet_leaf_2_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[6] ),
    .D(_01133_));
 sky130_as_sc_hs__dfxtp_2 _53028_ (.CLK(clknet_leaf_10_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[7] ),
    .D(_01134_));
 sky130_as_sc_hs__dfxtp_2 _53029_ (.CLK(clknet_leaf_8_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[8] ),
    .D(_01135_));
 sky130_as_sc_hs__dfxtp_2 _53030_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[9] ),
    .D(_01136_));
 sky130_as_sc_hs__dfxtp_2 _53031_ (.CLK(clknet_leaf_2_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[10] ),
    .D(_01137_));
 sky130_as_sc_hs__dfxtp_2 _53032_ (.CLK(clknet_leaf_8_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[11] ),
    .D(_01138_));
 sky130_as_sc_hs__dfxtp_2 _53033_ (.CLK(clknet_leaf_7_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[12] ),
    .D(_01139_));
 sky130_as_sc_hs__dfxtp_2 _53034_ (.CLK(clknet_leaf_2_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[13] ),
    .D(_01140_));
 sky130_as_sc_hs__dfxtp_2 _53035_ (.CLK(clknet_leaf_9_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[14] ),
    .D(_01141_));
 sky130_as_sc_hs__dfxtp_2 _53036_ (.CLK(clknet_leaf_2_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[15] ),
    .D(_01142_));
 sky130_as_sc_hs__dfxtp_2 _53037_ (.CLK(clknet_leaf_3_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[16] ),
    .D(_01143_));
 sky130_as_sc_hs__dfxtp_2 _53038_ (.CLK(clknet_leaf_2_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[17] ),
    .D(_01144_));
 sky130_as_sc_hs__dfxtp_2 _53039_ (.CLK(clknet_leaf_2_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[18] ),
    .D(_01145_));
 sky130_as_sc_hs__dfxtp_2 _53040_ (.CLK(clknet_leaf_5_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[19] ),
    .D(_01146_));
 sky130_as_sc_hs__dfxtp_2 _53041_ (.CLK(clknet_leaf_3_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[20] ),
    .D(_01147_));
 sky130_as_sc_hs__dfxtp_2 _53042_ (.CLK(clknet_leaf_11_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[21] ),
    .D(_01148_));
 sky130_as_sc_hs__dfxtp_2 _53043_ (.CLK(clknet_leaf_5_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[22] ),
    .D(_01149_));
 sky130_as_sc_hs__dfxtp_2 _53044_ (.CLK(clknet_leaf_10_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[23] ),
    .D(_01150_));
 sky130_as_sc_hs__dfxtp_2 _53045_ (.CLK(clknet_leaf_3_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[24] ),
    .D(_01151_));
 sky130_as_sc_hs__dfxtp_2 _53046_ (.CLK(clknet_leaf_4_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[25] ),
    .D(_01152_));
 sky130_as_sc_hs__dfxtp_2 _53047_ (.CLK(clknet_leaf_9_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[26] ),
    .D(_01153_));
 sky130_as_sc_hs__dfxtp_2 _53048_ (.CLK(clknet_leaf_7_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[27] ),
    .D(_01154_));
 sky130_as_sc_hs__dfxtp_2 _53049_ (.CLK(clknet_leaf_3_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[28] ),
    .D(_01155_));
 sky130_as_sc_hs__dfxtp_2 _53050_ (.CLK(clknet_leaf_5_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[29] ),
    .D(_01156_));
 sky130_as_sc_hs__dfxtp_2 _53051_ (.CLK(clknet_leaf_5_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[30] ),
    .D(_01157_));
 sky130_as_sc_hs__dfxtp_2 _53052_ (.CLK(clknet_leaf_203_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[31] ),
    .D(_01158_));
 sky130_as_sc_hs__dfxtp_2 _53053_ (.CLK(clknet_leaf_208_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[32] ),
    .D(_01159_));
 sky130_as_sc_hs__dfxtp_2 _53054_ (.CLK(clknet_leaf_207_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[33] ),
    .D(_01160_));
 sky130_as_sc_hs__dfxtp_2 _53055_ (.CLK(clknet_leaf_208_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[34] ),
    .D(_01161_));
 sky130_as_sc_hs__dfxtp_2 _53056_ (.CLK(clknet_leaf_208_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[35] ),
    .D(_01162_));
 sky130_as_sc_hs__dfxtp_2 _53057_ (.CLK(clknet_leaf_208_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[36] ),
    .D(_01163_));
 sky130_as_sc_hs__dfxtp_2 _53058_ (.CLK(clknet_leaf_208_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[37] ),
    .D(_01164_));
 sky130_as_sc_hs__dfxtp_2 _53059_ (.CLK(clknet_leaf_208_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[38] ),
    .D(_01165_));
 sky130_as_sc_hs__dfxtp_2 _53060_ (.CLK(clknet_leaf_210_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[39] ),
    .D(_01166_));
 sky130_as_sc_hs__dfxtp_2 _53061_ (.CLK(clknet_leaf_210_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[40] ),
    .D(_01167_));
 sky130_as_sc_hs__dfxtp_2 _53062_ (.CLK(clknet_leaf_210_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[41] ),
    .D(_01168_));
 sky130_as_sc_hs__dfxtp_2 _53063_ (.CLK(clknet_leaf_210_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[42] ),
    .D(_01169_));
 sky130_as_sc_hs__dfxtp_2 _53064_ (.CLK(clknet_leaf_210_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[43] ),
    .D(_01170_));
 sky130_as_sc_hs__dfxtp_2 _53065_ (.CLK(clknet_leaf_210_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[44] ),
    .D(_01171_));
 sky130_as_sc_hs__dfxtp_2 _53066_ (.CLK(clknet_leaf_211_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[45] ),
    .D(_01172_));
 sky130_as_sc_hs__dfxtp_2 _53067_ (.CLK(clknet_leaf_211_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[46] ),
    .D(_01173_));
 sky130_as_sc_hs__dfxtp_2 _53068_ (.CLK(clknet_leaf_212_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[47] ),
    .D(_01174_));
 sky130_as_sc_hs__dfxtp_2 _53069_ (.CLK(clknet_leaf_212_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[48] ),
    .D(_01175_));
 sky130_as_sc_hs__dfxtp_2 _53070_ (.CLK(clknet_leaf_212_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[49] ),
    .D(_01176_));
 sky130_as_sc_hs__dfxtp_2 _53071_ (.CLK(clknet_leaf_212_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[50] ),
    .D(_01177_));
 sky130_as_sc_hs__dfxtp_2 _53072_ (.CLK(clknet_leaf_214_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[51] ),
    .D(_01178_));
 sky130_as_sc_hs__dfxtp_2 _53073_ (.CLK(clknet_leaf_213_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[52] ),
    .D(_01179_));
 sky130_as_sc_hs__dfxtp_2 _53074_ (.CLK(clknet_leaf_213_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[53] ),
    .D(_01180_));
 sky130_as_sc_hs__dfxtp_2 _53075_ (.CLK(clknet_leaf_213_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[54] ),
    .D(_01181_));
 sky130_as_sc_hs__dfxtp_2 _53076_ (.CLK(clknet_leaf_213_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[55] ),
    .D(_01182_));
 sky130_as_sc_hs__dfxtp_2 _53077_ (.CLK(clknet_leaf_214_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[56] ),
    .D(_01183_));
 sky130_as_sc_hs__dfxtp_2 _53078_ (.CLK(clknet_leaf_214_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[57] ),
    .D(_01184_));
 sky130_as_sc_hs__dfxtp_2 _53079_ (.CLK(clknet_leaf_214_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[58] ),
    .D(_01185_));
 sky130_as_sc_hs__dfxtp_2 _53080_ (.CLK(clknet_leaf_215_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[59] ),
    .D(_01186_));
 sky130_as_sc_hs__dfxtp_2 _53081_ (.CLK(clknet_leaf_215_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[60] ),
    .D(_01187_));
 sky130_as_sc_hs__dfxtp_2 _53082_ (.CLK(clknet_leaf_215_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[61] ),
    .D(_01188_));
 sky130_as_sc_hs__dfxtp_2 _53083_ (.CLK(clknet_leaf_215_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[62] ),
    .D(_01189_));
 sky130_as_sc_hs__dfxtp_2 _53084_ (.CLK(clknet_leaf_205_wb_clk_i),
    .Q(\tholin_riscv.div_shifter[63] ),
    .D(_01190_));
 sky130_as_sc_hs__dfxtp_2 _53085_ (.CLK(clknet_leaf_192_wb_clk_i),
    .Q(\tholin_riscv.load_funct ),
    .D(net641));
 sky130_as_sc_hs__dfxtp_2 _53086_ (.CLK(clknet_leaf_156_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[0] ),
    .D(net1713));
 sky130_as_sc_hs__dfxtp_2 _53087_ (.CLK(clknet_leaf_156_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[1] ),
    .D(net771));
 sky130_as_sc_hs__dfxtp_2 _53088_ (.CLK(clknet_leaf_156_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[2] ),
    .D(net970));
 sky130_as_sc_hs__dfxtp_2 _53089_ (.CLK(clknet_leaf_156_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[3] ),
    .D(net1023));
 sky130_as_sc_hs__dfxtp_2 _53090_ (.CLK(clknet_leaf_156_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[4] ),
    .D(net825));
 sky130_as_sc_hs__dfxtp_2 _53091_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[5] ),
    .D(net854));
 sky130_as_sc_hs__dfxtp_2 _53092_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[6] ),
    .D(net1003));
 sky130_as_sc_hs__dfxtp_2 _53093_ (.CLK(clknet_leaf_165_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[7] ),
    .D(net1027));
 sky130_as_sc_hs__dfxtp_2 _53094_ (.CLK(clknet_leaf_166_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[8] ),
    .D(net1019));
 sky130_as_sc_hs__dfxtp_2 _53095_ (.CLK(clknet_leaf_165_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[9] ),
    .D(net950));
 sky130_as_sc_hs__dfxtp_2 _53096_ (.CLK(clknet_leaf_165_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[10] ),
    .D(net1052));
 sky130_as_sc_hs__dfxtp_2 _53097_ (.CLK(clknet_leaf_165_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[11] ),
    .D(net1015));
 sky130_as_sc_hs__dfxtp_2 _53098_ (.CLK(clknet_leaf_165_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[12] ),
    .D(net1126));
 sky130_as_sc_hs__dfxtp_2 _53099_ (.CLK(clknet_leaf_165_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[13] ),
    .D(net846));
 sky130_as_sc_hs__dfxtp_2 _53100_ (.CLK(clknet_leaf_165_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[14] ),
    .D(net946));
 sky130_as_sc_hs__dfxtp_2 _53101_ (.CLK(clknet_leaf_156_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[15] ),
    .D(net910));
 sky130_as_sc_hs__dfxtp_2 _53102_ (.CLK(clknet_leaf_165_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[16] ),
    .D(net862));
 sky130_as_sc_hs__dfxtp_2 _53103_ (.CLK(clknet_leaf_163_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[17] ),
    .D(net870));
 sky130_as_sc_hs__dfxtp_2 _53104_ (.CLK(clknet_leaf_163_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[18] ),
    .D(net898));
 sky130_as_sc_hs__dfxtp_2 _53105_ (.CLK(clknet_leaf_164_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[19] ),
    .D(net866));
 sky130_as_sc_hs__dfxtp_2 _53106_ (.CLK(clknet_leaf_164_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[20] ),
    .D(net1048));
 sky130_as_sc_hs__dfxtp_2 _53107_ (.CLK(clknet_leaf_164_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[21] ),
    .D(net1207));
 sky130_as_sc_hs__dfxtp_2 _53108_ (.CLK(clknet_leaf_167_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[22] ),
    .D(net906));
 sky130_as_sc_hs__dfxtp_2 _53109_ (.CLK(clknet_leaf_167_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[23] ),
    .D(net813));
 sky130_as_sc_hs__dfxtp_2 _53110_ (.CLK(clknet_leaf_166_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[24] ),
    .D(net918));
 sky130_as_sc_hs__dfxtp_2 _53111_ (.CLK(clknet_leaf_167_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[25] ),
    .D(net767));
 sky130_as_sc_hs__dfxtp_2 _53112_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[26] ),
    .D(net942));
 sky130_as_sc_hs__dfxtp_2 _53113_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[27] ),
    .D(net991));
 sky130_as_sc_hs__dfxtp_2 _53114_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[28] ),
    .D(net1092));
 sky130_as_sc_hs__dfxtp_2 _53115_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[29] ),
    .D(net1064));
 sky130_as_sc_hs__dfxtp_2 _53116_ (.CLK(clknet_leaf_184_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[30] ),
    .D(_01222_));
 sky130_as_sc_hs__dfxtp_2 _53117_ (.CLK(clknet_leaf_184_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre_ctr[31] ),
    .D(_01223_));
 sky130_as_sc_hs__dfxtp_2 _53118_ (.CLK(clknet_leaf_190_wb_clk_i),
    .Q(\tholin_riscv.cycle[0] ),
    .D(_01224_));
 sky130_as_sc_hs__dfxtp_2 _53119_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.cycle[1] ),
    .D(net1646));
 sky130_as_sc_hs__dfxtp_2 _53120_ (.CLK(clknet_leaf_180_wb_clk_i),
    .Q(\tholin_riscv.cycle[2] ),
    .D(_01226_));
 sky130_as_sc_hs__dfxtp_2 _53121_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.cycle[3] ),
    .D(_01227_));
 sky130_as_sc_hs__dfxtp_2 _53122_ (.CLK(clknet_leaf_199_wb_clk_i),
    .Q(\tholin_riscv.int_enabled ),
    .D(net759));
 sky130_as_sc_hs__dfxtp_2 _53123_ (.CLK(clknet_leaf_192_wb_clk_i),
    .Q(\tholin_riscv.ret_cycle[0] ),
    .D(_01229_));
 sky130_as_sc_hs__dfxtp_2 _53124_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.ret_cycle[1] ),
    .D(_01230_));
 sky130_as_sc_hs__dfxtp_2 _53125_ (.CLK(clknet_leaf_190_wb_clk_i),
    .Q(\tholin_riscv.io_size[0] ),
    .D(_01231_));
 sky130_as_sc_hs__dfxtp_2 _53126_ (.CLK(clknet_leaf_200_wb_clk_i),
    .Q(\tholin_riscv.io_size[1] ),
    .D(_01232_));
 sky130_as_sc_hs__dfxtp_2 _53127_ (.CLK(clknet_leaf_2_wb_clk_i),
    .Q(\tholin_riscv.Jimm[16] ),
    .D(_01233_));
 sky130_as_sc_hs__dfxtp_2 _53128_ (.CLK(clknet_leaf_127_wb_clk_i),
    .Q(\tholin_riscv.Jimm[17] ),
    .D(_01234_));
 sky130_as_sc_hs__dfxtp_2 _53129_ (.CLK(clknet_leaf_132_wb_clk_i),
    .Q(\tholin_riscv.Jimm[18] ),
    .D(_01235_));
 sky130_as_sc_hs__dfxtp_2 _53130_ (.CLK(clknet_leaf_7_wb_clk_i),
    .Q(\tholin_riscv.Jimm[19] ),
    .D(_01236_));
 sky130_as_sc_hs__dfxtp_2 _53131_ (.CLK(clknet_leaf_133_wb_clk_i),
    .Q(\tholin_riscv.Iimm[0] ),
    .D(_01237_));
 sky130_as_sc_hs__dfxtp_2 _53132_ (.CLK(clknet_leaf_196_wb_clk_i),
    .Q(\tholin_riscv.Iimm[1] ),
    .D(_01238_));
 sky130_as_sc_hs__dfxtp_2 _53133_ (.CLK(clknet_leaf_135_wb_clk_i),
    .Q(\tholin_riscv.Iimm[2] ),
    .D(_01239_));
 sky130_as_sc_hs__dfxtp_2 _53134_ (.CLK(clknet_leaf_6_wb_clk_i),
    .Q(\tholin_riscv.Iimm[3] ),
    .D(_01240_));
 sky130_as_sc_hs__dfxtp_2 _53135_ (.CLK(clknet_leaf_196_wb_clk_i),
    .Q(\tholin_riscv.Iimm[4] ),
    .D(_01241_));
 sky130_as_sc_hs__dfxtp_2 _53136_ (.CLK(clknet_leaf_193_wb_clk_i),
    .Q(\tholin_riscv.Bimm[5] ),
    .D(_01242_));
 sky130_as_sc_hs__dfxtp_2 _53137_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.Bimm[6] ),
    .D(_01243_));
 sky130_as_sc_hs__dfxtp_2 _53138_ (.CLK(clknet_leaf_197_wb_clk_i),
    .Q(\tholin_riscv.Bimm[7] ),
    .D(_01244_));
 sky130_as_sc_hs__dfxtp_2 _53139_ (.CLK(clknet_leaf_194_wb_clk_i),
    .Q(\tholin_riscv.Bimm[8] ),
    .D(_01245_));
 sky130_as_sc_hs__dfxtp_2 _53140_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.Bimm[9] ),
    .D(_01246_));
 sky130_as_sc_hs__dfxtp_2 _53141_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.Bimm[10] ),
    .D(_01247_));
 sky130_as_sc_hs__dfxtp_2 _53142_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.Bimm[12] ),
    .D(_01248_));
 sky130_as_sc_hs__dfxtp_2 _53143_ (.CLK(clknet_leaf_178_wb_clk_i),
    .Q(\tholin_riscv.is_write ),
    .D(_01249_));
 sky130_as_sc_hs__dfxtp_2 _53144_ (.CLK(clknet_leaf_189_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[0] ),
    .D(_01250_));
 sky130_as_sc_hs__dfxtp_2 _53145_ (.CLK(clknet_leaf_180_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[1] ),
    .D(_01251_));
 sky130_as_sc_hs__dfxtp_2 _53146_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[2] ),
    .D(_01252_));
 sky130_as_sc_hs__dfxtp_2 _53147_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[3] ),
    .D(_01253_));
 sky130_as_sc_hs__dfxtp_2 _53148_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[4] ),
    .D(_01254_));
 sky130_as_sc_hs__dfxtp_2 _53149_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[5] ),
    .D(_01255_));
 sky130_as_sc_hs__dfxtp_2 _53150_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[6] ),
    .D(_01256_));
 sky130_as_sc_hs__dfxtp_2 _53151_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[7] ),
    .D(_01257_));
 sky130_as_sc_hs__dfxtp_2 _53152_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[8] ),
    .D(_01258_));
 sky130_as_sc_hs__dfxtp_2 _53153_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[9] ),
    .D(_01259_));
 sky130_as_sc_hs__dfxtp_2 _53154_ (.CLK(clknet_leaf_211_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[10] ),
    .D(_01260_));
 sky130_as_sc_hs__dfxtp_2 _53155_ (.CLK(clknet_leaf_211_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[11] ),
    .D(_01261_));
 sky130_as_sc_hs__dfxtp_2 _53156_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[12] ),
    .D(_01262_));
 sky130_as_sc_hs__dfxtp_2 _53157_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[13] ),
    .D(_01263_));
 sky130_as_sc_hs__dfxtp_2 _53158_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[14] ),
    .D(_01264_));
 sky130_as_sc_hs__dfxtp_2 _53159_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[15] ),
    .D(_01265_));
 sky130_as_sc_hs__dfxtp_2 _53160_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[16] ),
    .D(_01266_));
 sky130_as_sc_hs__dfxtp_2 _53161_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[17] ),
    .D(_01267_));
 sky130_as_sc_hs__dfxtp_2 _53162_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[18] ),
    .D(_01268_));
 sky130_as_sc_hs__dfxtp_2 _53163_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[19] ),
    .D(_01269_));
 sky130_as_sc_hs__dfxtp_2 _53164_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[20] ),
    .D(_01270_));
 sky130_as_sc_hs__dfxtp_2 _53165_ (.CLK(clknet_leaf_210_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[21] ),
    .D(_01271_));
 sky130_as_sc_hs__dfxtp_2 _53166_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[22] ),
    .D(_01272_));
 sky130_as_sc_hs__dfxtp_2 _53167_ (.CLK(clknet_leaf_210_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[23] ),
    .D(_01273_));
 sky130_as_sc_hs__dfxtp_2 _53168_ (.CLK(clknet_leaf_211_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[24] ),
    .D(_01274_));
 sky130_as_sc_hs__dfxtp_2 _53169_ (.CLK(clknet_leaf_211_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[25] ),
    .D(_01275_));
 sky130_as_sc_hs__dfxtp_2 _53170_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[26] ),
    .D(_01276_));
 sky130_as_sc_hs__dfxtp_2 _53171_ (.CLK(clknet_leaf_211_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[27] ),
    .D(_01277_));
 sky130_as_sc_hs__dfxtp_2 _53172_ (.CLK(clknet_leaf_210_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[28] ),
    .D(_01278_));
 sky130_as_sc_hs__dfxtp_2 _53173_ (.CLK(clknet_leaf_211_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[29] ),
    .D(_01279_));
 sky130_as_sc_hs__dfxtp_2 _53174_ (.CLK(clknet_leaf_211_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[30] ),
    .D(_01280_));
 sky130_as_sc_hs__dfxtp_2 _53175_ (.CLK(clknet_leaf_211_wb_clk_i),
    .Q(\tholin_riscv.requested_addr[31] ),
    .D(_01281_));
 sky130_as_sc_hs__dfxtp_2 _53176_ (.CLK(clknet_leaf_218_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[0] ),
    .D(_01282_));
 sky130_as_sc_hs__dfxtp_2 _53177_ (.CLK(clknet_leaf_218_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[1] ),
    .D(_01283_));
 sky130_as_sc_hs__dfxtp_2 _53178_ (.CLK(clknet_leaf_215_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[2] ),
    .D(_01284_));
 sky130_as_sc_hs__dfxtp_2 _53179_ (.CLK(clknet_leaf_218_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[3] ),
    .D(_01285_));
 sky130_as_sc_hs__dfxtp_2 _53180_ (.CLK(clknet_leaf_216_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[4] ),
    .D(_01286_));
 sky130_as_sc_hs__dfxtp_2 _53181_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[5] ),
    .D(net1269));
 sky130_as_sc_hs__dfxtp_2 _53182_ (.CLK(clknet_leaf_178_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[6] ),
    .D(_01288_));
 sky130_as_sc_hs__dfxtp_2 _53183_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[7] ),
    .D(net1150));
 sky130_as_sc_hs__dfxtp_2 _53184_ (.CLK(clknet_leaf_178_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[8] ),
    .D(net1244));
 sky130_as_sc_hs__dfxtp_2 _53185_ (.CLK(clknet_leaf_178_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[9] ),
    .D(net1273));
 sky130_as_sc_hs__dfxtp_2 _53186_ (.CLK(clknet_leaf_215_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[10] ),
    .D(_01292_));
 sky130_as_sc_hs__dfxtp_2 _53187_ (.CLK(clknet_leaf_215_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[11] ),
    .D(_01293_));
 sky130_as_sc_hs__dfxtp_2 _53188_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[12] ),
    .D(_01294_));
 sky130_as_sc_hs__dfxtp_2 _53189_ (.CLK(clknet_leaf_218_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[13] ),
    .D(_01295_));
 sky130_as_sc_hs__dfxtp_2 _53190_ (.CLK(clknet_leaf_204_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[14] ),
    .D(_01296_));
 sky130_as_sc_hs__dfxtp_2 _53191_ (.CLK(clknet_leaf_215_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[15] ),
    .D(_01297_));
 sky130_as_sc_hs__dfxtp_2 _53192_ (.CLK(clknet_leaf_215_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[16] ),
    .D(_01298_));
 sky130_as_sc_hs__dfxtp_2 _53193_ (.CLK(clknet_leaf_204_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[17] ),
    .D(_01299_));
 sky130_as_sc_hs__dfxtp_2 _53194_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[18] ),
    .D(_01300_));
 sky130_as_sc_hs__dfxtp_2 _53195_ (.CLK(clknet_leaf_218_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[19] ),
    .D(_01301_));
 sky130_as_sc_hs__dfxtp_2 _53196_ (.CLK(clknet_leaf_204_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[20] ),
    .D(_01302_));
 sky130_as_sc_hs__dfxtp_2 _53197_ (.CLK(clknet_leaf_218_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[21] ),
    .D(_01303_));
 sky130_as_sc_hs__dfxtp_2 _53198_ (.CLK(clknet_leaf_215_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[22] ),
    .D(_01304_));
 sky130_as_sc_hs__dfxtp_2 _53199_ (.CLK(clknet_leaf_204_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[23] ),
    .D(_01305_));
 sky130_as_sc_hs__dfxtp_2 _53200_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[24] ),
    .D(net1154));
 sky130_as_sc_hs__dfxtp_2 _53201_ (.CLK(clknet_leaf_218_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[25] ),
    .D(_01307_));
 sky130_as_sc_hs__dfxtp_2 _53202_ (.CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[26] ),
    .D(_01308_));
 sky130_as_sc_hs__dfxtp_2 _53203_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[27] ),
    .D(_01309_));
 sky130_as_sc_hs__dfxtp_2 _53204_ (.CLK(clknet_leaf_203_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[28] ),
    .D(_01310_));
 sky130_as_sc_hs__dfxtp_2 _53205_ (.CLK(clknet_leaf_179_wb_clk_i),
    .Q(\tholin_riscv.intr_vec[29] ),
    .D(net1119));
 sky130_as_sc_hs__dfxtp_2 _53206_ (.CLK(clknet_leaf_145_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[0] ),
    .D(net1716));
 sky130_as_sc_hs__dfxtp_2 _53207_ (.CLK(clknet_leaf_144_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[1] ),
    .D(net750));
 sky130_as_sc_hs__dfxtp_2 _53208_ (.CLK(clknet_leaf_145_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[2] ),
    .D(net887));
 sky130_as_sc_hs__dfxtp_2 _53209_ (.CLK(clknet_leaf_144_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[3] ),
    .D(net966));
 sky130_as_sc_hs__dfxtp_2 _53210_ (.CLK(clknet_leaf_144_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[4] ),
    .D(net987));
 sky130_as_sc_hs__dfxtp_2 _53211_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[5] ),
    .D(net883));
 sky130_as_sc_hs__dfxtp_2 _53212_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[6] ),
    .D(net1112));
 sky130_as_sc_hs__dfxtp_2 _53213_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[7] ),
    .D(net930));
 sky130_as_sc_hs__dfxtp_2 _53214_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[8] ),
    .D(net1007));
 sky130_as_sc_hs__dfxtp_2 _53215_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[9] ),
    .D(net1011));
 sky130_as_sc_hs__dfxtp_2 _53216_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[10] ),
    .D(net983));
 sky130_as_sc_hs__dfxtp_2 _53217_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[11] ),
    .D(net979));
 sky130_as_sc_hs__dfxtp_2 _53218_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[12] ),
    .D(net1031));
 sky130_as_sc_hs__dfxtp_2 _53219_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[13] ),
    .D(net922));
 sky130_as_sc_hs__dfxtp_2 _53220_ (.CLK(clknet_leaf_154_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[14] ),
    .D(net999));
 sky130_as_sc_hs__dfxtp_2 _53221_ (.CLK(clknet_leaf_154_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[15] ),
    .D(net1068));
 sky130_as_sc_hs__dfxtp_2 _53222_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[16] ),
    .D(net1056));
 sky130_as_sc_hs__dfxtp_2 _53223_ (.CLK(clknet_leaf_154_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[17] ),
    .D(net938));
 sky130_as_sc_hs__dfxtp_2 _53224_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[18] ),
    .D(net902));
 sky130_as_sc_hs__dfxtp_2 _53225_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[19] ),
    .D(net1041));
 sky130_as_sc_hs__dfxtp_2 _53226_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[20] ),
    .D(net914));
 sky130_as_sc_hs__dfxtp_2 _53227_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[21] ),
    .D(net894));
 sky130_as_sc_hs__dfxtp_2 _53228_ (.CLK(clknet_leaf_142_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[22] ),
    .D(net934));
 sky130_as_sc_hs__dfxtp_2 _53229_ (.CLK(clknet_leaf_184_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[23] ),
    .D(net1037));
 sky130_as_sc_hs__dfxtp_2 _53230_ (.CLK(clknet_leaf_184_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[24] ),
    .D(net995));
 sky130_as_sc_hs__dfxtp_2 _53231_ (.CLK(clknet_leaf_184_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[25] ),
    .D(net763));
 sky130_as_sc_hs__dfxtp_2 _53232_ (.CLK(clknet_leaf_184_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[26] ),
    .D(net962));
 sky130_as_sc_hs__dfxtp_2 _53233_ (.CLK(clknet_leaf_142_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[27] ),
    .D(net1060));
 sky130_as_sc_hs__dfxtp_2 _53234_ (.CLK(clknet_leaf_142_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[28] ),
    .D(net1099));
 sky130_as_sc_hs__dfxtp_2 _53235_ (.CLK(clknet_leaf_142_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[29] ),
    .D(net958));
 sky130_as_sc_hs__dfxtp_2 _53236_ (.CLK(clknet_leaf_141_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[30] ),
    .D(net778));
 sky130_as_sc_hs__dfxtp_2 _53237_ (.CLK(clknet_leaf_142_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre_ctr[31] ),
    .D(_01343_));
 sky130_as_sc_hs__dfxtp_2 _53238_ (.CLK(clknet_leaf_169_wb_clk_i),
    .Q(\tholin_riscv.tmr1[0] ),
    .D(_01344_));
 sky130_as_sc_hs__dfxtp_2 _53239_ (.CLK(clknet_leaf_169_wb_clk_i),
    .Q(\tholin_riscv.tmr1[1] ),
    .D(net786));
 sky130_as_sc_hs__dfxtp_2 _53240_ (.CLK(clknet_leaf_169_wb_clk_i),
    .Q(\tholin_riscv.tmr1[2] ),
    .D(_01346_));
 sky130_as_sc_hs__dfxtp_2 _53241_ (.CLK(clknet_leaf_172_wb_clk_i),
    .Q(\tholin_riscv.tmr1[3] ),
    .D(_01347_));
 sky130_as_sc_hs__dfxtp_2 _53242_ (.CLK(clknet_leaf_172_wb_clk_i),
    .Q(\tholin_riscv.tmr1[4] ),
    .D(_01348_));
 sky130_as_sc_hs__dfxtp_2 _53243_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(\tholin_riscv.tmr1[5] ),
    .D(_01349_));
 sky130_as_sc_hs__dfxtp_2 _53244_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1[6] ),
    .D(_01350_));
 sky130_as_sc_hs__dfxtp_2 _53245_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1[7] ),
    .D(_01351_));
 sky130_as_sc_hs__dfxtp_2 _53246_ (.CLK(clknet_leaf_167_wb_clk_i),
    .Q(\tholin_riscv.tmr1[8] ),
    .D(_01352_));
 sky130_as_sc_hs__dfxtp_2 _53247_ (.CLK(clknet_leaf_167_wb_clk_i),
    .Q(\tholin_riscv.tmr1[9] ),
    .D(net1072));
 sky130_as_sc_hs__dfxtp_2 _53248_ (.CLK(clknet_leaf_164_wb_clk_i),
    .Q(\tholin_riscv.tmr1[10] ),
    .D(_01354_));
 sky130_as_sc_hs__dfxtp_2 _53249_ (.CLK(clknet_leaf_162_wb_clk_i),
    .Q(\tholin_riscv.tmr1[11] ),
    .D(_01355_));
 sky130_as_sc_hs__dfxtp_2 _53250_ (.CLK(clknet_leaf_162_wb_clk_i),
    .Q(\tholin_riscv.tmr1[12] ),
    .D(_01356_));
 sky130_as_sc_hs__dfxtp_2 _53251_ (.CLK(clknet_leaf_162_wb_clk_i),
    .Q(\tholin_riscv.tmr1[13] ),
    .D(_01357_));
 sky130_as_sc_hs__dfxtp_2 _53252_ (.CLK(clknet_leaf_161_wb_clk_i),
    .Q(\tholin_riscv.tmr1[14] ),
    .D(_01358_));
 sky130_as_sc_hs__dfxtp_2 _53253_ (.CLK(clknet_leaf_161_wb_clk_i),
    .Q(\tholin_riscv.tmr1[15] ),
    .D(_01359_));
 sky130_as_sc_hs__dfxtp_2 _53254_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(\tholin_riscv.tmr1[16] ),
    .D(net834));
 sky130_as_sc_hs__dfxtp_2 _53255_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(\tholin_riscv.tmr1[17] ),
    .D(_01361_));
 sky130_as_sc_hs__dfxtp_2 _53256_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(\tholin_riscv.tmr1[18] ),
    .D(_01362_));
 sky130_as_sc_hs__dfxtp_2 _53257_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(\tholin_riscv.tmr1[19] ),
    .D(_01363_));
 sky130_as_sc_hs__dfxtp_2 _53258_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1[20] ),
    .D(_01364_));
 sky130_as_sc_hs__dfxtp_2 _53259_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1[21] ),
    .D(_01365_));
 sky130_as_sc_hs__dfxtp_2 _53260_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1[22] ),
    .D(_01366_));
 sky130_as_sc_hs__dfxtp_2 _53261_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1[23] ),
    .D(_01367_));
 sky130_as_sc_hs__dfxtp_2 _53262_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1[24] ),
    .D(_01368_));
 sky130_as_sc_hs__dfxtp_2 _53263_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1[25] ),
    .D(_01369_));
 sky130_as_sc_hs__dfxtp_2 _53264_ (.CLK(clknet_leaf_182_wb_clk_i),
    .Q(\tholin_riscv.tmr1[26] ),
    .D(_01370_));
 sky130_as_sc_hs__dfxtp_2 _53265_ (.CLK(clknet_leaf_168_wb_clk_i),
    .Q(\tholin_riscv.tmr1[27] ),
    .D(_01371_));
 sky130_as_sc_hs__dfxtp_2 _53266_ (.CLK(clknet_leaf_167_wb_clk_i),
    .Q(\tholin_riscv.tmr1[28] ),
    .D(_01372_));
 sky130_as_sc_hs__dfxtp_2 _53267_ (.CLK(clknet_leaf_167_wb_clk_i),
    .Q(\tholin_riscv.tmr1[29] ),
    .D(_01373_));
 sky130_as_sc_hs__dfxtp_2 _53268_ (.CLK(clknet_leaf_167_wb_clk_i),
    .Q(\tholin_riscv.tmr1[30] ),
    .D(_01374_));
 sky130_as_sc_hs__dfxtp_2 _53269_ (.CLK(clknet_leaf_168_wb_clk_i),
    .Q(\tholin_riscv.tmr1[31] ),
    .D(_01375_));
 sky130_as_sc_hs__dfxtp_2 _53270_ (.CLK(clknet_leaf_169_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[0] ),
    .D(_01376_));
 sky130_as_sc_hs__dfxtp_2 _53271_ (.CLK(clknet_leaf_169_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[1] ),
    .D(_01377_));
 sky130_as_sc_hs__dfxtp_2 _53272_ (.CLK(clknet_leaf_172_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[2] ),
    .D(_01378_));
 sky130_as_sc_hs__dfxtp_2 _53273_ (.CLK(clknet_leaf_172_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[3] ),
    .D(_01379_));
 sky130_as_sc_hs__dfxtp_2 _53274_ (.CLK(clknet_leaf_172_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[4] ),
    .D(_01380_));
 sky130_as_sc_hs__dfxtp_2 _53275_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[5] ),
    .D(_01381_));
 sky130_as_sc_hs__dfxtp_2 _53276_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[6] ),
    .D(_01382_));
 sky130_as_sc_hs__dfxtp_2 _53277_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[7] ),
    .D(_01383_));
 sky130_as_sc_hs__dfxtp_2 _53278_ (.CLK(clknet_leaf_167_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[8] ),
    .D(_01384_));
 sky130_as_sc_hs__dfxtp_2 _53279_ (.CLK(clknet_leaf_167_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[9] ),
    .D(_01385_));
 sky130_as_sc_hs__dfxtp_2 _53280_ (.CLK(clknet_leaf_163_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[10] ),
    .D(_01386_));
 sky130_as_sc_hs__dfxtp_2 _53281_ (.CLK(clknet_leaf_164_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[11] ),
    .D(_01387_));
 sky130_as_sc_hs__dfxtp_2 _53282_ (.CLK(clknet_leaf_162_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[12] ),
    .D(_01388_));
 sky130_as_sc_hs__dfxtp_2 _53283_ (.CLK(clknet_leaf_162_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[13] ),
    .D(_01389_));
 sky130_as_sc_hs__dfxtp_2 _53284_ (.CLK(clknet_leaf_161_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[14] ),
    .D(_01390_));
 sky130_as_sc_hs__dfxtp_2 _53285_ (.CLK(clknet_leaf_161_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[15] ),
    .D(_01391_));
 sky130_as_sc_hs__dfxtp_2 _53286_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[16] ),
    .D(_01392_));
 sky130_as_sc_hs__dfxtp_2 _53287_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[17] ),
    .D(_01393_));
 sky130_as_sc_hs__dfxtp_2 _53288_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[18] ),
    .D(_01394_));
 sky130_as_sc_hs__dfxtp_2 _53289_ (.CLK(clknet_leaf_171_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[19] ),
    .D(_01395_));
 sky130_as_sc_hs__dfxtp_2 _53290_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[20] ),
    .D(_01396_));
 sky130_as_sc_hs__dfxtp_2 _53291_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[21] ),
    .D(_01397_));
 sky130_as_sc_hs__dfxtp_2 _53292_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[22] ),
    .D(_01398_));
 sky130_as_sc_hs__dfxtp_2 _53293_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[23] ),
    .D(_01399_));
 sky130_as_sc_hs__dfxtp_2 _53294_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[24] ),
    .D(_01400_));
 sky130_as_sc_hs__dfxtp_2 _53295_ (.CLK(clknet_leaf_170_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[25] ),
    .D(_01401_));
 sky130_as_sc_hs__dfxtp_2 _53296_ (.CLK(clknet_leaf_168_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[26] ),
    .D(_01402_));
 sky130_as_sc_hs__dfxtp_2 _53297_ (.CLK(clknet_leaf_168_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[27] ),
    .D(_01403_));
 sky130_as_sc_hs__dfxtp_2 _53298_ (.CLK(clknet_leaf_167_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[28] ),
    .D(_01404_));
 sky130_as_sc_hs__dfxtp_2 _53299_ (.CLK(clknet_leaf_167_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[29] ),
    .D(_01405_));
 sky130_as_sc_hs__dfxtp_2 _53300_ (.CLK(clknet_leaf_169_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[30] ),
    .D(_01406_));
 sky130_as_sc_hs__dfxtp_2 _53301_ (.CLK(clknet_leaf_168_wb_clk_i),
    .Q(\tholin_riscv.tmr1_top[31] ),
    .D(_01407_));
 sky130_as_sc_hs__dfxtp_2 _53302_ (.CLK(clknet_leaf_177_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[0] ),
    .D(_01408_));
 sky130_as_sc_hs__dfxtp_2 _53303_ (.CLK(clknet_leaf_177_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[1] ),
    .D(_01409_));
 sky130_as_sc_hs__dfxtp_2 _53304_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[2] ),
    .D(_01410_));
 sky130_as_sc_hs__dfxtp_2 _53305_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[3] ),
    .D(_01411_));
 sky130_as_sc_hs__dfxtp_2 _53306_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[4] ),
    .D(_01412_));
 sky130_as_sc_hs__dfxtp_2 _53307_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[5] ),
    .D(_01413_));
 sky130_as_sc_hs__dfxtp_2 _53308_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[6] ),
    .D(_01414_));
 sky130_as_sc_hs__dfxtp_2 _53309_ (.CLK(clknet_leaf_174_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[7] ),
    .D(_01415_));
 sky130_as_sc_hs__dfxtp_2 _53310_ (.CLK(clknet_leaf_182_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[8] ),
    .D(_01416_));
 sky130_as_sc_hs__dfxtp_2 _53311_ (.CLK(clknet_leaf_182_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[9] ),
    .D(_01417_));
 sky130_as_sc_hs__dfxtp_2 _53312_ (.CLK(clknet_leaf_168_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[10] ),
    .D(_01418_));
 sky130_as_sc_hs__dfxtp_2 _53313_ (.CLK(clknet_leaf_169_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[11] ),
    .D(_01419_));
 sky130_as_sc_hs__dfxtp_2 _53314_ (.CLK(clknet_leaf_173_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[12] ),
    .D(_01420_));
 sky130_as_sc_hs__dfxtp_2 _53315_ (.CLK(clknet_leaf_172_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[13] ),
    .D(_01421_));
 sky130_as_sc_hs__dfxtp_2 _53316_ (.CLK(clknet_leaf_174_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[14] ),
    .D(_01422_));
 sky130_as_sc_hs__dfxtp_2 _53317_ (.CLK(clknet_leaf_174_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[15] ),
    .D(_01423_));
 sky130_as_sc_hs__dfxtp_2 _53318_ (.CLK(clknet_leaf_174_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[16] ),
    .D(_01424_));
 sky130_as_sc_hs__dfxtp_2 _53319_ (.CLK(clknet_leaf_174_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[17] ),
    .D(_01425_));
 sky130_as_sc_hs__dfxtp_2 _53320_ (.CLK(clknet_leaf_172_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[18] ),
    .D(_01426_));
 sky130_as_sc_hs__dfxtp_2 _53321_ (.CLK(clknet_leaf_172_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[19] ),
    .D(_01427_));
 sky130_as_sc_hs__dfxtp_2 _53322_ (.CLK(clknet_leaf_177_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[20] ),
    .D(_01428_));
 sky130_as_sc_hs__dfxtp_2 _53323_ (.CLK(clknet_leaf_177_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[21] ),
    .D(_01429_));
 sky130_as_sc_hs__dfxtp_2 _53324_ (.CLK(clknet_leaf_174_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[22] ),
    .D(_01430_));
 sky130_as_sc_hs__dfxtp_2 _53325_ (.CLK(clknet_leaf_173_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[23] ),
    .D(_01431_));
 sky130_as_sc_hs__dfxtp_2 _53326_ (.CLK(clknet_leaf_173_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[24] ),
    .D(_01432_));
 sky130_as_sc_hs__dfxtp_2 _53327_ (.CLK(clknet_leaf_177_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[25] ),
    .D(_01433_));
 sky130_as_sc_hs__dfxtp_2 _53328_ (.CLK(clknet_leaf_178_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[26] ),
    .D(_01434_));
 sky130_as_sc_hs__dfxtp_2 _53329_ (.CLK(clknet_leaf_178_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[27] ),
    .D(_01435_));
 sky130_as_sc_hs__dfxtp_2 _53330_ (.CLK(clknet_leaf_178_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[28] ),
    .D(_01436_));
 sky130_as_sc_hs__dfxtp_2 _53331_ (.CLK(clknet_leaf_178_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[29] ),
    .D(_01437_));
 sky130_as_sc_hs__dfxtp_2 _53332_ (.CLK(clknet_leaf_182_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[30] ),
    .D(_01438_));
 sky130_as_sc_hs__dfxtp_2 _53333_ (.CLK(clknet_leaf_182_wb_clk_i),
    .Q(\tholin_riscv.tmr0_top[31] ),
    .D(_01439_));
 sky130_as_sc_hs__dfxtp_2 _53334_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[0] ),
    .D(net1188));
 sky130_as_sc_hs__dfxtp_2 _53335_ (.CLK(clknet_leaf_156_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[1] ),
    .D(net1379));
 sky130_as_sc_hs__dfxtp_2 _53336_ (.CLK(clknet_leaf_156_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[2] ),
    .D(_01442_));
 sky130_as_sc_hs__dfxtp_2 _53337_ (.CLK(clknet_leaf_156_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[3] ),
    .D(_01443_));
 sky130_as_sc_hs__dfxtp_2 _53338_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[4] ),
    .D(_01444_));
 sky130_as_sc_hs__dfxtp_2 _53339_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[5] ),
    .D(_01445_));
 sky130_as_sc_hs__dfxtp_2 _53340_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[6] ),
    .D(_01446_));
 sky130_as_sc_hs__dfxtp_2 _53341_ (.CLK(clknet_leaf_184_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[7] ),
    .D(_01447_));
 sky130_as_sc_hs__dfxtp_2 _53342_ (.CLK(clknet_leaf_166_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[8] ),
    .D(net1482));
 sky130_as_sc_hs__dfxtp_2 _53343_ (.CLK(clknet_leaf_166_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[9] ),
    .D(_01449_));
 sky130_as_sc_hs__dfxtp_2 _53344_ (.CLK(clknet_leaf_166_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[10] ),
    .D(_01450_));
 sky130_as_sc_hs__dfxtp_2 _53345_ (.CLK(clknet_leaf_166_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[11] ),
    .D(_01451_));
 sky130_as_sc_hs__dfxtp_2 _53346_ (.CLK(clknet_leaf_166_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[12] ),
    .D(_01452_));
 sky130_as_sc_hs__dfxtp_2 _53347_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[13] ),
    .D(_01453_));
 sky130_as_sc_hs__dfxtp_2 _53348_ (.CLK(clknet_leaf_164_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[14] ),
    .D(_01454_));
 sky130_as_sc_hs__dfxtp_2 _53349_ (.CLK(clknet_leaf_156_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[15] ),
    .D(_01455_));
 sky130_as_sc_hs__dfxtp_2 _53350_ (.CLK(clknet_leaf_156_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[16] ),
    .D(_01456_));
 sky130_as_sc_hs__dfxtp_2 _53351_ (.CLK(clknet_leaf_163_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[17] ),
    .D(_01457_));
 sky130_as_sc_hs__dfxtp_2 _53352_ (.CLK(clknet_leaf_163_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[18] ),
    .D(_01458_));
 sky130_as_sc_hs__dfxtp_2 _53353_ (.CLK(clknet_leaf_164_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[19] ),
    .D(_01459_));
 sky130_as_sc_hs__dfxtp_2 _53354_ (.CLK(clknet_leaf_164_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[20] ),
    .D(_01460_));
 sky130_as_sc_hs__dfxtp_2 _53355_ (.CLK(clknet_leaf_164_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[21] ),
    .D(_01461_));
 sky130_as_sc_hs__dfxtp_2 _53356_ (.CLK(clknet_leaf_166_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[22] ),
    .D(_01462_));
 sky130_as_sc_hs__dfxtp_2 _53357_ (.CLK(clknet_leaf_167_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[23] ),
    .D(_01463_));
 sky130_as_sc_hs__dfxtp_2 _53358_ (.CLK(clknet_leaf_166_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[24] ),
    .D(_01464_));
 sky130_as_sc_hs__dfxtp_2 _53359_ (.CLK(clknet_leaf_182_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[25] ),
    .D(net1418));
 sky130_as_sc_hs__dfxtp_2 _53360_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[26] ),
    .D(net1583));
 sky130_as_sc_hs__dfxtp_2 _53361_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[27] ),
    .D(_01467_));
 sky130_as_sc_hs__dfxtp_2 _53362_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[28] ),
    .D(_01468_));
 sky130_as_sc_hs__dfxtp_2 _53363_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[29] ),
    .D(net1558));
 sky130_as_sc_hs__dfxtp_2 _53364_ (.CLK(clknet_leaf_184_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[30] ),
    .D(net1472));
 sky130_as_sc_hs__dfxtp_2 _53365_ (.CLK(clknet_leaf_183_wb_clk_i),
    .Q(\tholin_riscv.tmr1_pre[31] ),
    .D(net1505));
 sky130_as_sc_hs__dfxtp_2 _53366_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[0] ),
    .D(net1134));
 sky130_as_sc_hs__dfxtp_2 _53367_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[1] ),
    .D(net1465));
 sky130_as_sc_hs__dfxtp_2 _53368_ (.CLK(clknet_leaf_145_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[2] ),
    .D(_01474_));
 sky130_as_sc_hs__dfxtp_2 _53369_ (.CLK(clknet_leaf_144_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[3] ),
    .D(_01475_));
 sky130_as_sc_hs__dfxtp_2 _53370_ (.CLK(clknet_leaf_144_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[4] ),
    .D(_01476_));
 sky130_as_sc_hs__dfxtp_2 _53371_ (.CLK(clknet_leaf_144_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[5] ),
    .D(_01477_));
 sky130_as_sc_hs__dfxtp_2 _53372_ (.CLK(clknet_leaf_141_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[6] ),
    .D(_01478_));
 sky130_as_sc_hs__dfxtp_2 _53373_ (.CLK(clknet_leaf_141_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[7] ),
    .D(net1407));
 sky130_as_sc_hs__dfxtp_2 _53374_ (.CLK(clknet_leaf_141_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[8] ),
    .D(net1262));
 sky130_as_sc_hs__dfxtp_2 _53375_ (.CLK(clknet_leaf_141_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[9] ),
    .D(net1333));
 sky130_as_sc_hs__dfxtp_2 _53376_ (.CLK(clknet_leaf_141_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[10] ),
    .D(net1414));
 sky130_as_sc_hs__dfxtp_2 _53377_ (.CLK(clknet_leaf_142_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[11] ),
    .D(net1489));
 sky130_as_sc_hs__dfxtp_2 _53378_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[12] ),
    .D(_01484_));
 sky130_as_sc_hs__dfxtp_2 _53379_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[13] ),
    .D(_01485_));
 sky130_as_sc_hs__dfxtp_2 _53380_ (.CLK(clknet_leaf_143_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[14] ),
    .D(net1532));
 sky130_as_sc_hs__dfxtp_2 _53381_ (.CLK(clknet_leaf_154_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[15] ),
    .D(_01487_));
 sky130_as_sc_hs__dfxtp_2 _53382_ (.CLK(clknet_leaf_154_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[16] ),
    .D(_01488_));
 sky130_as_sc_hs__dfxtp_2 _53383_ (.CLK(clknet_leaf_154_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[17] ),
    .D(_01489_));
 sky130_as_sc_hs__dfxtp_2 _53384_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[18] ),
    .D(_01490_));
 sky130_as_sc_hs__dfxtp_2 _53385_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[19] ),
    .D(_01491_));
 sky130_as_sc_hs__dfxtp_2 _53386_ (.CLK(clknet_leaf_142_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[20] ),
    .D(_01492_));
 sky130_as_sc_hs__dfxtp_2 _53387_ (.CLK(clknet_leaf_155_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[21] ),
    .D(_01493_));
 sky130_as_sc_hs__dfxtp_2 _53388_ (.CLK(clknet_leaf_142_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[22] ),
    .D(_01494_));
 sky130_as_sc_hs__dfxtp_2 _53389_ (.CLK(clknet_leaf_184_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[23] ),
    .D(_01495_));
 sky130_as_sc_hs__dfxtp_2 _53390_ (.CLK(clknet_leaf_184_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[24] ),
    .D(_01496_));
 sky130_as_sc_hs__dfxtp_2 _53391_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[25] ),
    .D(net1367));
 sky130_as_sc_hs__dfxtp_2 _53392_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[26] ),
    .D(net1587));
 sky130_as_sc_hs__dfxtp_2 _53393_ (.CLK(clknet_leaf_184_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[27] ),
    .D(_01499_));
 sky130_as_sc_hs__dfxtp_2 _53394_ (.CLK(clknet_leaf_184_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[28] ),
    .D(_01500_));
 sky130_as_sc_hs__dfxtp_2 _53395_ (.CLK(clknet_leaf_185_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[29] ),
    .D(net1554));
 sky130_as_sc_hs__dfxtp_2 _53396_ (.CLK(clknet_leaf_141_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[30] ),
    .D(net1437));
 sky130_as_sc_hs__dfxtp_2 _53397_ (.CLK(clknet_leaf_140_wb_clk_i),
    .Q(\tholin_riscv.tmr0_pre[31] ),
    .D(_01503_));
 sky130_as_sc_hs__dfxtp_2 _53398_ (.CLK(clknet_leaf_178_wb_clk_i),
    .Q(\tholin_riscv.tmr0[0] ),
    .D(_01504_));
 sky130_as_sc_hs__dfxtp_2 _53399_ (.CLK(clknet_leaf_178_wb_clk_i),
    .Q(\tholin_riscv.tmr0[1] ),
    .D(net782));
 sky130_as_sc_hs__dfxtp_2 _53400_ (.CLK(clknet_leaf_177_wb_clk_i),
    .Q(\tholin_riscv.tmr0[2] ),
    .D(_01506_));
 sky130_as_sc_hs__dfxtp_2 _53401_ (.CLK(clknet_leaf_177_wb_clk_i),
    .Q(\tholin_riscv.tmr0[3] ),
    .D(_01507_));
 sky130_as_sc_hs__dfxtp_2 _53402_ (.CLK(clknet_leaf_176_wb_clk_i),
    .Q(\tholin_riscv.tmr0[4] ),
    .D(_01508_));
 sky130_as_sc_hs__dfxtp_2 _53403_ (.CLK(clknet_leaf_175_wb_clk_i),
    .Q(\tholin_riscv.tmr0[5] ),
    .D(_01509_));
 sky130_as_sc_hs__dfxtp_2 _53404_ (.CLK(clknet_leaf_174_wb_clk_i),
    .Q(\tholin_riscv.tmr0[6] ),
    .D(_01510_));
 sky130_as_sc_hs__dfxtp_2 _53405_ (.CLK(clknet_leaf_174_wb_clk_i),
    .Q(\tholin_riscv.tmr0[7] ),
    .D(_01511_));
 sky130_as_sc_hs__dfxtp_2 _53406_ (.CLK(clknet_leaf_182_wb_clk_i),
    .Q(\tholin_riscv.tmr0[8] ),
    .D(_01512_));
 sky130_as_sc_hs__dfxtp_2 _53407_ (.CLK(clknet_leaf_182_wb_clk_i),
    .Q(\tholin_riscv.tmr0[9] ),
    .D(_01513_));
 sky130_as_sc_hs__dfxtp_2 _53408_ (.CLK(clknet_leaf_168_wb_clk_i),
    .Q(\tholin_riscv.tmr0[10] ),
    .D(_01514_));
 sky130_as_sc_hs__dfxtp_2 _53409_ (.CLK(clknet_leaf_173_wb_clk_i),
    .Q(\tholin_riscv.tmr0[11] ),
    .D(_01515_));
 sky130_as_sc_hs__dfxtp_2 _53410_ (.CLK(clknet_leaf_173_wb_clk_i),
    .Q(\tholin_riscv.tmr0[12] ),
    .D(_01516_));
 sky130_as_sc_hs__dfxtp_2 _53411_ (.CLK(clknet_leaf_172_wb_clk_i),
    .Q(\tholin_riscv.tmr0[13] ),
    .D(_01517_));
 sky130_as_sc_hs__dfxtp_2 _53412_ (.CLK(clknet_leaf_174_wb_clk_i),
    .Q(\tholin_riscv.tmr0[14] ),
    .D(_01518_));
 sky130_as_sc_hs__dfxtp_2 _53413_ (.CLK(clknet_leaf_174_wb_clk_i),
    .Q(\tholin_riscv.tmr0[15] ),
    .D(_01519_));
 sky130_as_sc_hs__dfxtp_2 _53414_ (.CLK(clknet_leaf_172_wb_clk_i),
    .Q(\tholin_riscv.tmr0[16] ),
    .D(net879));
 sky130_as_sc_hs__dfxtp_2 _53415_ (.CLK(clknet_leaf_174_wb_clk_i),
    .Q(\tholin_riscv.tmr0[17] ),
    .D(_01521_));
 sky130_as_sc_hs__dfxtp_2 _53416_ (.CLK(clknet_leaf_172_wb_clk_i),
    .Q(\tholin_riscv.tmr0[18] ),
    .D(_01522_));
 sky130_as_sc_hs__dfxtp_2 _53417_ (.CLK(clknet_leaf_172_wb_clk_i),
    .Q(\tholin_riscv.tmr0[19] ),
    .D(_01523_));
 sky130_as_sc_hs__dfxtp_2 _53418_ (.CLK(clknet_leaf_177_wb_clk_i),
    .Q(\tholin_riscv.tmr0[20] ),
    .D(_01524_));
 sky130_as_sc_hs__dfxtp_2 _53419_ (.CLK(clknet_leaf_177_wb_clk_i),
    .Q(\tholin_riscv.tmr0[21] ),
    .D(_01525_));
 sky130_as_sc_hs__dfxtp_2 _53420_ (.CLK(clknet_leaf_173_wb_clk_i),
    .Q(\tholin_riscv.tmr0[22] ),
    .D(net975));
 sky130_as_sc_hs__dfxtp_2 _53421_ (.CLK(clknet_leaf_173_wb_clk_i),
    .Q(\tholin_riscv.tmr0[23] ),
    .D(_01527_));
 sky130_as_sc_hs__dfxtp_2 _53422_ (.CLK(clknet_leaf_173_wb_clk_i),
    .Q(\tholin_riscv.tmr0[24] ),
    .D(_01528_));
 sky130_as_sc_hs__dfxtp_2 _53423_ (.CLK(clknet_leaf_173_wb_clk_i),
    .Q(\tholin_riscv.tmr0[25] ),
    .D(_01529_));
 sky130_as_sc_hs__dfxtp_2 _53424_ (.CLK(clknet_leaf_178_wb_clk_i),
    .Q(\tholin_riscv.tmr0[26] ),
    .D(_01530_));
 sky130_as_sc_hs__dfxtp_2 _53425_ (.CLK(clknet_leaf_178_wb_clk_i),
    .Q(\tholin_riscv.tmr0[27] ),
    .D(_01531_));
 sky130_as_sc_hs__dfxtp_2 _53426_ (.CLK(clknet_leaf_177_wb_clk_i),
    .Q(\tholin_riscv.tmr0[28] ),
    .D(_01532_));
 sky130_as_sc_hs__dfxtp_2 _53427_ (.CLK(clknet_leaf_182_wb_clk_i),
    .Q(\tholin_riscv.tmr0[29] ),
    .D(_01533_));
 sky130_as_sc_hs__dfxtp_2 _53428_ (.CLK(clknet_leaf_182_wb_clk_i),
    .Q(\tholin_riscv.tmr0[30] ),
    .D(_01534_));
 sky130_as_sc_hs__dfxtp_2 _53429_ (.CLK(clknet_leaf_182_wb_clk_i),
    .Q(\tholin_riscv.tmr0[31] ),
    .D(_01535_));
 sky130_as_sc_hs__dfxtp_2 _53430_ (.CLK(clknet_leaf_195_wb_clk_i),
    .Q(\tholin_riscv.PCE[0] ),
    .D(_01536_));
 sky130_as_sc_hs__dfxtp_2 _53431_ (.CLK(clknet_leaf_198_wb_clk_i),
    .Q(\tholin_riscv.PCE[1] ),
    .D(_01537_));
 sky130_as_sc_hs__dfxtp_2 _53432_ (.CLK(clknet_leaf_101_wb_clk_i),
    .Q(\tholin_riscv.PCE[2] ),
    .D(_01538_));
 sky130_as_sc_hs__dfxtp_2 _53433_ (.CLK(clknet_leaf_147_wb_clk_i),
    .Q(\tholin_riscv.PCE[3] ),
    .D(_01539_));
 sky130_as_sc_hs__dfxtp_2 _53434_ (.CLK(clknet_leaf_151_wb_clk_i),
    .Q(\tholin_riscv.PCE[4] ),
    .D(_01540_));
 sky130_as_sc_hs__dfxtp_2 _53435_ (.CLK(clknet_leaf_199_wb_clk_i),
    .Q(\tholin_riscv.PCE[5] ),
    .D(_01541_));
 sky130_as_sc_hs__dfxtp_2 _53436_ (.CLK(clknet_leaf_122_wb_clk_i),
    .Q(\tholin_riscv.PCE[6] ),
    .D(_01542_));
 sky130_as_sc_hs__dfxtp_2 _53437_ (.CLK(clknet_leaf_114_wb_clk_i),
    .Q(\tholin_riscv.PCE[7] ),
    .D(_01543_));
 sky130_as_sc_hs__dfxtp_2 _53438_ (.CLK(clknet_leaf_156_wb_clk_i),
    .Q(\tholin_riscv.PCE[8] ),
    .D(_01544_));
 sky130_as_sc_hs__dfxtp_2 _53439_ (.CLK(clknet_leaf_199_wb_clk_i),
    .Q(\tholin_riscv.PCE[9] ),
    .D(_01545_));
 sky130_as_sc_hs__dfxtp_2 _53440_ (.CLK(clknet_leaf_148_wb_clk_i),
    .Q(\tholin_riscv.PCE[10] ),
    .D(_01546_));
 sky130_as_sc_hs__dfxtp_2 _53441_ (.CLK(clknet_leaf_124_wb_clk_i),
    .Q(\tholin_riscv.PCE[11] ),
    .D(_01547_));
 sky130_as_sc_hs__dfxtp_2 _53442_ (.CLK(clknet_leaf_117_wb_clk_i),
    .Q(\tholin_riscv.PCE[12] ),
    .D(_01548_));
 sky130_as_sc_hs__dfxtp_2 _53443_ (.CLK(clknet_leaf_147_wb_clk_i),
    .Q(\tholin_riscv.PCE[13] ),
    .D(_01549_));
 sky130_as_sc_hs__dfxtp_2 _53444_ (.CLK(clknet_leaf_148_wb_clk_i),
    .Q(\tholin_riscv.PCE[14] ),
    .D(_01550_));
 sky130_as_sc_hs__dfxtp_2 _53445_ (.CLK(clknet_leaf_126_wb_clk_i),
    .Q(\tholin_riscv.PCE[15] ),
    .D(_01551_));
 sky130_as_sc_hs__dfxtp_2 _53446_ (.CLK(clknet_leaf_102_wb_clk_i),
    .Q(\tholin_riscv.PCE[16] ),
    .D(_01552_));
 sky130_as_sc_hs__dfxtp_2 _53447_ (.CLK(clknet_leaf_148_wb_clk_i),
    .Q(\tholin_riscv.PCE[17] ),
    .D(_01553_));
 sky130_as_sc_hs__dfxtp_2 _53448_ (.CLK(clknet_leaf_150_wb_clk_i),
    .Q(\tholin_riscv.PCE[18] ),
    .D(_01554_));
 sky130_as_sc_hs__dfxtp_2 _53449_ (.CLK(clknet_leaf_120_wb_clk_i),
    .Q(\tholin_riscv.PCE[19] ),
    .D(_01555_));
 sky130_as_sc_hs__dfxtp_2 _53450_ (.CLK(clknet_leaf_117_wb_clk_i),
    .Q(\tholin_riscv.PCE[20] ),
    .D(_01556_));
 sky130_as_sc_hs__dfxtp_2 _53451_ (.CLK(clknet_leaf_99_wb_clk_i),
    .Q(\tholin_riscv.PCE[21] ),
    .D(_01557_));
 sky130_as_sc_hs__dfxtp_2 _53452_ (.CLK(clknet_leaf_106_wb_clk_i),
    .Q(\tholin_riscv.PCE[22] ),
    .D(_01558_));
 sky130_as_sc_hs__dfxtp_2 _53453_ (.CLK(clknet_leaf_118_wb_clk_i),
    .Q(\tholin_riscv.PCE[23] ),
    .D(_01559_));
 sky130_as_sc_hs__dfxtp_2 _53454_ (.CLK(clknet_leaf_148_wb_clk_i),
    .Q(\tholin_riscv.PCE[24] ),
    .D(_01560_));
 sky130_as_sc_hs__dfxtp_2 _53455_ (.CLK(clknet_leaf_139_wb_clk_i),
    .Q(\tholin_riscv.PCE[25] ),
    .D(_01561_));
 sky130_as_sc_hs__dfxtp_2 _53456_ (.CLK(clknet_leaf_110_wb_clk_i),
    .Q(\tholin_riscv.PCE[26] ),
    .D(_01562_));
 sky130_as_sc_hs__dfxtp_2 _53457_ (.CLK(clknet_leaf_148_wb_clk_i),
    .Q(\tholin_riscv.PCE[27] ),
    .D(_01563_));
 sky130_as_sc_hs__dfxtp_2 _53458_ (.CLK(clknet_leaf_98_wb_clk_i),
    .Q(\tholin_riscv.PCE[28] ),
    .D(_01564_));
 sky130_as_sc_hs__dfxtp_2 _53459_ (.CLK(clknet_leaf_117_wb_clk_i),
    .Q(\tholin_riscv.PCE[29] ),
    .D(_01565_));
 sky130_as_sc_hs__dfxtp_2 _53460_ (.CLK(clknet_leaf_120_wb_clk_i),
    .Q(\tholin_riscv.PCE[30] ),
    .D(_01566_));
 sky130_as_sc_hs__dfxtp_2 _53461_ (.CLK(clknet_leaf_147_wb_clk_i),
    .Q(\tholin_riscv.PCE[31] ),
    .D(_01567_));
 sky130_as_sc_hs__dfxtp_2 _53462_ (.CLK(clknet_leaf_187_wb_clk_i),
    .Q(\tholin_riscv.last_io_state ),
    .D(_01568_));
 sky130_as_sc_hs__dfxtp_2 _53463_ (.CLK(clknet_leaf_189_wb_clk_i),
    .Q(\tholin_riscv.current_irq[0] ),
    .D(net604));
 sky130_as_sc_hs__dfxtp_2 _53464_ (.CLK(clknet_leaf_110_wb_clk_i),
    .Q(\tholin_riscv.current_irq[1] ),
    .D(_01570_));
 sky130_as_sc_hs__dfxtp_2 _53465_ (.CLK(clknet_leaf_188_wb_clk_i),
    .Q(\tholin_riscv.irqs[0] ),
    .D(net550));
 sky130_as_sc_hs__dfxtp_2 _53466_ (.CLK(clknet_leaf_181_wb_clk_i),
    .Q(\tholin_riscv.irqs[1] ),
    .D(net553));
 sky130_as_sc_hs__dfxtp_2 _53467_ (.CLK(clknet_leaf_188_wb_clk_i),
    .Q(\tholin_riscv.irqs[2] ),
    .D(net1720));
 sky130_as_sc_hs__dfxtp_2 _53468_ (.CLK(clknet_leaf_181_wb_clk_i),
    .Q(\tholin_riscv.timer_int_enable ),
    .D(_01574_));
 sky130_as_sc_hs__dfxtp_2 _53469_ (.CLK(clknet_leaf_188_wb_clk_i),
    .Q(\tholin_riscv.uart_int_enable ),
    .D(_01575_));
 sky130_as_sc_hs__dfxtp_2 _53470_ (.CLK(clknet_leaf_188_wb_clk_i),
    .Q(\tholin_riscv.io_int_enable ),
    .D(_01576_));
 sky130_as_sc_hs__dfxtp_2 _53471_ (.CLK(clknet_leaf_160_wb_clk_i),
    .Q(net60),
    .D(_01577_));
 sky130_as_sc_hs__dfxtp_2 _53472_ (.CLK(clknet_leaf_160_wb_clk_i),
    .Q(net61),
    .D(_01578_));
 sky130_as_sc_hs__dfxtp_2 _53473_ (.CLK(clknet_leaf_159_wb_clk_i),
    .Q(net62),
    .D(_01579_));
 sky130_as_sc_hs__dfxtp_2 _53474_ (.CLK(clknet_leaf_159_wb_clk_i),
    .Q(net64),
    .D(_01580_));
 sky130_as_sc_hs__dfxtp_2 _53475_ (.CLK(clknet_leaf_159_wb_clk_i),
    .Q(net65),
    .D(_01581_));
 sky130_as_sc_hs__dfxtp_2 _53476_ (.CLK(clknet_leaf_159_wb_clk_i),
    .Q(net66),
    .D(_01582_));
 sky130_as_sc_hs__dfxtp_2 _53477_ (.CLK(clknet_leaf_146_wb_clk_i),
    .Q(\tholin_riscv.PORT_dir[0] ),
    .D(_01583_));
 sky130_as_sc_hs__dfxtp_2 _53478_ (.CLK(clknet_leaf_146_wb_clk_i),
    .Q(\tholin_riscv.PORT_dir[1] ),
    .D(_01584_));
 sky130_as_sc_hs__dfxtp_2 _53479_ (.CLK(clknet_leaf_96_wb_clk_i),
    .Q(\tholin_riscv.PORT_dir[2] ),
    .D(_01585_));
 sky130_as_sc_hs__dfxtp_2 _53480_ (.CLK(clknet_leaf_96_wb_clk_i),
    .Q(\tholin_riscv.PORT_dir[3] ),
    .D(_01586_));
 sky130_as_sc_hs__dfxtp_2 _53481_ (.CLK(clknet_leaf_96_wb_clk_i),
    .Q(\tholin_riscv.PORT_dir[4] ),
    .D(_01587_));
 sky130_as_sc_hs__dfxtp_2 _53482_ (.CLK(clknet_leaf_96_wb_clk_i),
    .Q(\tholin_riscv.PORT_dir[5] ),
    .D(_01588_));
 sky130_as_sc_hs__dfxtp_2 _53483_ (.CLK(clknet_leaf_130_wb_clk_i),
    .Q(\tholin_riscv.regs[9][0] ),
    .D(net680));
 sky130_as_sc_hs__dfxtp_2 _53484_ (.CLK(clknet_leaf_128_wb_clk_i),
    .Q(\tholin_riscv.regs[9][1] ),
    .D(_01590_));
 sky130_as_sc_hs__dfxtp_2 _53485_ (.CLK(clknet_leaf_64_wb_clk_i),
    .Q(\tholin_riscv.regs[9][2] ),
    .D(_01591_));
 sky130_as_sc_hs__dfxtp_2 _53486_ (.CLK(clknet_leaf_55_wb_clk_i),
    .Q(\tholin_riscv.regs[9][3] ),
    .D(_01592_));
 sky130_as_sc_hs__dfxtp_2 _53487_ (.CLK(clknet_leaf_104_wb_clk_i),
    .Q(\tholin_riscv.regs[9][4] ),
    .D(_01593_));
 sky130_as_sc_hs__dfxtp_2 _53488_ (.CLK(clknet_leaf_60_wb_clk_i),
    .Q(\tholin_riscv.regs[9][5] ),
    .D(_01594_));
 sky130_as_sc_hs__dfxtp_2 _53489_ (.CLK(clknet_leaf_61_wb_clk_i),
    .Q(\tholin_riscv.regs[9][6] ),
    .D(_01595_));
 sky130_as_sc_hs__dfxtp_2 _53490_ (.CLK(clknet_leaf_51_wb_clk_i),
    .Q(\tholin_riscv.regs[9][7] ),
    .D(_01596_));
 sky130_as_sc_hs__dfxtp_2 _53491_ (.CLK(clknet_leaf_83_wb_clk_i),
    .Q(\tholin_riscv.regs[9][8] ),
    .D(_01597_));
 sky130_as_sc_hs__dfxtp_2 _53492_ (.CLK(clknet_leaf_44_wb_clk_i),
    .Q(\tholin_riscv.regs[9][9] ),
    .D(_01598_));
 sky130_as_sc_hs__dfxtp_2 _53493_ (.CLK(clknet_leaf_48_wb_clk_i),
    .Q(\tholin_riscv.regs[9][10] ),
    .D(_01599_));
 sky130_as_sc_hs__dfxtp_2 _53494_ (.CLK(clknet_leaf_31_wb_clk_i),
    .Q(\tholin_riscv.regs[9][11] ),
    .D(_01600_));
 sky130_as_sc_hs__dfxtp_2 _53495_ (.CLK(clknet_leaf_32_wb_clk_i),
    .Q(\tholin_riscv.regs[9][12] ),
    .D(_01601_));
 sky130_as_sc_hs__dfxtp_2 _53496_ (.CLK(clknet_leaf_25_wb_clk_i),
    .Q(\tholin_riscv.regs[9][13] ),
    .D(_01602_));
 sky130_as_sc_hs__dfxtp_2 _53497_ (.CLK(clknet_leaf_14_wb_clk_i),
    .Q(\tholin_riscv.regs[9][14] ),
    .D(_01603_));
 sky130_as_sc_hs__dfxtp_2 _53498_ (.CLK(clknet_leaf_16_wb_clk_i),
    .Q(\tholin_riscv.regs[9][15] ),
    .D(_01604_));
 sky130_as_sc_hs__dfxtp_2 _53499_ (.CLK(clknet_leaf_145_wb_clk_i),
    .Q(\tholin_riscv.regs[9][16] ),
    .D(_01605_));
 sky130_as_sc_hs__dfxtp_2 _53500_ (.CLK(clknet_leaf_115_wb_clk_i),
    .Q(\tholin_riscv.regs[9][17] ),
    .D(_01606_));
 sky130_as_sc_hs__dfxtp_2 _53501_ (.CLK(clknet_leaf_118_wb_clk_i),
    .Q(\tholin_riscv.regs[9][18] ),
    .D(_01607_));
 sky130_as_sc_hs__dfxtp_2 _53502_ (.CLK(clknet_leaf_106_wb_clk_i),
    .Q(\tholin_riscv.regs[9][19] ),
    .D(_01608_));
 sky130_as_sc_hs__dfxtp_2 _53503_ (.CLK(clknet_leaf_105_wb_clk_i),
    .Q(\tholin_riscv.regs[9][20] ),
    .D(_01609_));
 sky130_as_sc_hs__dfxtp_2 _53504_ (.CLK(clknet_leaf_113_wb_clk_i),
    .Q(\tholin_riscv.regs[9][21] ),
    .D(_01610_));
 sky130_as_sc_hs__dfxtp_2 _53505_ (.CLK(clknet_leaf_104_wb_clk_i),
    .Q(\tholin_riscv.regs[9][22] ),
    .D(_01611_));
 sky130_as_sc_hs__dfxtp_2 _53506_ (.CLK(clknet_leaf_94_wb_clk_i),
    .Q(\tholin_riscv.regs[9][23] ),
    .D(_01612_));
 sky130_as_sc_hs__dfxtp_2 _53507_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[9][24] ),
    .D(_01613_));
 sky130_as_sc_hs__dfxtp_2 _53508_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[9][25] ),
    .D(_01614_));
 sky130_as_sc_hs__dfxtp_2 _53509_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[9][26] ),
    .D(_01615_));
 sky130_as_sc_hs__dfxtp_2 _53510_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[9][27] ),
    .D(_01616_));
 sky130_as_sc_hs__dfxtp_2 _53511_ (.CLK(clknet_leaf_23_wb_clk_i),
    .Q(\tholin_riscv.regs[9][28] ),
    .D(_01617_));
 sky130_as_sc_hs__dfxtp_2 _53512_ (.CLK(clknet_leaf_35_wb_clk_i),
    .Q(\tholin_riscv.regs[9][29] ),
    .D(_01618_));
 sky130_as_sc_hs__dfxtp_2 _53513_ (.CLK(clknet_leaf_96_wb_clk_i),
    .Q(\tholin_riscv.regs[9][30] ),
    .D(_01619_));
 sky130_as_sc_hs__dfxtp_2 _53514_ (.CLK(clknet_leaf_147_wb_clk_i),
    .Q(\tholin_riscv.regs[9][31] ),
    .D(_01620_));
 sky130_as_sc_hs__dfxtp_2 _53515_ (.CLK(clknet_leaf_180_wb_clk_i),
    .Q(\tholin_riscv.mul_delay ),
    .D(net598));
 sky130_as_sc_hs__dfxtp_2 _53516_ (.CLK(clknet_leaf_130_wb_clk_i),
    .Q(\tholin_riscv.regs[1][0] ),
    .D(net725));
 sky130_as_sc_hs__dfxtp_2 _53517_ (.CLK(clknet_leaf_128_wb_clk_i),
    .Q(\tholin_riscv.regs[1][1] ),
    .D(_01623_));
 sky130_as_sc_hs__dfxtp_2 _53518_ (.CLK(clknet_leaf_66_wb_clk_i),
    .Q(\tholin_riscv.regs[1][2] ),
    .D(_01624_));
 sky130_as_sc_hs__dfxtp_2 _53519_ (.CLK(clknet_leaf_13_wb_clk_i),
    .Q(\tholin_riscv.regs[1][3] ),
    .D(_01625_));
 sky130_as_sc_hs__dfxtp_2 _53520_ (.CLK(clknet_leaf_184_wb_clk_i),
    .Q(\tholin_riscv.regs[1][4] ),
    .D(_01626_));
 sky130_as_sc_hs__dfxtp_2 _53521_ (.CLK(clknet_leaf_58_wb_clk_i),
    .Q(\tholin_riscv.regs[1][5] ),
    .D(_01627_));
 sky130_as_sc_hs__dfxtp_2 _53522_ (.CLK(clknet_leaf_60_wb_clk_i),
    .Q(\tholin_riscv.regs[1][6] ),
    .D(_01628_));
 sky130_as_sc_hs__dfxtp_2 _53523_ (.CLK(clknet_leaf_50_wb_clk_i),
    .Q(\tholin_riscv.regs[1][7] ),
    .D(_01629_));
 sky130_as_sc_hs__dfxtp_2 _53524_ (.CLK(clknet_leaf_83_wb_clk_i),
    .Q(\tholin_riscv.regs[1][8] ),
    .D(_01630_));
 sky130_as_sc_hs__dfxtp_2 _53525_ (.CLK(clknet_leaf_44_wb_clk_i),
    .Q(\tholin_riscv.regs[1][9] ),
    .D(_01631_));
 sky130_as_sc_hs__dfxtp_2 _53526_ (.CLK(clknet_leaf_47_wb_clk_i),
    .Q(\tholin_riscv.regs[1][10] ),
    .D(_01632_));
 sky130_as_sc_hs__dfxtp_2 _53527_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[1][11] ),
    .D(_01633_));
 sky130_as_sc_hs__dfxtp_2 _53528_ (.CLK(clknet_leaf_37_wb_clk_i),
    .Q(\tholin_riscv.regs[1][12] ),
    .D(_01634_));
 sky130_as_sc_hs__dfxtp_2 _53529_ (.CLK(clknet_leaf_33_wb_clk_i),
    .Q(\tholin_riscv.regs[1][13] ),
    .D(_01635_));
 sky130_as_sc_hs__dfxtp_2 _53530_ (.CLK(clknet_leaf_12_wb_clk_i),
    .Q(\tholin_riscv.regs[1][14] ),
    .D(_01636_));
 sky130_as_sc_hs__dfxtp_2 _53531_ (.CLK(clknet_leaf_14_wb_clk_i),
    .Q(\tholin_riscv.regs[1][15] ),
    .D(_01637_));
 sky130_as_sc_hs__dfxtp_2 _53532_ (.CLK(clknet_leaf_115_wb_clk_i),
    .Q(\tholin_riscv.regs[1][16] ),
    .D(_01638_));
 sky130_as_sc_hs__dfxtp_2 _53533_ (.CLK(clknet_leaf_103_wb_clk_i),
    .Q(\tholin_riscv.regs[1][17] ),
    .D(_01639_));
 sky130_as_sc_hs__dfxtp_2 _53534_ (.CLK(clknet_leaf_77_wb_clk_i),
    .Q(\tholin_riscv.regs[1][18] ),
    .D(_01640_));
 sky130_as_sc_hs__dfxtp_2 _53535_ (.CLK(clknet_leaf_105_wb_clk_i),
    .Q(\tholin_riscv.regs[1][19] ),
    .D(_01641_));
 sky130_as_sc_hs__dfxtp_2 _53536_ (.CLK(clknet_leaf_114_wb_clk_i),
    .Q(\tholin_riscv.regs[1][20] ),
    .D(_01642_));
 sky130_as_sc_hs__dfxtp_2 _53537_ (.CLK(clknet_leaf_116_wb_clk_i),
    .Q(\tholin_riscv.regs[1][21] ),
    .D(_01643_));
 sky130_as_sc_hs__dfxtp_2 _53538_ (.CLK(clknet_leaf_113_wb_clk_i),
    .Q(\tholin_riscv.regs[1][22] ),
    .D(_01644_));
 sky130_as_sc_hs__dfxtp_2 _53539_ (.CLK(clknet_leaf_117_wb_clk_i),
    .Q(\tholin_riscv.regs[1][23] ),
    .D(_01645_));
 sky130_as_sc_hs__dfxtp_2 _53540_ (.CLK(clknet_leaf_34_wb_clk_i),
    .Q(\tholin_riscv.regs[1][24] ),
    .D(_01646_));
 sky130_as_sc_hs__dfxtp_2 _53541_ (.CLK(clknet_leaf_20_wb_clk_i),
    .Q(\tholin_riscv.regs[1][25] ),
    .D(_01647_));
 sky130_as_sc_hs__dfxtp_2 _53542_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[1][26] ),
    .D(_01648_));
 sky130_as_sc_hs__dfxtp_2 _53543_ (.CLK(clknet_leaf_25_wb_clk_i),
    .Q(\tholin_riscv.regs[1][27] ),
    .D(_01649_));
 sky130_as_sc_hs__dfxtp_2 _53544_ (.CLK(clknet_leaf_24_wb_clk_i),
    .Q(\tholin_riscv.regs[1][28] ),
    .D(_01650_));
 sky130_as_sc_hs__dfxtp_2 _53545_ (.CLK(clknet_leaf_36_wb_clk_i),
    .Q(\tholin_riscv.regs[1][29] ),
    .D(_01651_));
 sky130_as_sc_hs__dfxtp_2 _53546_ (.CLK(clknet_leaf_117_wb_clk_i),
    .Q(\tholin_riscv.regs[1][30] ),
    .D(_01652_));
 sky130_as_sc_hs__dfxtp_2 _53547_ (.CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\tholin_riscv.regs[1][31] ),
    .D(_01653_));
 sky130_as_sc_hs__dfxtp_2 _53548_ (.CLK(clknet_leaf_197_wb_clk_i),
    .Q(\tholin_riscv.PC[2] ),
    .D(_01654_));
 sky130_as_sc_hs__dfxtp_2 _53549_ (.CLK(clknet_leaf_197_wb_clk_i),
    .Q(\tholin_riscv.PC[3] ),
    .D(_01655_));
 sky130_as_sc_hs__dfxtp_2 _53550_ (.CLK(clknet_leaf_197_wb_clk_i),
    .Q(\tholin_riscv.PC[4] ),
    .D(_01656_));
 sky130_as_sc_hs__dfxtp_2 _53551_ (.CLK(clknet_leaf_197_wb_clk_i),
    .Q(\tholin_riscv.PC[5] ),
    .D(_01657_));
 sky130_as_sc_hs__dfxtp_2 _53552_ (.CLK(clknet_leaf_197_wb_clk_i),
    .Q(\tholin_riscv.PC[6] ),
    .D(_01658_));
 sky130_as_sc_hs__dfxtp_2 _53553_ (.CLK(clknet_leaf_197_wb_clk_i),
    .Q(\tholin_riscv.PC[7] ),
    .D(_01659_));
 sky130_as_sc_hs__dfxtp_2 _53554_ (.CLK(clknet_leaf_197_wb_clk_i),
    .Q(\tholin_riscv.PC[8] ),
    .D(_01660_));
 sky130_as_sc_hs__dfxtp_2 _53555_ (.CLK(clknet_leaf_199_wb_clk_i),
    .Q(\tholin_riscv.PC[9] ),
    .D(_01661_));
 sky130_as_sc_hs__dfxtp_2 _53556_ (.CLK(clknet_leaf_199_wb_clk_i),
    .Q(\tholin_riscv.PC[10] ),
    .D(_01662_));
 sky130_as_sc_hs__dfxtp_2 _53557_ (.CLK(clknet_leaf_198_wb_clk_i),
    .Q(\tholin_riscv.PC[11] ),
    .D(_01663_));
 sky130_as_sc_hs__dfxtp_2 _53558_ (.CLK(clknet_leaf_202_wb_clk_i),
    .Q(\tholin_riscv.PC[12] ),
    .D(_01664_));
 sky130_as_sc_hs__dfxtp_2 _53559_ (.CLK(clknet_leaf_198_wb_clk_i),
    .Q(\tholin_riscv.PC[13] ),
    .D(_01665_));
 sky130_as_sc_hs__dfxtp_2 _53560_ (.CLK(clknet_leaf_198_wb_clk_i),
    .Q(\tholin_riscv.PC[14] ),
    .D(_01666_));
 sky130_as_sc_hs__dfxtp_2 _53561_ (.CLK(clknet_leaf_197_wb_clk_i),
    .Q(\tholin_riscv.PC[15] ),
    .D(_01667_));
 sky130_as_sc_hs__dfxtp_2 _53562_ (.CLK(clknet_leaf_4_wb_clk_i),
    .Q(\tholin_riscv.PC[16] ),
    .D(_01668_));
 sky130_as_sc_hs__dfxtp_2 _53563_ (.CLK(clknet_leaf_4_wb_clk_i),
    .Q(\tholin_riscv.PC[17] ),
    .D(_01669_));
 sky130_as_sc_hs__dfxtp_2 _53564_ (.CLK(clknet_leaf_5_wb_clk_i),
    .Q(\tholin_riscv.PC[18] ),
    .D(_01670_));
 sky130_as_sc_hs__dfxtp_2 _53565_ (.CLK(clknet_leaf_5_wb_clk_i),
    .Q(\tholin_riscv.PC[19] ),
    .D(_01671_));
 sky130_as_sc_hs__dfxtp_2 _53566_ (.CLK(clknet_leaf_5_wb_clk_i),
    .Q(\tholin_riscv.PC[20] ),
    .D(_01672_));
 sky130_as_sc_hs__dfxtp_2 _53567_ (.CLK(clknet_leaf_196_wb_clk_i),
    .Q(\tholin_riscv.PC[21] ),
    .D(_01673_));
 sky130_as_sc_hs__dfxtp_2 _53568_ (.CLK(clknet_leaf_196_wb_clk_i),
    .Q(\tholin_riscv.PC[22] ),
    .D(_01674_));
 sky130_as_sc_hs__dfxtp_2 _53569_ (.CLK(clknet_leaf_196_wb_clk_i),
    .Q(\tholin_riscv.PC[23] ),
    .D(_01675_));
 sky130_as_sc_hs__dfxtp_2 _53570_ (.CLK(clknet_leaf_195_wb_clk_i),
    .Q(\tholin_riscv.PC[24] ),
    .D(_01676_));
 sky130_as_sc_hs__dfxtp_2 _53571_ (.CLK(clknet_leaf_195_wb_clk_i),
    .Q(\tholin_riscv.PC[25] ),
    .D(_01677_));
 sky130_as_sc_hs__dfxtp_2 _53572_ (.CLK(clknet_leaf_194_wb_clk_i),
    .Q(\tholin_riscv.PC[26] ),
    .D(_01678_));
 sky130_as_sc_hs__dfxtp_2 _53573_ (.CLK(clknet_leaf_194_wb_clk_i),
    .Q(\tholin_riscv.PC[27] ),
    .D(_01679_));
 sky130_as_sc_hs__dfxtp_2 _53574_ (.CLK(clknet_leaf_194_wb_clk_i),
    .Q(\tholin_riscv.PC[28] ),
    .D(_01680_));
 sky130_as_sc_hs__dfxtp_2 _53575_ (.CLK(clknet_leaf_194_wb_clk_i),
    .Q(\tholin_riscv.PC[29] ),
    .D(_01681_));
 sky130_as_sc_hs__dfxtp_2 _53576_ (.CLK(clknet_leaf_191_wb_clk_i),
    .Q(\tholin_riscv.PC[30] ),
    .D(_01682_));
 sky130_as_sc_hs__dfxtp_2 _53577_ (.CLK(clknet_leaf_191_wb_clk_i),
    .Q(\tholin_riscv.PC[31] ),
    .D(_01683_));
 sky130_as_sc_hs__dfxtp_2 _53578_ (.CLK(clknet_leaf_133_wb_clk_i),
    .Q(_00000_),
    .D(_01684_));
 sky130_as_sc_hs__dfxtp_2 _53579_ (.CLK(clknet_leaf_5_wb_clk_i),
    .Q(_00001_),
    .D(_01685_));
 sky130_as_sc_hs__dfxtp_2 _53580_ (.CLK(clknet_leaf_135_wb_clk_i),
    .Q(_00002_),
    .D(_01686_));
 sky130_as_sc_hs__dfxtp_2 _53581_ (.CLK(clknet_leaf_6_wb_clk_i),
    .Q(_00003_),
    .D(_01687_));
 sky130_as_sc_hs__dfxtp_2 _53582_ (.CLK(clknet_leaf_6_wb_clk_i),
    .Q(_00004_),
    .D(_01688_));
 sky130_as_sc_hs__dfxtp_2 _53583_ (.CLK(clknet_leaf_131_wb_clk_i),
    .Q(\tholin_riscv.regs[29][0] ),
    .D(net671));
 sky130_as_sc_hs__dfxtp_2 _53584_ (.CLK(clknet_leaf_126_wb_clk_i),
    .Q(\tholin_riscv.regs[29][1] ),
    .D(_01690_));
 sky130_as_sc_hs__dfxtp_2 _53585_ (.CLK(clknet_leaf_63_wb_clk_i),
    .Q(\tholin_riscv.regs[29][2] ),
    .D(_01691_));
 sky130_as_sc_hs__dfxtp_2 _53586_ (.CLK(clknet_leaf_55_wb_clk_i),
    .Q(\tholin_riscv.regs[29][3] ),
    .D(_01692_));
 sky130_as_sc_hs__dfxtp_2 _53587_ (.CLK(clknet_leaf_148_wb_clk_i),
    .Q(\tholin_riscv.regs[29][4] ),
    .D(_01693_));
 sky130_as_sc_hs__dfxtp_2 _53588_ (.CLK(clknet_leaf_54_wb_clk_i),
    .Q(\tholin_riscv.regs[29][5] ),
    .D(_01694_));
 sky130_as_sc_hs__dfxtp_2 _53589_ (.CLK(clknet_leaf_62_wb_clk_i),
    .Q(\tholin_riscv.regs[29][6] ),
    .D(_01695_));
 sky130_as_sc_hs__dfxtp_2 _53590_ (.CLK(clknet_leaf_52_wb_clk_i),
    .Q(\tholin_riscv.regs[29][7] ),
    .D(_01696_));
 sky130_as_sc_hs__dfxtp_2 _53591_ (.CLK(clknet_leaf_80_wb_clk_i),
    .Q(\tholin_riscv.regs[29][8] ),
    .D(_01697_));
 sky130_as_sc_hs__dfxtp_2 _53592_ (.CLK(clknet_leaf_44_wb_clk_i),
    .Q(\tholin_riscv.regs[29][9] ),
    .D(_01698_));
 sky130_as_sc_hs__dfxtp_2 _53593_ (.CLK(clknet_leaf_49_wb_clk_i),
    .Q(\tholin_riscv.regs[29][10] ),
    .D(_01699_));
 sky130_as_sc_hs__dfxtp_2 _53594_ (.CLK(clknet_leaf_30_wb_clk_i),
    .Q(\tholin_riscv.regs[29][11] ),
    .D(_01700_));
 sky130_as_sc_hs__dfxtp_2 _53595_ (.CLK(clknet_leaf_26_wb_clk_i),
    .Q(\tholin_riscv.regs[29][12] ),
    .D(_01701_));
 sky130_as_sc_hs__dfxtp_2 _53596_ (.CLK(clknet_leaf_28_wb_clk_i),
    .Q(\tholin_riscv.regs[29][13] ),
    .D(_01702_));
 sky130_as_sc_hs__dfxtp_2 _53597_ (.CLK(clknet_leaf_19_wb_clk_i),
    .Q(\tholin_riscv.regs[29][14] ),
    .D(_01703_));
 sky130_as_sc_hs__dfxtp_2 _53598_ (.CLK(clknet_leaf_18_wb_clk_i),
    .Q(\tholin_riscv.regs[29][15] ),
    .D(_01704_));
 sky130_as_sc_hs__dfxtp_2 _53599_ (.CLK(clknet_leaf_108_wb_clk_i),
    .Q(\tholin_riscv.regs[29][16] ),
    .D(_01705_));
 sky130_as_sc_hs__dfxtp_2 _53600_ (.CLK(clknet_leaf_107_wb_clk_i),
    .Q(\tholin_riscv.regs[29][17] ),
    .D(_01706_));
 sky130_as_sc_hs__dfxtp_2 _53601_ (.CLK(clknet_leaf_103_wb_clk_i),
    .Q(\tholin_riscv.regs[29][18] ),
    .D(_01707_));
 sky130_as_sc_hs__dfxtp_2 _53602_ (.CLK(clknet_leaf_106_wb_clk_i),
    .Q(\tholin_riscv.regs[29][19] ),
    .D(_01708_));
 sky130_as_sc_hs__dfxtp_2 _53603_ (.CLK(clknet_leaf_117_wb_clk_i),
    .Q(\tholin_riscv.regs[29][20] ),
    .D(_01709_));
 sky130_as_sc_hs__dfxtp_2 _53604_ (.CLK(clknet_leaf_106_wb_clk_i),
    .Q(\tholin_riscv.regs[29][21] ),
    .D(_01710_));
 sky130_as_sc_hs__dfxtp_2 _53605_ (.CLK(clknet_leaf_102_wb_clk_i),
    .Q(\tholin_riscv.regs[29][22] ),
    .D(_01711_));
 sky130_as_sc_hs__dfxtp_2 _53606_ (.CLK(clknet_leaf_114_wb_clk_i),
    .Q(\tholin_riscv.regs[29][23] ),
    .D(_01712_));
 sky130_as_sc_hs__dfxtp_2 _53607_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[29][24] ),
    .D(_01713_));
 sky130_as_sc_hs__dfxtp_2 _53608_ (.CLK(clknet_leaf_79_wb_clk_i),
    .Q(\tholin_riscv.regs[29][25] ),
    .D(_01714_));
 sky130_as_sc_hs__dfxtp_2 _53609_ (.CLK(clknet_leaf_87_wb_clk_i),
    .Q(\tholin_riscv.regs[29][26] ),
    .D(_01715_));
 sky130_as_sc_hs__dfxtp_2 _53610_ (.CLK(clknet_leaf_92_wb_clk_i),
    .Q(\tholin_riscv.regs[29][27] ),
    .D(_01716_));
 sky130_as_sc_hs__dfxtp_2 _53611_ (.CLK(clknet_leaf_90_wb_clk_i),
    .Q(\tholin_riscv.regs[29][28] ),
    .D(_01717_));
 sky130_as_sc_hs__dfxtp_2 _53612_ (.CLK(clknet_leaf_40_wb_clk_i),
    .Q(\tholin_riscv.regs[29][29] ),
    .D(_01718_));
 sky130_as_sc_hs__dfxtp_2 _53613_ (.CLK(clknet_leaf_124_wb_clk_i),
    .Q(\tholin_riscv.regs[29][30] ),
    .D(_01719_));
 sky130_as_sc_hs__dfxtp_2 _53614_ (.CLK(clknet_leaf_134_wb_clk_i),
    .Q(\tholin_riscv.regs[29][31] ),
    .D(_01720_));
 sky130_as_sc_hs__buff_2 _53629_ (.A(net124),
    .Y(net23));
 sky130_as_sc_hs__buff_2 _53630_ (.A(net124),
    .Y(net30));
 sky130_as_sc_hs__buff_2 _53631_ (.A(net124),
    .Y(net34));
 sky130_as_sc_hs__buff_2 _53632_ (.A(net124),
    .Y(net38));
 sky130_as_sc_hs__buff_2 _53633_ (.A(net124),
    .Y(net39));
 sky130_as_sc_hs__buff_2 _53634_ (.A(net124),
    .Y(net40));
 sky130_as_sc_hs__buff_2 _53635_ (.A(net124),
    .Y(net41));
 sky130_as_sc_hs__buff_2 _53636_ (.A(net124),
    .Y(net42));
 sky130_as_sc_hs__buff_2 _53637_ (.A(net124),
    .Y(net43));
 sky130_as_sc_hs__buff_2 _53638_ (.A(net124),
    .Y(net44));
 sky130_as_sc_hs__buff_2 _53639_ (.A(net124),
    .Y(net24));
 sky130_as_sc_hs__buff_2 _53640_ (.A(net124),
    .Y(net25));
 sky130_as_sc_hs__buff_2 _53641_ (.A(net124),
    .Y(net26));
 sky130_as_sc_hs__buff_2 _53642_ (.A(net124),
    .Y(net27));
 sky130_as_sc_hs__buff_2 _53643_ (.A(net124),
    .Y(net28));
 sky130_as_sc_hs__buff_2 _53644_ (.A(net124),
    .Y(net54));
 sky130_as_sc_hs__clkbuff_11 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .Y(clknet_0_wb_clk_i));
 sky130_as_sc_hs__clkbuff_8 clkbuf_2_0_0_wb_clk_i (.Y(clknet_2_0_0_wb_clk_i),
    .A(clknet_0_wb_clk_i));
 sky130_as_sc_hs__clkbuff_8 clkbuf_2_1_0_wb_clk_i (.Y(clknet_2_1_0_wb_clk_i),
    .A(clknet_0_wb_clk_i));
 sky130_as_sc_hs__clkbuff_8 clkbuf_2_2_0_wb_clk_i (.Y(clknet_2_2_0_wb_clk_i),
    .A(clknet_0_wb_clk_i));
 sky130_as_sc_hs__clkbuff_8 clkbuf_2_3_0_wb_clk_i (.Y(clknet_2_3_0_wb_clk_i),
    .A(clknet_0_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_0__f_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .Y(clknet_4_0__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_10__f_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .Y(clknet_4_10__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_11__f_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .Y(clknet_4_11__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_12__f_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .Y(clknet_4_12__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_13__f_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .Y(clknet_4_13__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_14__f_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .Y(clknet_4_14__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_15__f_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .Y(clknet_4_15__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_1__f_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .Y(clknet_4_1__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_2__f_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .Y(clknet_4_2__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_3__f_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .Y(clknet_4_3__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_4__f_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .Y(clknet_4_4__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_5__f_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .Y(clknet_4_5__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_6__f_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .Y(clknet_4_6__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_7__f_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .Y(clknet_4_7__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_8__f_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .Y(clknet_4_8__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_4_9__f_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .Y(clknet_4_9__leaf_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_100_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_100_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_101_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_101_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_102_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_102_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_103_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_103_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_104_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_104_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_105_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_105_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_106_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_106_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_107_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .Y(clknet_leaf_107_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_108_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .Y(clknet_leaf_108_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_109_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_109_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_10_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_10_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_110_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .Y(clknet_leaf_110_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_111_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .Y(clknet_leaf_111_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_112_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .Y(clknet_leaf_112_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_113_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .Y(clknet_leaf_113_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_114_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .Y(clknet_leaf_114_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_115_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_115_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_116_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_116_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_117_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .Y(clknet_leaf_117_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_118_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .Y(clknet_leaf_118_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_119_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .Y(clknet_leaf_119_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_11_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_11_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_120_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .Y(clknet_leaf_120_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_121_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .Y(clknet_leaf_121_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_122_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_122_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_123_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_123_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_124_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_124_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_125_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_125_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_126_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_126_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_127_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_127_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_128_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_128_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_129_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_129_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_12_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_12_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_130_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_130_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_131_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .Y(clknet_leaf_131_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_132_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_132_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_133_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_133_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_134_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_134_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_135_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_135_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_136_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_136_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_137_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_137_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_138_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_138_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_139_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_139_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_13_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_13_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_140_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_140_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_141_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_141_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_142_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_142_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_143_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_143_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_144_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_144_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_145_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_145_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_146_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_146_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_147_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_147_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_148_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_148_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_149_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_149_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_14_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_14_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_150_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_150_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_151_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_151_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_152_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_152_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_153_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .Y(clknet_leaf_153_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_154_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .Y(clknet_leaf_154_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_155_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .Y(clknet_leaf_155_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_156_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .Y(clknet_leaf_156_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_157_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .Y(clknet_leaf_157_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_158_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .Y(clknet_leaf_158_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_159_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .Y(clknet_leaf_159_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_15_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_15_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_160_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .Y(clknet_leaf_160_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_161_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .Y(clknet_leaf_161_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_162_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .Y(clknet_leaf_162_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_163_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .Y(clknet_leaf_163_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_164_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .Y(clknet_leaf_164_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_165_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .Y(clknet_leaf_165_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_166_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .Y(clknet_leaf_166_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_167_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .Y(clknet_leaf_167_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_168_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .Y(clknet_leaf_168_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_169_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .Y(clknet_leaf_169_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_16_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_16_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_170_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .Y(clknet_leaf_170_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_171_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .Y(clknet_leaf_171_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_172_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .Y(clknet_leaf_172_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_173_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .Y(clknet_leaf_173_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_174_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .Y(clknet_leaf_174_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_175_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .Y(clknet_leaf_175_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_176_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .Y(clknet_leaf_176_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_177_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .Y(clknet_leaf_177_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_178_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .Y(clknet_leaf_178_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_179_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .Y(clknet_leaf_179_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_17_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_17_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_180_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .Y(clknet_leaf_180_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_181_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .Y(clknet_leaf_181_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_182_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .Y(clknet_leaf_182_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_183_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .Y(clknet_leaf_183_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_184_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .Y(clknet_leaf_184_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_185_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_185_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_186_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_186_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_187_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_187_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_188_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .Y(clknet_leaf_188_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_189_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .Y(clknet_leaf_189_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_18_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_18_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_190_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .Y(clknet_leaf_190_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_191_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .Y(clknet_leaf_191_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_192_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_192_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_193_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .Y(clknet_leaf_193_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_194_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .Y(clknet_leaf_194_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_195_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .Y(clknet_leaf_195_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_196_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .Y(clknet_leaf_196_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_197_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .Y(clknet_leaf_197_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_198_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .Y(clknet_leaf_198_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_199_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .Y(clknet_leaf_199_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_19_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_19_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_1_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .Y(clknet_leaf_1_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_200_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .Y(clknet_leaf_200_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_202_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .Y(clknet_leaf_202_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_203_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .Y(clknet_leaf_203_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_204_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .Y(clknet_leaf_204_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_205_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .Y(clknet_leaf_205_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_206_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .Y(clknet_leaf_206_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_207_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .Y(clknet_leaf_207_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_208_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .Y(clknet_leaf_208_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_209_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .Y(clknet_leaf_209_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_20_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_20_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_210_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .Y(clknet_leaf_210_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_211_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .Y(clknet_leaf_211_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_212_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .Y(clknet_leaf_212_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_213_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .Y(clknet_leaf_213_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_214_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .Y(clknet_leaf_214_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_215_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .Y(clknet_leaf_215_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_216_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .Y(clknet_leaf_216_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_218_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .Y(clknet_leaf_218_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_21_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_21_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_22_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_22_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_23_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_23_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_24_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_24_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_25_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_25_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_26_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_26_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_27_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_27_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_28_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_28_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_29_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_29_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_2_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .Y(clknet_leaf_2_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_30_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_30_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_31_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_31_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_32_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_32_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_33_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_33_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_34_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_34_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_35_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_35_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_36_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_36_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_37_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_37_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_38_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_38_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_39_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_39_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_3_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .Y(clknet_leaf_3_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_40_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_40_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_41_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_41_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_42_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_42_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_43_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_43_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_44_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_44_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_45_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_45_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_46_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_46_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_47_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_47_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_48_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_48_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_49_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_49_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_4_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .Y(clknet_leaf_4_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_50_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_50_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_51_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .Y(clknet_leaf_51_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_52_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_52_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_53_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_53_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_54_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_54_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_55_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_55_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_56_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_56_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_57_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_57_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_58_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_58_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_59_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_59_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_5_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .Y(clknet_leaf_5_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_60_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_60_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_61_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_61_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_62_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_62_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_63_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_63_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_64_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_64_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_65_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_65_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_66_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_66_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_67_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_67_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_68_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_68_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_69_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_69_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_6_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_6_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_70_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_70_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_71_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_71_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_72_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_72_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_73_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_73_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_74_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_74_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_75_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .Y(clknet_leaf_75_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_77_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .Y(clknet_leaf_77_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_78_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .Y(clknet_leaf_78_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_79_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .Y(clknet_leaf_79_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_7_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_7_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_80_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .Y(clknet_leaf_80_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_81_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .Y(clknet_leaf_81_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_82_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_82_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_83_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_83_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_84_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .Y(clknet_leaf_84_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_85_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .Y(clknet_leaf_85_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_86_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_86_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_87_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .Y(clknet_leaf_87_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_88_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .Y(clknet_leaf_88_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_89_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .Y(clknet_leaf_89_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_8_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .Y(clknet_leaf_8_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_90_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .Y(clknet_leaf_90_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_91_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .Y(clknet_leaf_91_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_92_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .Y(clknet_leaf_92_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_93_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_93_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_94_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_94_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_96_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_96_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_97_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_97_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_98_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_98_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_99_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .Y(clknet_leaf_99_wb_clk_i));
 sky130_as_sc_hs__clkbuff_11 clkbuf_leaf_9_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .Y(clknet_leaf_9_wb_clk_i));
 sky130_as_sc_hs__clkbuff_8 fanout100 (.Y(net100),
    .A(_15290_));
 sky130_as_sc_hs__clkbuff_11 fanout101 (.A(_15290_),
    .Y(net101));
 sky130_as_sc_hs__clkbuff_11 fanout102 (.A(_15290_),
    .Y(net102));
 sky130_as_sc_hs__clkbuff_8 fanout103 (.Y(net103),
    .A(_19961_));
 sky130_as_sc_hs__clkbuff_8 fanout104 (.Y(net104),
    .A(_19961_));
 sky130_as_sc_hs__clkbuff_8 fanout105 (.Y(net105),
    .A(net106));
 sky130_as_sc_hs__clkbuff_8 fanout106 (.Y(net106),
    .A(_19930_));
 sky130_as_sc_hs__buff_11 fanout107 (.A(net109),
    .Y(net107));
 sky130_as_sc_hs__buff_4 fanout108 (.A(net109),
    .Y(net108));
 sky130_as_sc_hs__clkbuff_8 fanout109 (.Y(net109),
    .A(_06562_));
 sky130_as_sc_hs__buff_11 fanout110 (.A(net111),
    .Y(net110));
 sky130_as_sc_hs__buff_11 fanout111 (.A(_06555_),
    .Y(net111));
 sky130_as_sc_hs__clkbuff_11 fanout112 (.A(net113),
    .Y(net112));
 sky130_as_sc_hs__buff_11 fanout113 (.A(_22167_),
    .Y(net113));
 sky130_as_sc_hs__clkbuff_8 fanout114 (.Y(net114),
    .A(net115));
 sky130_as_sc_hs__buff_4 fanout115 (.A(net116),
    .Y(net115));
 sky130_as_sc_hs__clkbuff_11 fanout116 (.A(_20825_),
    .Y(net116));
 sky130_as_sc_hs__buff_11 fanout117 (.A(_06914_),
    .Y(net117));
 sky130_as_sc_hs__buff_11 fanout118 (.A(net119),
    .Y(net118));
 sky130_as_sc_hs__buff_11 fanout119 (.A(_06523_),
    .Y(net119));
 sky130_as_sc_hs__clkbuff_11 fanout120 (.A(net121),
    .Y(net120));
 sky130_as_sc_hs__clkbuff_8 fanout121 (.Y(net121),
    .A(_23691_));
 sky130_as_sc_hs__clkbuff_11 fanout122 (.A(net123),
    .Y(net122));
 sky130_as_sc_hs__clkbuff_11 fanout123 (.A(_23534_),
    .Y(net123));
 sky130_as_sc_hs__buff_11 fanout124 (.A(net29),
    .Y(net124));
 sky130_as_sc_hs__clkbuff_11 fanout125 (.A(_13061_),
    .Y(net125));
 sky130_as_sc_hs__clkbuff_11 fanout126 (.A(net127),
    .Y(net126));
 sky130_as_sc_hs__clkbuff_11 fanout127 (.A(_05518_),
    .Y(net127));
 sky130_as_sc_hs__clkbuff_8 fanout128 (.Y(net128),
    .A(_02387_));
 sky130_as_sc_hs__clkbuff_8 fanout129 (.Y(net129),
    .A(_02387_));
 sky130_as_sc_hs__clkbuff_8 fanout130 (.Y(net130),
    .A(net131));
 sky130_as_sc_hs__buff_4 fanout131 (.A(_16428_),
    .Y(net131));
 sky130_as_sc_hs__buff_11 fanout132 (.A(net134),
    .Y(net132));
 sky130_as_sc_hs__buff_4 fanout133 (.A(net134),
    .Y(net133));
 sky130_as_sc_hs__buff_11 fanout134 (.A(_15287_),
    .Y(net134));
 sky130_as_sc_hs__buff_11 fanout135 (.A(net136),
    .Y(net135));
 sky130_as_sc_hs__buff_11 fanout136 (.A(_19989_),
    .Y(net136));
 sky130_as_sc_hs__buff_11 fanout137 (.A(_19758_),
    .Y(net137));
 sky130_as_sc_hs__buff_11 fanout138 (.A(net139),
    .Y(net138));
 sky130_as_sc_hs__buff_11 fanout139 (.A(_06163_),
    .Y(net139));
 sky130_as_sc_hs__clkbuff_8 fanout140 (.Y(net140),
    .A(_05926_));
 sky130_as_sc_hs__buff_11 fanout141 (.A(net142),
    .Y(net141));
 sky130_as_sc_hs__buff_11 fanout142 (.A(_05510_),
    .Y(net142));
 sky130_as_sc_hs__buff_11 fanout143 (.A(net144),
    .Y(net143));
 sky130_as_sc_hs__buff_11 fanout144 (.A(net145),
    .Y(net144));
 sky130_as_sc_hs__clkbuff_8 fanout145 (.Y(net145),
    .A(_19934_));
 sky130_as_sc_hs__buff_4 fanout146 (.A(net147),
    .Y(net146));
 sky130_as_sc_hs__buff_2 fanout147 (.A(net148),
    .Y(net147));
 sky130_as_sc_hs__clkbuff_4 fanout148 (.A(_18407_),
    .Y(net148));
 sky130_as_sc_hs__clkbuff_8 fanout149 (.Y(net149),
    .A(_05515_));
 sky130_as_sc_hs__buff_11 fanout150 (.A(net151),
    .Y(net150));
 sky130_as_sc_hs__buff_11 fanout151 (.A(_19538_),
    .Y(net151));
 sky130_as_sc_hs__buff_11 fanout152 (.A(net153),
    .Y(net152));
 sky130_as_sc_hs__buff_11 fanout153 (.A(net156),
    .Y(net153));
 sky130_as_sc_hs__buff_11 fanout154 (.A(net156),
    .Y(net154));
 sky130_as_sc_hs__buff_11 fanout155 (.A(net156),
    .Y(net155));
 sky130_as_sc_hs__buff_11 fanout156 (.A(_19537_),
    .Y(net156));
 sky130_as_sc_hs__buff_11 fanout157 (.A(net160),
    .Y(net157));
 sky130_as_sc_hs__buff_11 fanout158 (.A(net160),
    .Y(net158));
 sky130_as_sc_hs__buff_11 fanout159 (.A(net160),
    .Y(net159));
 sky130_as_sc_hs__buff_11 fanout160 (.A(_19536_),
    .Y(net160));
 sky130_as_sc_hs__buff_11 fanout161 (.A(net165),
    .Y(net161));
 sky130_as_sc_hs__buff_11 fanout162 (.A(net165),
    .Y(net162));
 sky130_as_sc_hs__buff_11 fanout163 (.A(net165),
    .Y(net163));
 sky130_as_sc_hs__buff_11 fanout164 (.A(net165),
    .Y(net164));
 sky130_as_sc_hs__buff_11 fanout165 (.A(_19536_),
    .Y(net165));
 sky130_as_sc_hs__buff_11 fanout166 (.A(net167),
    .Y(net166));
 sky130_as_sc_hs__buff_11 fanout167 (.A(net173),
    .Y(net167));
 sky130_as_sc_hs__buff_11 fanout168 (.A(net173),
    .Y(net168));
 sky130_as_sc_hs__clkbuff_11 fanout169 (.A(net173),
    .Y(net169));
 sky130_as_sc_hs__buff_11 fanout170 (.A(net172),
    .Y(net170));
 sky130_as_sc_hs__buff_11 fanout171 (.A(net172),
    .Y(net171));
 sky130_as_sc_hs__clkbuff_8 fanout172 (.Y(net172),
    .A(net173));
 sky130_as_sc_hs__buff_11 fanout173 (.A(_19535_),
    .Y(net173));
 sky130_as_sc_hs__buff_11 fanout174 (.A(net186),
    .Y(net174));
 sky130_as_sc_hs__clkbuff_11 fanout175 (.A(net186),
    .Y(net175));
 sky130_as_sc_hs__buff_11 fanout176 (.A(net179),
    .Y(net176));
 sky130_as_sc_hs__buff_11 fanout177 (.A(net178),
    .Y(net177));
 sky130_as_sc_hs__clkbuff_8 fanout178 (.Y(net178),
    .A(net179));
 sky130_as_sc_hs__clkbuff_8 fanout179 (.Y(net179),
    .A(net186));
 sky130_as_sc_hs__buff_11 fanout180 (.A(net186),
    .Y(net180));
 sky130_as_sc_hs__buff_4 fanout181 (.A(net182),
    .Y(net181));
 sky130_as_sc_hs__buff_11 fanout182 (.A(net186),
    .Y(net182));
 sky130_as_sc_hs__buff_11 fanout183 (.A(net186),
    .Y(net183));
 sky130_as_sc_hs__clkbuff_8 fanout184 (.Y(net184),
    .A(net186));
 sky130_as_sc_hs__buff_11 fanout185 (.A(net186),
    .Y(net185));
 sky130_as_sc_hs__buff_11 fanout186 (.A(_19535_),
    .Y(net186));
 sky130_as_sc_hs__clkbuff_8 fanout187 (.Y(net187),
    .A(net190));
 sky130_as_sc_hs__clkbuff_8 fanout188 (.Y(net188),
    .A(net190));
 sky130_as_sc_hs__buff_4 fanout189 (.A(net190),
    .Y(net189));
 sky130_as_sc_hs__buff_4 fanout190 (.A(_19534_),
    .Y(net190));
 sky130_as_sc_hs__clkbuff_8 fanout191 (.Y(net191),
    .A(net195));
 sky130_as_sc_hs__clkbuff_4 fanout192 (.A(net195),
    .Y(net192));
 sky130_as_sc_hs__clkbuff_8 fanout193 (.Y(net193),
    .A(net195));
 sky130_as_sc_hs__buff_2 fanout194 (.A(net195),
    .Y(net194));
 sky130_as_sc_hs__clkbuff_8 fanout195 (.Y(net195),
    .A(_19534_));
 sky130_as_sc_hs__clkbuff_8 fanout196 (.Y(net196),
    .A(_19534_));
 sky130_as_sc_hs__clkbuff_8 fanout197 (.Y(net197),
    .A(net198));
 sky130_as_sc_hs__clkbuff_8 fanout198 (.Y(net198),
    .A(_19534_));
 sky130_as_sc_hs__clkbuff_8 fanout199 (.Y(net199),
    .A(net200));
 sky130_as_sc_hs__clkbuff_8 fanout200 (.Y(net200),
    .A(_19534_));
 sky130_as_sc_hs__clkbuff_8 fanout201 (.Y(net201),
    .A(net210));
 sky130_as_sc_hs__buff_4 fanout202 (.A(net210),
    .Y(net202));
 sky130_as_sc_hs__clkbuff_8 fanout203 (.Y(net203),
    .A(net210));
 sky130_as_sc_hs__clkbuff_8 fanout204 (.Y(net204),
    .A(net206));
 sky130_as_sc_hs__clkbuff_8 fanout205 (.Y(net205),
    .A(net206));
 sky130_as_sc_hs__buff_4 fanout206 (.A(net210),
    .Y(net206));
 sky130_as_sc_hs__clkbuff_8 fanout207 (.Y(net207),
    .A(net208));
 sky130_as_sc_hs__clkbuff_8 fanout208 (.Y(net208),
    .A(net209));
 sky130_as_sc_hs__clkbuff_8 fanout209 (.Y(net209),
    .A(net210));
 sky130_as_sc_hs__buff_4 fanout210 (.A(_19485_),
    .Y(net210));
 sky130_as_sc_hs__buff_11 fanout211 (.A(net219),
    .Y(net211));
 sky130_as_sc_hs__buff_11 fanout212 (.A(net213),
    .Y(net212));
 sky130_as_sc_hs__buff_11 fanout213 (.A(net214),
    .Y(net213));
 sky130_as_sc_hs__buff_11 fanout214 (.A(net219),
    .Y(net214));
 sky130_as_sc_hs__buff_11 fanout215 (.A(net219),
    .Y(net215));
 sky130_as_sc_hs__clkbuff_8 fanout216 (.Y(net216),
    .A(net219));
 sky130_as_sc_hs__buff_11 fanout217 (.A(net219),
    .Y(net217));
 sky130_as_sc_hs__clkbuff_8 fanout218 (.Y(net218),
    .A(net219));
 sky130_as_sc_hs__buff_11 fanout219 (.A(net230),
    .Y(net219));
 sky130_as_sc_hs__buff_11 fanout220 (.A(net221),
    .Y(net220));
 sky130_as_sc_hs__buff_11 fanout221 (.A(net224),
    .Y(net221));
 sky130_as_sc_hs__buff_11 fanout222 (.A(net223),
    .Y(net222));
 sky130_as_sc_hs__buff_11 fanout223 (.A(net224),
    .Y(net223));
 sky130_as_sc_hs__clkbuff_11 fanout224 (.A(net230),
    .Y(net224));
 sky130_as_sc_hs__buff_11 fanout225 (.A(net227),
    .Y(net225));
 sky130_as_sc_hs__clkbuff_8 fanout226 (.Y(net226),
    .A(net227));
 sky130_as_sc_hs__buff_11 fanout227 (.A(net230),
    .Y(net227));
 sky130_as_sc_hs__buff_11 fanout228 (.A(net229),
    .Y(net228));
 sky130_as_sc_hs__buff_11 fanout229 (.A(net230),
    .Y(net229));
 sky130_as_sc_hs__buff_11 fanout230 (.A(_19484_),
    .Y(net230));
 sky130_as_sc_hs__buff_11 fanout231 (.A(net232),
    .Y(net231));
 sky130_as_sc_hs__buff_11 fanout232 (.A(_19483_),
    .Y(net232));
 sky130_as_sc_hs__buff_11 fanout233 (.A(_19483_),
    .Y(net233));
 sky130_as_sc_hs__clkbuff_11 fanout234 (.A(_19483_),
    .Y(net234));
 sky130_as_sc_hs__buff_11 fanout235 (.A(net239),
    .Y(net235));
 sky130_as_sc_hs__buff_11 fanout236 (.A(net239),
    .Y(net236));
 sky130_as_sc_hs__buff_11 fanout237 (.A(net238),
    .Y(net237));
 sky130_as_sc_hs__buff_11 fanout238 (.A(net239),
    .Y(net238));
 sky130_as_sc_hs__clkbuff_11 fanout239 (.A(_19483_),
    .Y(net239));
 sky130_as_sc_hs__buff_11 fanout240 (.A(net244),
    .Y(net240));
 sky130_as_sc_hs__buff_11 fanout241 (.A(net244),
    .Y(net241));
 sky130_as_sc_hs__buff_11 fanout242 (.A(net244),
    .Y(net242));
 sky130_as_sc_hs__buff_11 fanout243 (.A(net244),
    .Y(net243));
 sky130_as_sc_hs__buff_11 fanout244 (.A(_19482_),
    .Y(net244));
 sky130_as_sc_hs__buff_11 fanout245 (.A(net246),
    .Y(net245));
 sky130_as_sc_hs__buff_11 fanout246 (.A(_19481_),
    .Y(net246));
 sky130_as_sc_hs__buff_11 fanout247 (.A(net248),
    .Y(net247));
 sky130_as_sc_hs__clkbuff_11 fanout248 (.A(_00004_),
    .Y(net248));
 sky130_as_sc_hs__buff_11 fanout249 (.A(net250),
    .Y(net249));
 sky130_as_sc_hs__buff_11 fanout250 (.A(_00003_),
    .Y(net250));
 sky130_as_sc_hs__buff_11 fanout251 (.A(net253),
    .Y(net251));
 sky130_as_sc_hs__buff_11 fanout252 (.A(net253),
    .Y(net252));
 sky130_as_sc_hs__buff_11 fanout253 (.A(_00003_),
    .Y(net253));
 sky130_as_sc_hs__buff_11 fanout254 (.A(net255),
    .Y(net254));
 sky130_as_sc_hs__buff_11 fanout255 (.A(net256),
    .Y(net255));
 sky130_as_sc_hs__buff_11 fanout256 (.A(_00002_),
    .Y(net256));
 sky130_as_sc_hs__buff_11 fanout257 (.A(net259),
    .Y(net257));
 sky130_as_sc_hs__buff_11 fanout258 (.A(net259),
    .Y(net258));
 sky130_as_sc_hs__clkbuff_11 fanout259 (.A(_00002_),
    .Y(net259));
 sky130_as_sc_hs__buff_11 fanout260 (.A(net262),
    .Y(net260));
 sky130_as_sc_hs__buff_11 fanout261 (.A(net262),
    .Y(net261));
 sky130_as_sc_hs__buff_11 fanout262 (.A(_00002_),
    .Y(net262));
 sky130_as_sc_hs__buff_11 fanout263 (.A(net282),
    .Y(net263));
 sky130_as_sc_hs__buff_11 fanout264 (.A(net282),
    .Y(net264));
 sky130_as_sc_hs__buff_11 fanout265 (.A(net282),
    .Y(net265));
 sky130_as_sc_hs__clkbuff_11 fanout266 (.A(net282),
    .Y(net266));
 sky130_as_sc_hs__buff_11 fanout267 (.A(net269),
    .Y(net267));
 sky130_as_sc_hs__buff_11 fanout268 (.A(net269),
    .Y(net268));
 sky130_as_sc_hs__buff_11 fanout269 (.A(net282),
    .Y(net269));
 sky130_as_sc_hs__buff_11 fanout270 (.A(net275),
    .Y(net270));
 sky130_as_sc_hs__buff_11 fanout271 (.A(net275),
    .Y(net271));
 sky130_as_sc_hs__buff_11 fanout272 (.A(net275),
    .Y(net272));
 sky130_as_sc_hs__buff_11 fanout273 (.A(net274),
    .Y(net273));
 sky130_as_sc_hs__clkbuff_11 fanout274 (.A(net275),
    .Y(net274));
 sky130_as_sc_hs__buff_11 fanout275 (.A(net282),
    .Y(net275));
 sky130_as_sc_hs__buff_11 fanout276 (.A(net277),
    .Y(net276));
 sky130_as_sc_hs__buff_11 fanout277 (.A(net281),
    .Y(net277));
 sky130_as_sc_hs__buff_11 fanout278 (.A(net281),
    .Y(net278));
 sky130_as_sc_hs__clkbuff_8 fanout279 (.Y(net279),
    .A(net281));
 sky130_as_sc_hs__buff_11 fanout280 (.A(net281),
    .Y(net280));
 sky130_as_sc_hs__buff_11 fanout281 (.A(net282),
    .Y(net281));
 sky130_as_sc_hs__buff_11 fanout282 (.A(_00001_),
    .Y(net282));
 sky130_as_sc_hs__clkbuff_11 fanout283 (.A(net291),
    .Y(net283));
 sky130_as_sc_hs__buff_4 fanout284 (.A(net291),
    .Y(net284));
 sky130_as_sc_hs__clkbuff_8 fanout285 (.Y(net285),
    .A(net286));
 sky130_as_sc_hs__clkbuff_8 fanout286 (.Y(net286),
    .A(net291));
 sky130_as_sc_hs__clkbuff_11 fanout287 (.A(net291),
    .Y(net287));
 sky130_as_sc_hs__buff_4 fanout288 (.A(net291),
    .Y(net288));
 sky130_as_sc_hs__clkbuff_8 fanout289 (.Y(net289),
    .A(net291));
 sky130_as_sc_hs__buff_4 fanout290 (.A(net291),
    .Y(net290));
 sky130_as_sc_hs__clkbuff_8 fanout291 (.Y(net291),
    .A(net292));
 sky130_as_sc_hs__clkbuff_8 fanout292 (.Y(net292),
    .A(_00000_));
 sky130_as_sc_hs__clkbuff_11 fanout293 (.A(net307),
    .Y(net293));
 sky130_as_sc_hs__buff_4 fanout294 (.A(net295),
    .Y(net294));
 sky130_as_sc_hs__clkbuff_8 fanout295 (.Y(net295),
    .A(net307));
 sky130_as_sc_hs__clkbuff_8 fanout296 (.Y(net296),
    .A(net307));
 sky130_as_sc_hs__clkbuff_8 fanout297 (.Y(net297),
    .A(net298));
 sky130_as_sc_hs__clkbuff_8 fanout298 (.Y(net298),
    .A(net307));
 sky130_as_sc_hs__clkbuff_11 fanout299 (.A(net307),
    .Y(net299));
 sky130_as_sc_hs__buff_4 fanout300 (.A(net307),
    .Y(net300));
 sky130_as_sc_hs__clkbuff_8 fanout301 (.Y(net301),
    .A(net307));
 sky130_as_sc_hs__clkbuff_4 fanout302 (.A(net307),
    .Y(net302));
 sky130_as_sc_hs__clkbuff_8 fanout303 (.Y(net303),
    .A(net306));
 sky130_as_sc_hs__clkbuff_4 fanout304 (.A(net306),
    .Y(net304));
 sky130_as_sc_hs__clkbuff_8 fanout305 (.Y(net305),
    .A(net306));
 sky130_as_sc_hs__buff_4 fanout306 (.A(net307),
    .Y(net306));
 sky130_as_sc_hs__clkbuff_11 fanout307 (.A(_00000_),
    .Y(net307));
 sky130_as_sc_hs__clkbuff_8 fanout308 (.Y(net308),
    .A(net311));
 sky130_as_sc_hs__clkbuff_8 fanout309 (.Y(net309),
    .A(net310));
 sky130_as_sc_hs__buff_4 fanout310 (.A(net311),
    .Y(net310));
 sky130_as_sc_hs__clkbuff_4 fanout311 (.A(net333),
    .Y(net311));
 sky130_as_sc_hs__clkbuff_8 fanout312 (.Y(net312),
    .A(net313));
 sky130_as_sc_hs__clkbuff_8 fanout313 (.Y(net313),
    .A(net333));
 sky130_as_sc_hs__clkbuff_8 fanout314 (.Y(net314),
    .A(net320));
 sky130_as_sc_hs__clkbuff_8 fanout315 (.Y(net315),
    .A(net320));
 sky130_as_sc_hs__clkbuff_8 fanout316 (.Y(net316),
    .A(net320));
 sky130_as_sc_hs__clkbuff_4 fanout317 (.A(net320),
    .Y(net317));
 sky130_as_sc_hs__clkbuff_8 fanout318 (.Y(net318),
    .A(net319));
 sky130_as_sc_hs__clkbuff_8 fanout319 (.Y(net319),
    .A(net320));
 sky130_as_sc_hs__clkbuff_8 fanout320 (.Y(net320),
    .A(net333));
 sky130_as_sc_hs__clkbuff_8 fanout321 (.Y(net321),
    .A(net323));
 sky130_as_sc_hs__clkbuff_4 fanout322 (.A(net323),
    .Y(net322));
 sky130_as_sc_hs__clkbuff_8 fanout323 (.Y(net323),
    .A(net333));
 sky130_as_sc_hs__clkbuff_8 fanout324 (.Y(net324),
    .A(net326));
 sky130_as_sc_hs__clkbuff_8 fanout325 (.Y(net325),
    .A(net326));
 sky130_as_sc_hs__buff_4 fanout326 (.A(net333),
    .Y(net326));
 sky130_as_sc_hs__clkbuff_8 fanout327 (.Y(net327),
    .A(net329));
 sky130_as_sc_hs__clkbuff_8 fanout328 (.Y(net328),
    .A(net329));
 sky130_as_sc_hs__buff_4 fanout329 (.A(net332),
    .Y(net329));
 sky130_as_sc_hs__clkbuff_8 fanout330 (.Y(net330),
    .A(net332));
 sky130_as_sc_hs__clkbuff_8 fanout331 (.Y(net331),
    .A(net332));
 sky130_as_sc_hs__buff_4 fanout332 (.A(net333),
    .Y(net332));
 sky130_as_sc_hs__clkbuff_8 fanout333 (.Y(net333),
    .A(_00000_));
 sky130_as_sc_hs__clkbuff_11 fanout334 (.A(\tholin_riscv.Bimm[12] ),
    .Y(net334));
 sky130_as_sc_hs__buff_11 fanout335 (.A(net336),
    .Y(net335));
 sky130_as_sc_hs__buff_11 fanout336 (.A(\tholin_riscv.Jimm[19] ),
    .Y(net336));
 sky130_as_sc_hs__buff_11 fanout337 (.A(net341),
    .Y(net337));
 sky130_as_sc_hs__buff_11 fanout338 (.A(net341),
    .Y(net338));
 sky130_as_sc_hs__buff_11 fanout339 (.A(net341),
    .Y(net339));
 sky130_as_sc_hs__buff_11 fanout340 (.A(net341),
    .Y(net340));
 sky130_as_sc_hs__buff_11 fanout341 (.A(\tholin_riscv.Jimm[18] ),
    .Y(net341));
 sky130_as_sc_hs__buff_11 fanout342 (.A(net343),
    .Y(net342));
 sky130_as_sc_hs__buff_11 fanout343 (.A(\tholin_riscv.Jimm[17] ),
    .Y(net343));
 sky130_as_sc_hs__buff_11 fanout344 (.A(\tholin_riscv.Jimm[17] ),
    .Y(net344));
 sky130_as_sc_hs__buff_11 fanout345 (.A(\tholin_riscv.Jimm[17] ),
    .Y(net345));
 sky130_as_sc_hs__buff_11 fanout346 (.A(\tholin_riscv.Jimm[17] ),
    .Y(net346));
 sky130_as_sc_hs__buff_11 fanout347 (.A(\tholin_riscv.Jimm[17] ),
    .Y(net347));
 sky130_as_sc_hs__buff_11 fanout348 (.A(net350),
    .Y(net348));
 sky130_as_sc_hs__buff_11 fanout349 (.A(net350),
    .Y(net349));
 sky130_as_sc_hs__buff_11 fanout350 (.A(\tholin_riscv.Jimm[17] ),
    .Y(net350));
 sky130_as_sc_hs__buff_11 fanout351 (.A(net359),
    .Y(net351));
 sky130_as_sc_hs__buff_11 fanout352 (.A(net354),
    .Y(net352));
 sky130_as_sc_hs__clkbuff_8 fanout353 (.Y(net353),
    .A(net354));
 sky130_as_sc_hs__buff_11 fanout354 (.A(net359),
    .Y(net354));
 sky130_as_sc_hs__buff_11 fanout355 (.A(net359),
    .Y(net355));
 sky130_as_sc_hs__clkbuff_11 fanout356 (.A(net359),
    .Y(net356));
 sky130_as_sc_hs__buff_11 fanout357 (.A(net358),
    .Y(net357));
 sky130_as_sc_hs__buff_11 fanout358 (.A(net359),
    .Y(net358));
 sky130_as_sc_hs__buff_11 fanout359 (.A(\tholin_riscv.Jimm[16] ),
    .Y(net359));
 sky130_as_sc_hs__buff_11 fanout360 (.A(net370),
    .Y(net360));
 sky130_as_sc_hs__buff_11 fanout361 (.A(net370),
    .Y(net361));
 sky130_as_sc_hs__buff_11 fanout362 (.A(net363),
    .Y(net362));
 sky130_as_sc_hs__buff_11 fanout363 (.A(net370),
    .Y(net363));
 sky130_as_sc_hs__buff_11 fanout364 (.A(net365),
    .Y(net364));
 sky130_as_sc_hs__buff_11 fanout365 (.A(net370),
    .Y(net365));
 sky130_as_sc_hs__buff_11 fanout366 (.A(net370),
    .Y(net366));
 sky130_as_sc_hs__buff_11 fanout367 (.A(net369),
    .Y(net367));
 sky130_as_sc_hs__buff_4 fanout368 (.A(net369),
    .Y(net368));
 sky130_as_sc_hs__buff_11 fanout369 (.A(net370),
    .Y(net369));
 sky130_as_sc_hs__buff_11 fanout370 (.A(\tholin_riscv.Jimm[16] ),
    .Y(net370));
 sky130_as_sc_hs__clkbuff_8 fanout371 (.Y(net371),
    .A(\tholin_riscv.io_size[1] ));
 sky130_as_sc_hs__clkbuff_8 fanout372 (.Y(net372),
    .A(net373));
 sky130_as_sc_hs__buff_4 fanout373 (.A(net410),
    .Y(net373));
 sky130_as_sc_hs__clkbuff_8 fanout374 (.Y(net374),
    .A(net377));
 sky130_as_sc_hs__clkbuff_8 fanout375 (.Y(net375),
    .A(net377));
 sky130_as_sc_hs__buff_4 fanout376 (.A(net377),
    .Y(net376));
 sky130_as_sc_hs__buff_4 fanout377 (.A(net382),
    .Y(net377));
 sky130_as_sc_hs__clkbuff_8 fanout378 (.Y(net378),
    .A(net382));
 sky130_as_sc_hs__clkbuff_4 fanout379 (.A(net382),
    .Y(net379));
 sky130_as_sc_hs__clkbuff_8 fanout380 (.Y(net380),
    .A(net381));
 sky130_as_sc_hs__clkbuff_8 fanout381 (.Y(net381),
    .A(net382));
 sky130_as_sc_hs__buff_11 fanout382 (.A(net410),
    .Y(net382));
 sky130_as_sc_hs__clkbuff_8 fanout383 (.Y(net383),
    .A(net384));
 sky130_as_sc_hs__clkbuff_8 fanout384 (.Y(net384),
    .A(net410));
 sky130_as_sc_hs__clkbuff_8 fanout385 (.Y(net385),
    .A(net410));
 sky130_as_sc_hs__clkbuff_8 fanout386 (.Y(net386),
    .A(net410));
 sky130_as_sc_hs__clkbuff_8 fanout387 (.Y(net387),
    .A(net388));
 sky130_as_sc_hs__clkbuff_8 fanout388 (.Y(net388),
    .A(net394));
 sky130_as_sc_hs__clkbuff_8 fanout389 (.Y(net389),
    .A(net394));
 sky130_as_sc_hs__clkbuff_8 fanout390 (.Y(net390),
    .A(net394));
 sky130_as_sc_hs__buff_4 fanout391 (.A(net394),
    .Y(net391));
 sky130_as_sc_hs__clkbuff_8 fanout392 (.Y(net392),
    .A(net393));
 sky130_as_sc_hs__clkbuff_8 fanout393 (.Y(net393),
    .A(net394));
 sky130_as_sc_hs__clkbuff_8 fanout394 (.Y(net394),
    .A(net410));
 sky130_as_sc_hs__clkbuff_8 fanout395 (.Y(net395),
    .A(net396));
 sky130_as_sc_hs__clkbuff_8 fanout396 (.Y(net396),
    .A(net409));
 sky130_as_sc_hs__clkbuff_8 fanout397 (.Y(net397),
    .A(net400));
 sky130_as_sc_hs__clkbuff_8 fanout398 (.Y(net398),
    .A(net400));
 sky130_as_sc_hs__clkbuff_4 fanout399 (.A(net400),
    .Y(net399));
 sky130_as_sc_hs__buff_4 fanout400 (.A(net409),
    .Y(net400));
 sky130_as_sc_hs__clkbuff_8 fanout401 (.Y(net401),
    .A(net408));
 sky130_as_sc_hs__buff_4 fanout402 (.A(net408),
    .Y(net402));
 sky130_as_sc_hs__clkbuff_8 fanout403 (.Y(net403),
    .A(net404));
 sky130_as_sc_hs__clkbuff_8 fanout404 (.Y(net404),
    .A(net408));
 sky130_as_sc_hs__clkbuff_8 fanout405 (.Y(net405),
    .A(net408));
 sky130_as_sc_hs__clkbuff_4 fanout406 (.A(net408),
    .Y(net406));
 sky130_as_sc_hs__clkbuff_8 fanout407 (.Y(net407),
    .A(net408));
 sky130_as_sc_hs__clkbuff_8 fanout408 (.Y(net408),
    .A(net409));
 sky130_as_sc_hs__buff_4 fanout409 (.A(net410),
    .Y(net409));
 sky130_as_sc_hs__buff_11 fanout410 (.A(\tholin_riscv.Jimm[15] ),
    .Y(net410));
 sky130_as_sc_hs__clkbuff_11 fanout411 (.A(net1798),
    .Y(net411));
 sky130_as_sc_hs__buff_11 fanout412 (.A(net413),
    .Y(net412));
 sky130_as_sc_hs__buff_11 fanout413 (.A(_21568_),
    .Y(net413));
 sky130_as_sc_hs__clkbuff_8 fanout414 (.Y(net414),
    .A(net415));
 sky130_as_sc_hs__clkbuff_8 fanout415 (.Y(net415),
    .A(_06551_));
 sky130_as_sc_hs__buff_11 fanout416 (.A(net417),
    .Y(net416));
 sky130_as_sc_hs__clkbuff_8 fanout417 (.Y(net417),
    .A(_05513_));
 sky130_as_sc_hs__clkbuff_8 fanout418 (.Y(net418),
    .A(_02550_));
 sky130_as_sc_hs__clkbuff_11 fanout419 (.A(net420),
    .Y(net419));
 sky130_as_sc_hs__buff_11 fanout420 (.A(_02481_),
    .Y(net420));
 sky130_as_sc_hs__clkbuff_8 fanout421 (.Y(net421),
    .A(net422));
 sky130_as_sc_hs__clkbuff_8 fanout422 (.Y(net422),
    .A(_01730_));
 sky130_as_sc_hs__clkbuff_8 fanout423 (.Y(net423),
    .A(net424));
 sky130_as_sc_hs__buff_11 fanout424 (.A(_25874_),
    .Y(net424));
 sky130_as_sc_hs__clkbuff_8 fanout425 (.Y(net425),
    .A(net426));
 sky130_as_sc_hs__clkbuff_11 fanout426 (.A(_25494_),
    .Y(net426));
 sky130_as_sc_hs__clkbuff_11 fanout427 (.A(net428),
    .Y(net427));
 sky130_as_sc_hs__buff_11 fanout428 (.A(_25281_),
    .Y(net428));
 sky130_as_sc_hs__clkbuff_11 fanout429 (.A(net430),
    .Y(net429));
 sky130_as_sc_hs__buff_11 fanout430 (.A(_25255_),
    .Y(net430));
 sky130_as_sc_hs__clkbuff_11 fanout431 (.A(net432),
    .Y(net431));
 sky130_as_sc_hs__buff_11 fanout432 (.A(_25140_),
    .Y(net432));
 sky130_as_sc_hs__clkbuff_8 fanout433 (.Y(net433),
    .A(_25035_));
 sky130_as_sc_hs__clkbuff_8 fanout434 (.Y(net434),
    .A(_24904_));
 sky130_as_sc_hs__clkbuff_8 fanout435 (.Y(net435),
    .A(_24904_));
 sky130_as_sc_hs__clkbuff_8 fanout436 (.Y(net436),
    .A(net437));
 sky130_as_sc_hs__clkbuff_8 fanout437 (.Y(net437),
    .A(_24820_));
 sky130_as_sc_hs__clkbuff_11 fanout438 (.A(net439),
    .Y(net438));
 sky130_as_sc_hs__buff_11 fanout439 (.A(_24795_),
    .Y(net439));
 sky130_as_sc_hs__clkbuff_8 fanout440 (.Y(net440),
    .A(_24780_));
 sky130_as_sc_hs__clkbuff_8 fanout441 (.Y(net441),
    .A(_24780_));
 sky130_as_sc_hs__clkbuff_8 fanout442 (.Y(net442),
    .A(net443));
 sky130_as_sc_hs__clkbuff_8 fanout443 (.Y(net443),
    .A(_24742_));
 sky130_as_sc_hs__clkbuff_8 fanout444 (.Y(net444),
    .A(_24723_));
 sky130_as_sc_hs__clkbuff_8 fanout445 (.Y(net445),
    .A(_24723_));
 sky130_as_sc_hs__clkbuff_11 fanout446 (.A(net447),
    .Y(net446));
 sky130_as_sc_hs__buff_11 fanout447 (.A(_24622_),
    .Y(net447));
 sky130_as_sc_hs__clkbuff_8 fanout448 (.Y(net448),
    .A(net449));
 sky130_as_sc_hs__clkbuff_11 fanout449 (.A(_24596_),
    .Y(net449));
 sky130_as_sc_hs__clkbuff_8 fanout450 (.Y(net450),
    .A(net451));
 sky130_as_sc_hs__clkbuff_11 fanout451 (.A(_24585_),
    .Y(net451));
 sky130_as_sc_hs__clkbuff_11 fanout452 (.A(_24580_),
    .Y(net452));
 sky130_as_sc_hs__clkbuff_8 fanout453 (.Y(net453),
    .A(_24580_));
 sky130_as_sc_hs__clkbuff_8 fanout454 (.Y(net454),
    .A(_24561_));
 sky130_as_sc_hs__clkbuff_8 fanout455 (.Y(net455),
    .A(_24561_));
 sky130_as_sc_hs__clkbuff_8 fanout456 (.Y(net456),
    .A(net457));
 sky130_as_sc_hs__clkbuff_8 fanout457 (.Y(net457),
    .A(_24479_));
 sky130_as_sc_hs__clkbuff_11 fanout458 (.A(_24244_),
    .Y(net458));
 sky130_as_sc_hs__clkbuff_8 fanout459 (.Y(net459),
    .A(_24244_));
 sky130_as_sc_hs__clkbuff_8 fanout460 (.Y(net460),
    .A(_24234_));
 sky130_as_sc_hs__clkbuff_8 fanout461 (.Y(net461),
    .A(_24234_));
 sky130_as_sc_hs__clkbuff_8 fanout462 (.Y(net462),
    .A(net463));
 sky130_as_sc_hs__clkbuff_11 fanout463 (.A(_24221_),
    .Y(net463));
 sky130_as_sc_hs__clkbuff_8 fanout464 (.Y(net464),
    .A(net465));
 sky130_as_sc_hs__clkbuff_11 fanout465 (.A(_24210_),
    .Y(net465));
 sky130_as_sc_hs__clkbuff_8 fanout466 (.Y(net466),
    .A(_24198_));
 sky130_as_sc_hs__buff_4 fanout467 (.A(_24198_),
    .Y(net467));
 sky130_as_sc_hs__clkbuff_8 fanout468 (.Y(net468),
    .A(_24123_));
 sky130_as_sc_hs__buff_4 fanout469 (.A(_24123_),
    .Y(net469));
 sky130_as_sc_hs__clkbuff_8 fanout470 (.Y(net470),
    .A(net471));
 sky130_as_sc_hs__clkbuff_11 fanout471 (.A(_24047_),
    .Y(net471));
 sky130_as_sc_hs__clkbuff_8 fanout472 (.Y(net472),
    .A(net473));
 sky130_as_sc_hs__clkbuff_11 fanout473 (.A(_23680_),
    .Y(net473));
 sky130_as_sc_hs__clkbuff_8 fanout474 (.Y(net474),
    .A(net475));
 sky130_as_sc_hs__buff_11 fanout475 (.A(_23657_),
    .Y(net475));
 sky130_as_sc_hs__clkbuff_11 fanout476 (.A(_23650_),
    .Y(net476));
 sky130_as_sc_hs__clkbuff_11 fanout477 (.A(_23650_),
    .Y(net477));
 sky130_as_sc_hs__clkbuff_11 fanout478 (.A(net479),
    .Y(net478));
 sky130_as_sc_hs__buff_11 fanout479 (.A(_23643_),
    .Y(net479));
 sky130_as_sc_hs__clkbuff_8 fanout480 (.Y(net480),
    .A(net481));
 sky130_as_sc_hs__clkbuff_11 fanout481 (.A(_23629_),
    .Y(net481));
 sky130_as_sc_hs__clkbuff_8 fanout482 (.Y(net482),
    .A(_23624_));
 sky130_as_sc_hs__buff_4 fanout483 (.A(_23624_),
    .Y(net483));
 sky130_as_sc_hs__clkbuff_8 fanout484 (.Y(net484),
    .A(net485));
 sky130_as_sc_hs__buff_4 fanout485 (.A(net487),
    .Y(net485));
 sky130_as_sc_hs__clkbuff_8 fanout486 (.Y(net486),
    .A(net487));
 sky130_as_sc_hs__clkbuff_8 fanout487 (.Y(net487),
    .A(net496));
 sky130_as_sc_hs__clkbuff_8 fanout488 (.Y(net488),
    .A(net489));
 sky130_as_sc_hs__buff_4 fanout489 (.A(net496),
    .Y(net489));
 sky130_as_sc_hs__clkbuff_8 fanout490 (.Y(net490),
    .A(net492));
 sky130_as_sc_hs__clkbuff_11 fanout491 (.A(net492),
    .Y(net491));
 sky130_as_sc_hs__clkbuff_8 fanout492 (.Y(net492),
    .A(net496));
 sky130_as_sc_hs__clkbuff_8 fanout493 (.Y(net493),
    .A(net494));
 sky130_as_sc_hs__clkbuff_8 fanout494 (.Y(net494),
    .A(net495));
 sky130_as_sc_hs__clkbuff_8 fanout495 (.Y(net495),
    .A(net496));
 sky130_as_sc_hs__clkbuff_8 fanout496 (.Y(net496),
    .A(net524));
 sky130_as_sc_hs__clkbuff_8 fanout497 (.Y(net497),
    .A(net499));
 sky130_as_sc_hs__clkbuff_8 fanout498 (.Y(net498),
    .A(net499));
 sky130_as_sc_hs__clkbuff_8 fanout499 (.Y(net499),
    .A(net524));
 sky130_as_sc_hs__clkbuff_8 fanout500 (.Y(net500),
    .A(net502));
 sky130_as_sc_hs__buff_4 fanout501 (.A(net502),
    .Y(net501));
 sky130_as_sc_hs__clkbuff_8 fanout502 (.Y(net502),
    .A(net524));
 sky130_as_sc_hs__clkbuff_8 fanout503 (.Y(net503),
    .A(net504));
 sky130_as_sc_hs__clkbuff_8 fanout504 (.Y(net504),
    .A(net524));
 sky130_as_sc_hs__clkbuff_11 fanout505 (.A(net509),
    .Y(net505));
 sky130_as_sc_hs__clkbuff_8 fanout506 (.Y(net506),
    .A(net509));
 sky130_as_sc_hs__clkbuff_8 fanout507 (.Y(net507),
    .A(net509));
 sky130_as_sc_hs__clkbuff_8 fanout508 (.Y(net508),
    .A(net509));
 sky130_as_sc_hs__clkbuff_8 fanout509 (.Y(net509),
    .A(net514));
 sky130_as_sc_hs__clkbuff_8 fanout510 (.Y(net510),
    .A(net511));
 sky130_as_sc_hs__clkbuff_8 fanout511 (.Y(net511),
    .A(net514));
 sky130_as_sc_hs__clkbuff_8 fanout512 (.Y(net512),
    .A(net514));
 sky130_as_sc_hs__buff_4 fanout513 (.A(net514),
    .Y(net513));
 sky130_as_sc_hs__buff_11 fanout514 (.A(net524),
    .Y(net514));
 sky130_as_sc_hs__clkbuff_8 fanout515 (.Y(net515),
    .A(net517));
 sky130_as_sc_hs__clkbuff_8 fanout516 (.Y(net516),
    .A(net517));
 sky130_as_sc_hs__clkbuff_8 fanout517 (.Y(net517),
    .A(net522));
 sky130_as_sc_hs__clkbuff_8 fanout518 (.Y(net518),
    .A(net522));
 sky130_as_sc_hs__clkbuff_8 fanout519 (.Y(net519),
    .A(net520));
 sky130_as_sc_hs__clkbuff_8 fanout520 (.Y(net520),
    .A(net522));
 sky130_as_sc_hs__clkbuff_8 fanout521 (.Y(net521),
    .A(net522));
 sky130_as_sc_hs__clkbuff_8 fanout522 (.Y(net522),
    .A(net523));
 sky130_as_sc_hs__clkbuff_8 fanout523 (.Y(net523),
    .A(net524));
 sky130_as_sc_hs__buff_11 fanout524 (.A(net22),
    .Y(net524));
 sky130_as_sc_hs__clkbuff_8 fanout525 (.Y(net525),
    .A(net526));
 sky130_as_sc_hs__clkbuff_8 fanout526 (.Y(net526),
    .A(net22));
 sky130_as_sc_hs__buff_11 fanout527 (.A(net22),
    .Y(net527));
 sky130_as_sc_hs__clkbuff_8 fanout74 (.Y(net74),
    .A(net75));
 sky130_as_sc_hs__clkbuff_11 fanout75 (.A(_02725_),
    .Y(net75));
 sky130_as_sc_hs__buff_11 fanout76 (.A(net77),
    .Y(net76));
 sky130_as_sc_hs__buff_11 fanout77 (.A(_13479_),
    .Y(net77));
 sky130_as_sc_hs__clkbuff_11 fanout78 (.A(net79),
    .Y(net78));
 sky130_as_sc_hs__buff_11 fanout79 (.A(_24698_),
    .Y(net79));
 sky130_as_sc_hs__buff_11 fanout80 (.A(_18135_),
    .Y(net80));
 sky130_as_sc_hs__buff_11 fanout81 (.A(_17404_),
    .Y(net81));
 sky130_as_sc_hs__clkbuff_8 fanout82 (.Y(net82),
    .A(_05945_));
 sky130_as_sc_hs__clkbuff_11 fanout83 (.A(_24939_),
    .Y(net83));
 sky130_as_sc_hs__clkbuff_11 fanout84 (.A(_24939_),
    .Y(net84));
 sky130_as_sc_hs__clkbuff_11 fanout85 (.A(_24591_),
    .Y(net85));
 sky130_as_sc_hs__clkbuff_8 fanout86 (.Y(net86),
    .A(_24591_));
 sky130_as_sc_hs__clkbuff_8 fanout87 (.Y(net87),
    .A(net88));
 sky130_as_sc_hs__clkbuff_8 fanout88 (.Y(net88),
    .A(_24550_));
 sky130_as_sc_hs__clkbuff_8 fanout89 (.Y(net89),
    .A(_24537_));
 sky130_as_sc_hs__clkbuff_11 fanout90 (.A(_24128_),
    .Y(net90));
 sky130_as_sc_hs__clkbuff_8 fanout91 (.Y(net91),
    .A(_24128_));
 sky130_as_sc_hs__clkbuff_8 fanout92 (.Y(net92),
    .A(net93));
 sky130_as_sc_hs__clkbuff_8 fanout93 (.Y(net93),
    .A(_18129_));
 sky130_as_sc_hs__clkbuff_8 fanout94 (.Y(net94),
    .A(_17897_));
 sky130_as_sc_hs__clkbuff_8 fanout95 (.Y(net95),
    .A(_17897_));
 sky130_as_sc_hs__clkbuff_8 fanout96 (.Y(net96),
    .A(net97));
 sky130_as_sc_hs__clkbuff_4 fanout97 (.A(net98),
    .Y(net97));
 sky130_as_sc_hs__buff_4 fanout98 (.A(_17398_),
    .Y(net98));
 sky130_as_sc_hs__clkbuff_8 fanout99 (.Y(net99),
    .A(net100));
 sky130_as_sc_hs__buff_2 hold1 (.A(\tholin_riscv.tmr1_pre_ctr[0] ),
    .Y(net542));
 sky130_as_sc_hs__buff_2 hold10 (.A(net1609),
    .Y(net551));
 sky130_as_sc_hs__buff_2 hold100 (.A(_01191_),
    .Y(net641));
 sky130_as_sc_hs__buff_2 hold1000 (.A(_17021_),
    .Y(net1541));
 sky130_as_sc_hs__buff_2 hold1001 (.A(\tholin_riscv.tmr1_pre[20] ),
    .Y(net1542));
 sky130_as_sc_hs__buff_2 hold1002 (.A(_17861_),
    .Y(net1543));
 sky130_as_sc_hs__buff_2 hold1003 (.A(_17863_),
    .Y(net1544));
 sky130_as_sc_hs__buff_2 hold1004 (.A(\tholin_riscv.tmr0_pre[5] ),
    .Y(net1545));
 sky130_as_sc_hs__buff_2 hold1005 (.A(_17914_),
    .Y(net1546));
 sky130_as_sc_hs__buff_2 hold1006 (.A(_17916_),
    .Y(net1547));
 sky130_as_sc_hs__buff_2 hold1007 (.A(\tholin_riscv.intr_vec[17] ),
    .Y(net1548));
 sky130_as_sc_hs__buff_2 hold1008 (.A(_17028_),
    .Y(net1549));
 sky130_as_sc_hs__buff_2 hold1009 (.A(_17030_),
    .Y(net1550));
 sky130_as_sc_hs__buff_2 hold101 (.A(net1789),
    .Y(net642));
 sky130_as_sc_hs__buff_2 hold1010 (.A(\tholin_riscv.tmr0_pre[29] ),
    .Y(net1551));
 sky130_as_sc_hs__buff_2 hold1011 (.A(_17985_),
    .Y(net1552));
 sky130_as_sc_hs__buff_2 hold1012 (.A(_17987_),
    .Y(net1553));
 sky130_as_sc_hs__buff_2 hold1013 (.A(_01501_),
    .Y(net1554));
 sky130_as_sc_hs__buff_2 hold1014 (.A(\tholin_riscv.tmr1_pre[29] ),
    .Y(net1555));
 sky130_as_sc_hs__buff_2 hold1015 (.A(_17888_),
    .Y(net1556));
 sky130_as_sc_hs__buff_2 hold1016 (.A(_17890_),
    .Y(net1557));
 sky130_as_sc_hs__buff_2 hold1017 (.A(_01469_),
    .Y(net1558));
 sky130_as_sc_hs__buff_2 hold1018 (.A(\tholin_riscv.tmr1_pre[28] ),
    .Y(net1559));
 sky130_as_sc_hs__buff_2 hold1019 (.A(_17885_),
    .Y(net1560));
 sky130_as_sc_hs__buff_2 hold102 (.A(_15282_),
    .Y(net643));
 sky130_as_sc_hs__buff_2 hold1020 (.A(_17887_),
    .Y(net1561));
 sky130_as_sc_hs__buff_2 hold1021 (.A(\tholin_riscv.requested_addr[26] ),
    .Y(net1562));
 sky130_as_sc_hs__buff_2 hold1022 (.A(_16945_),
    .Y(net1563));
 sky130_as_sc_hs__buff_2 hold1023 (.A(_16946_),
    .Y(net1564));
 sky130_as_sc_hs__buff_2 hold1024 (.A(\tholin_riscv.requested_addr[10] ),
    .Y(net1565));
 sky130_as_sc_hs__buff_2 hold1025 (.A(_16849_),
    .Y(net1566));
 sky130_as_sc_hs__buff_2 hold1026 (.A(_16850_),
    .Y(net1567));
 sky130_as_sc_hs__buff_2 hold1027 (.A(\tholin_riscv.tmr0_pre[22] ),
    .Y(net1568));
 sky130_as_sc_hs__buff_2 hold1028 (.A(_17964_),
    .Y(net1569));
 sky130_as_sc_hs__buff_2 hold1029 (.A(_17966_),
    .Y(net1570));
 sky130_as_sc_hs__buff_2 hold103 (.A(_01087_),
    .Y(net644));
 sky130_as_sc_hs__buff_2 hold1030 (.A(\tholin_riscv.requested_addr[30] ),
    .Y(net1571));
 sky130_as_sc_hs__buff_2 hold1031 (.A(_16969_),
    .Y(net1572));
 sky130_as_sc_hs__buff_2 hold1032 (.A(_16970_),
    .Y(net1573));
 sky130_as_sc_hs__buff_2 hold1033 (.A(\tholin_riscv.requested_addr[19] ),
    .Y(net1574));
 sky130_as_sc_hs__buff_2 hold1034 (.A(_16903_),
    .Y(net1575));
 sky130_as_sc_hs__buff_2 hold1035 (.A(_16904_),
    .Y(net1576));
 sky130_as_sc_hs__buff_2 hold1036 (.A(\tholin_riscv.tmr1_pre[9] ),
    .Y(net1577));
 sky130_as_sc_hs__buff_2 hold1037 (.A(_17829_),
    .Y(net1578));
 sky130_as_sc_hs__buff_2 hold1038 (.A(_17831_),
    .Y(net1579));
 sky130_as_sc_hs__buff_2 hold1039 (.A(\tholin_riscv.tmr1_pre[26] ),
    .Y(net1580));
 sky130_as_sc_hs__buff_2 hold104 (.A(net1790),
    .Y(net645));
 sky130_as_sc_hs__buff_2 hold1040 (.A(_17879_),
    .Y(net1581));
 sky130_as_sc_hs__buff_2 hold1041 (.A(_17881_),
    .Y(net1582));
 sky130_as_sc_hs__buff_2 hold1042 (.A(_01466_),
    .Y(net1583));
 sky130_as_sc_hs__buff_2 hold1043 (.A(\tholin_riscv.tmr0_pre[26] ),
    .Y(net1584));
 sky130_as_sc_hs__buff_2 hold1044 (.A(_17976_),
    .Y(net1585));
 sky130_as_sc_hs__buff_2 hold1045 (.A(_17978_),
    .Y(net1586));
 sky130_as_sc_hs__buff_2 hold1046 (.A(_01498_),
    .Y(net1587));
 sky130_as_sc_hs__buff_2 hold1047 (.A(\tholin_riscv.tmr1_pre[10] ),
    .Y(net1588));
 sky130_as_sc_hs__buff_2 hold1048 (.A(_17832_),
    .Y(net1589));
 sky130_as_sc_hs__buff_2 hold1049 (.A(\tholin_riscv.requested_addr[15] ),
    .Y(net1590));
 sky130_as_sc_hs__buff_2 hold105 (.A(_15278_),
    .Y(net646));
 sky130_as_sc_hs__buff_2 hold1050 (.A(_16879_),
    .Y(net1591));
 sky130_as_sc_hs__buff_2 hold1051 (.A(_16880_),
    .Y(net1592));
 sky130_as_sc_hs__buff_2 hold1052 (.A(\tholin_riscv.intr_vec[26] ),
    .Y(net1593));
 sky130_as_sc_hs__buff_2 hold1053 (.A(_17055_),
    .Y(net1594));
 sky130_as_sc_hs__buff_2 hold1054 (.A(\tholin_riscv.requested_addr[1] ),
    .Y(net1595));
 sky130_as_sc_hs__buff_2 hold1055 (.A(_16795_),
    .Y(net1596));
 sky130_as_sc_hs__buff_4 hold1056 (.A(\tholin_riscv.instr[1] ),
    .Y(net1597));
 sky130_as_sc_hs__buff_2 hold1057 (.A(\tholin_riscv.requested_addr[16] ),
    .Y(net1598));
 sky130_as_sc_hs__buff_2 hold1058 (.A(_16885_),
    .Y(net1599));
 sky130_as_sc_hs__buff_2 hold1059 (.A(\tholin_riscv.requested_addr[25] ),
    .Y(net1600));
 sky130_as_sc_hs__buff_2 hold106 (.A(_01085_),
    .Y(net647));
 sky130_as_sc_hs__buff_2 hold1060 (.A(_16939_),
    .Y(net1601));
 sky130_as_sc_hs__buff_2 hold1061 (.A(\tholin_riscv.io_int_enable ),
    .Y(net1602));
 sky130_as_sc_hs__buff_2 hold1062 (.A(\tholin_riscv.requested_addr[21] ),
    .Y(net1603));
 sky130_as_sc_hs__buff_2 hold1063 (.A(_16915_),
    .Y(net1604));
 sky130_as_sc_hs__buff_2 hold1064 (.A(\tholin_riscv.requested_addr[24] ),
    .Y(net1605));
 sky130_as_sc_hs__buff_2 hold1065 (.A(_16933_),
    .Y(net1606));
 sky130_as_sc_hs__buff_2 hold1066 (.A(\tholin_riscv.uart.div_counter[12] ),
    .Y(net1607));
 sky130_as_sc_hs__buff_2 hold1067 (.A(_14761_),
    .Y(net1608));
 sky130_as_sc_hs__buff_2 hold1068 (.A(\tholin_riscv.timer_int_enable ),
    .Y(net1609));
 sky130_as_sc_hs__buff_2 hold1069 (.A(\tholin_riscv.requested_addr[12] ),
    .Y(net1610));
 sky130_as_sc_hs__buff_2 hold107 (.A(net1797),
    .Y(net648));
 sky130_as_sc_hs__buff_2 hold1070 (.A(_16861_),
    .Y(net1611));
 sky130_as_sc_hs__buff_2 hold1071 (.A(\tholin_riscv.requested_addr[9] ),
    .Y(net1612));
 sky130_as_sc_hs__buff_2 hold1072 (.A(_16843_),
    .Y(net1613));
 sky130_as_sc_hs__buff_2 hold1073 (.A(\tholin_riscv.requested_addr[29] ),
    .Y(net1614));
 sky130_as_sc_hs__buff_2 hold1074 (.A(_16963_),
    .Y(net1615));
 sky130_as_sc_hs__buff_2 hold1075 (.A(\tholin_riscv.requested_addr[20] ),
    .Y(net1616));
 sky130_as_sc_hs__buff_2 hold1076 (.A(_16909_),
    .Y(net1617));
 sky130_as_sc_hs__buff_2 hold1077 (.A(\tholin_riscv.requested_addr[13] ),
    .Y(net1618));
 sky130_as_sc_hs__buff_2 hold1078 (.A(_16867_),
    .Y(net1619));
 sky130_as_sc_hs__buff_2 hold1079 (.A(\tholin_riscv.uart.div_counter[11] ),
    .Y(net1620));
 sky130_as_sc_hs__buff_2 hold108 (.A(_15262_),
    .Y(net649));
 sky130_as_sc_hs__buff_2 hold1080 (.A(_14755_),
    .Y(net1621));
 sky130_as_sc_hs__buff_2 hold1081 (.A(\tholin_riscv.requested_addr[28] ),
    .Y(net1622));
 sky130_as_sc_hs__buff_2 hold1082 (.A(_16957_),
    .Y(net1623));
 sky130_as_sc_hs__buff_2 hold1083 (.A(\tholin_riscv.uart.div_counter[10] ),
    .Y(net1624));
 sky130_as_sc_hs__buff_2 hold1084 (.A(_14749_),
    .Y(net1625));
 sky130_as_sc_hs__buff_2 hold1085 (.A(\tholin_riscv.uart.div_counter[9] ),
    .Y(net1626));
 sky130_as_sc_hs__buff_2 hold1086 (.A(_14743_),
    .Y(net1627));
 sky130_as_sc_hs__buff_2 hold1087 (.A(\tholin_riscv.instr[3] ),
    .Y(net1628));
 sky130_as_sc_hs__buff_2 hold1088 (.A(_21148_),
    .Y(net1629));
 sky130_as_sc_hs__buff_2 hold1089 (.A(\tholin_riscv.PC[0] ),
    .Y(net1630));
 sky130_as_sc_hs__buff_2 hold109 (.A(_01081_),
    .Y(net650));
 sky130_as_sc_hs__buff_2 hold1090 (.A(_13556_),
    .Y(net1631));
 sky130_as_sc_hs__buff_2 hold1091 (.A(\tholin_riscv.requested_addr[17] ),
    .Y(net1632));
 sky130_as_sc_hs__buff_2 hold1092 (.A(_16891_),
    .Y(net1633));
 sky130_as_sc_hs__buff_2 hold1093 (.A(\tholin_riscv.instr[4] ),
    .Y(net1634));
 sky130_as_sc_hs__buff_2 hold1094 (.A(_21249_),
    .Y(net1635));
 sky130_as_sc_hs__buff_2 hold1095 (.A(\tholin_riscv.uart.div_counter[13] ),
    .Y(net1636));
 sky130_as_sc_hs__buff_2 hold1096 (.A(_14767_),
    .Y(net1637));
 sky130_as_sc_hs__buff_2 hold1097 (.A(\tholin_riscv.requested_addr[8] ),
    .Y(net1638));
 sky130_as_sc_hs__buff_2 hold1098 (.A(_16837_),
    .Y(net1639));
 sky130_as_sc_hs__buff_2 hold1099 (.A(\tholin_riscv.instr[2] ),
    .Y(net1640));
 sky130_as_sc_hs__buff_2 hold11 (.A(_18582_),
    .Y(net552));
 sky130_as_sc_hs__buff_2 hold110 (.A(net1801),
    .Y(net651));
 sky130_as_sc_hs__buff_2 hold1100 (.A(_21044_),
    .Y(net1641));
 sky130_as_sc_hs__buff_2 hold1101 (.A(\tholin_riscv.PC[1] ),
    .Y(net1642));
 sky130_as_sc_hs__buff_2 hold1102 (.A(_13078_),
    .Y(net1643));
 sky130_as_sc_hs__buff_2 hold1103 (.A(\tholin_riscv.cycle[1] ),
    .Y(net1644));
 sky130_as_sc_hs__buff_2 hold1104 (.A(_16394_),
    .Y(net1645));
 sky130_as_sc_hs__buff_2 hold1105 (.A(_01225_),
    .Y(net1646));
 sky130_as_sc_hs__buff_2 hold1106 (.A(\tholin_riscv.uart.div_counter[0] ),
    .Y(net1647));
 sky130_as_sc_hs__buff_2 hold1107 (.A(_14632_),
    .Y(net1648));
 sky130_as_sc_hs__buff_2 hold1108 (.A(_14691_),
    .Y(net1649));
 sky130_as_sc_hs__buff_2 hold1109 (.A(net61),
    .Y(net1650));
 sky130_as_sc_hs__buff_2 hold111 (.A(_13282_),
    .Y(net652));
 sky130_as_sc_hs__buff_2 hold1110 (.A(_18600_),
    .Y(net1651));
 sky130_as_sc_hs__buff_2 hold1111 (.A(net62),
    .Y(net1652));
 sky130_as_sc_hs__buff_2 hold1112 (.A(_18603_),
    .Y(net1653));
 sky130_as_sc_hs__buff_2 hold1113 (.A(\tholin_riscv.instr[5] ),
    .Y(net1654));
 sky130_as_sc_hs__buff_2 hold1114 (.A(net60),
    .Y(net1655));
 sky130_as_sc_hs__buff_2 hold1115 (.A(_18597_),
    .Y(net1656));
 sky130_as_sc_hs__buff_2 hold1116 (.A(net64),
    .Y(net1657));
 sky130_as_sc_hs__buff_2 hold1117 (.A(_18606_),
    .Y(net1658));
 sky130_as_sc_hs__buff_2 hold1118 (.A(net65),
    .Y(net1659));
 sky130_as_sc_hs__buff_2 hold1119 (.A(_18609_),
    .Y(net1660));
 sky130_as_sc_hs__buff_2 hold112 (.A(_00310_),
    .Y(net653));
 sky130_as_sc_hs__buff_2 hold1120 (.A(\tholin_riscv.PC[5] ),
    .Y(net1661));
 sky130_as_sc_hs__buff_2 hold1121 (.A(_18860_),
    .Y(net1662));
 sky130_as_sc_hs__buff_2 hold1122 (.A(\tholin_riscv.PC[10] ),
    .Y(net1663));
 sky130_as_sc_hs__buff_2 hold1123 (.A(_18961_),
    .Y(net1664));
 sky130_as_sc_hs__buff_2 hold1124 (.A(\tholin_riscv.uart.receive_div_counter[0] ),
    .Y(net1665));
 sky130_as_sc_hs__buff_2 hold1125 (.A(_14970_),
    .Y(net1666));
 sky130_as_sc_hs__buff_2 hold1126 (.A(\tholin_riscv.PC[4] ),
    .Y(net1667));
 sky130_as_sc_hs__buff_2 hold1127 (.A(_18840_),
    .Y(net1668));
 sky130_as_sc_hs__buff_2 hold1128 (.A(\tholin_riscv.PC[8] ),
    .Y(net1669));
 sky130_as_sc_hs__buff_2 hold1129 (.A(_18920_),
    .Y(net1670));
 sky130_as_sc_hs__buff_2 hold113 (.A(net1800),
    .Y(net654));
 sky130_as_sc_hs__buff_2 hold1130 (.A(net66),
    .Y(net1671));
 sky130_as_sc_hs__buff_2 hold1131 (.A(_18612_),
    .Y(net1672));
 sky130_as_sc_hs__buff_2 hold1132 (.A(\tholin_riscv.PC[6] ),
    .Y(net1673));
 sky130_as_sc_hs__buff_2 hold1133 (.A(\tholin_riscv.PC[11] ),
    .Y(net1674));
 sky130_as_sc_hs__buff_2 hold1134 (.A(_18984_),
    .Y(net1675));
 sky130_as_sc_hs__buff_2 hold1135 (.A(\tholin_riscv.PC[9] ),
    .Y(net1676));
 sky130_as_sc_hs__buff_2 hold1136 (.A(_18941_),
    .Y(net1677));
 sky130_as_sc_hs__buff_2 hold1137 (.A(\tholin_riscv.Jimm[12] ),
    .Y(net1678));
 sky130_as_sc_hs__buff_2 hold1138 (.A(\tholin_riscv.PC[13] ),
    .Y(net1679));
 sky130_as_sc_hs__buff_2 hold1139 (.A(\tholin_riscv.PC[3] ),
    .Y(net1680));
 sky130_as_sc_hs__buff_2 hold114 (.A(_12953_),
    .Y(net655));
 sky130_as_sc_hs__buff_2 hold1140 (.A(\tholin_riscv.PC[14] ),
    .Y(net1681));
 sky130_as_sc_hs__buff_2 hold1141 (.A(\tholin_riscv.spi.div_counter[0] ),
    .Y(net1682));
 sky130_as_sc_hs__buff_2 hold1142 (.A(\tholin_riscv.PC[27] ),
    .Y(net1683));
 sky130_as_sc_hs__buff_2 hold1143 (.A(\tholin_riscv.instr[1] ),
    .Y(net1684));
 sky130_as_sc_hs__buff_2 hold1144 (.A(net1597),
    .Y(net1685));
 sky130_as_sc_hs__buff_2 hold1145 (.A(\tholin_riscv.PC[23] ),
    .Y(net1686));
 sky130_as_sc_hs__buff_2 hold1146 (.A(\tholin_riscv.PC[7] ),
    .Y(net1687));
 sky130_as_sc_hs__buff_2 hold1147 (.A(\tholin_riscv.Bimm[11] ),
    .Y(net1688));
 sky130_as_sc_hs__buff_2 hold1148 (.A(\tholin_riscv.PC[24] ),
    .Y(net1689));
 sky130_as_sc_hs__buff_2 hold1149 (.A(\tholin_riscv.Jimm[13] ),
    .Y(net1690));
 sky130_as_sc_hs__buff_2 hold115 (.A(_00181_),
    .Y(net656));
 sky130_as_sc_hs__buff_2 hold1150 (.A(\tholin_riscv.requested_addr[0] ),
    .Y(net1691));
 sky130_as_sc_hs__buff_2 hold1151 (.A(\tholin_riscv.PC[15] ),
    .Y(net1692));
 sky130_as_sc_hs__buff_2 hold1152 (.A(\tholin_riscv.PC[26] ),
    .Y(net1693));
 sky130_as_sc_hs__buff_2 hold1153 (.A(\tholin_riscv.uart.counter[0] ),
    .Y(net1694));
 sky130_as_sc_hs__buff_2 hold1154 (.A(\tholin_riscv.PC[25] ),
    .Y(net1695));
 sky130_as_sc_hs__buff_2 hold1155 (.A(\tholin_riscv.PC[28] ),
    .Y(net1696));
 sky130_as_sc_hs__buff_2 hold1156 (.A(\tholin_riscv.PC[29] ),
    .Y(net1697));
 sky130_as_sc_hs__buff_2 hold1157 (.A(\tholin_riscv.PC[18] ),
    .Y(net1698));
 sky130_as_sc_hs__buff_2 hold1158 (.A(\tholin_riscv.uart.receive_counter[2] ),
    .Y(net1699));
 sky130_as_sc_hs__buff_2 hold1159 (.A(\tholin_riscv.PC[17] ),
    .Y(net1700));
 sky130_as_sc_hs__buff_2 hold116 (.A(net1812),
    .Y(net657));
 sky130_as_sc_hs__buff_2 hold1160 (.A(\tholin_riscv.PC[16] ),
    .Y(net1701));
 sky130_as_sc_hs__buff_2 hold1161 (.A(\tholin_riscv.PC[20] ),
    .Y(net1702));
 sky130_as_sc_hs__buff_2 hold1162 (.A(\tholin_riscv.requested_addr[6] ),
    .Y(net1703));
 sky130_as_sc_hs__buff_2 hold1163 (.A(\tholin_riscv.PC[22] ),
    .Y(net1704));
 sky130_as_sc_hs__buff_2 hold1164 (.A(\tholin_riscv.cycle[0] ),
    .Y(net1705));
 sky130_as_sc_hs__buff_2 hold1165 (.A(\tholin_riscv.PC[12] ),
    .Y(net1706));
 sky130_as_sc_hs__buff_2 hold1166 (.A(\tholin_riscv.PC[21] ),
    .Y(net1707));
 sky130_as_sc_hs__buff_2 hold1167 (.A(\tholin_riscv.PC[19] ),
    .Y(net1708));
 sky130_as_sc_hs__buff_2 hold1168 (.A(\tholin_riscv.uart.counter[1] ),
    .Y(net1709));
 sky130_as_sc_hs__buff_2 hold1169 (.A(\tholin_riscv.Bimm[1] ),
    .Y(net1710));
 sky130_as_sc_hs__buff_2 hold117 (.A(_13958_),
    .Y(net658));
 sky130_as_sc_hs__buff_2 hold1170 (.A(net542),
    .Y(net1711));
 sky130_as_sc_hs__buff_2 hold1171 (.A(_01192_),
    .Y(net1712));
 sky130_as_sc_hs__buff_2 hold1172 (.A(net543),
    .Y(net1713));
 sky130_as_sc_hs__buff_2 hold1173 (.A(net544),
    .Y(net1714));
 sky130_as_sc_hs__buff_2 hold1174 (.A(_01312_),
    .Y(net1715));
 sky130_as_sc_hs__buff_2 hold1175 (.A(net545),
    .Y(net1716));
 sky130_as_sc_hs__buff_2 hold1176 (.A(\tholin_riscv.uart.has_byte ),
    .Y(net1717));
 sky130_as_sc_hs__buff_2 hold1177 (.A(net546),
    .Y(net1718));
 sky130_as_sc_hs__buff_2 hold1178 (.A(_01573_),
    .Y(net1719));
 sky130_as_sc_hs__buff_2 hold1179 (.A(net547),
    .Y(net1720));
 sky130_as_sc_hs__buff_2 hold118 (.A(_00663_),
    .Y(net659));
 sky130_as_sc_hs__buff_2 hold1180 (.A(\tholin_riscv.irqs[1] ),
    .Y(net1721));
 sky130_as_sc_hs__buff_2 hold1181 (.A(_19529_),
    .Y(net1722));
 sky130_as_sc_hs__buff_2 hold1182 (.A(\tholin_riscv.uart.receive_buff[4] ),
    .Y(net1723));
 sky130_as_sc_hs__buff_2 hold1183 (.A(net554),
    .Y(net1724));
 sky130_as_sc_hs__buff_2 hold1184 (.A(_00975_),
    .Y(net1725));
 sky130_as_sc_hs__buff_2 hold1185 (.A(net556),
    .Y(net1726));
 sky130_as_sc_hs__buff_2 hold1186 (.A(\tholin_riscv.spi.data_in_buff[7] ),
    .Y(net1727));
 sky130_as_sc_hs__buff_2 hold1187 (.A(net557),
    .Y(net1728));
 sky130_as_sc_hs__buff_2 hold1188 (.A(_01044_),
    .Y(net1729));
 sky130_as_sc_hs__buff_2 hold1189 (.A(net559),
    .Y(net1730));
 sky130_as_sc_hs__buff_2 hold119 (.A(net1805),
    .Y(net660));
 sky130_as_sc_hs__buff_2 hold1190 (.A(\tholin_riscv.spi.data_in_buff[3] ),
    .Y(net1731));
 sky130_as_sc_hs__buff_2 hold1191 (.A(net560),
    .Y(net1732));
 sky130_as_sc_hs__buff_2 hold1192 (.A(_01040_),
    .Y(net1733));
 sky130_as_sc_hs__buff_2 hold1193 (.A(net562),
    .Y(net1734));
 sky130_as_sc_hs__buff_2 hold1194 (.A(\tholin_riscv.uart.dout[7] ),
    .Y(net1735));
 sky130_as_sc_hs__buff_2 hold1195 (.A(_14804_),
    .Y(net1736));
 sky130_as_sc_hs__buff_2 hold1196 (.A(\tholin_riscv.spi.dout[2] ),
    .Y(net1737));
 sky130_as_sc_hs__buff_2 hold1197 (.A(_15110_),
    .Y(net1738));
 sky130_as_sc_hs__buff_2 hold1198 (.A(_01039_),
    .Y(net1739));
 sky130_as_sc_hs__buff_2 hold1199 (.A(\tholin_riscv.spi.dout[5] ),
    .Y(net1740));
 sky130_as_sc_hs__buff_2 hold12 (.A(_01572_),
    .Y(net553));
 sky130_as_sc_hs__buff_2 hold120 (.A(_13759_),
    .Y(net661));
 sky130_as_sc_hs__buff_2 hold1200 (.A(_15119_),
    .Y(net1741));
 sky130_as_sc_hs__buff_2 hold1201 (.A(_01042_),
    .Y(net1742));
 sky130_as_sc_hs__buff_2 hold1202 (.A(net565),
    .Y(net1743));
 sky130_as_sc_hs__buff_2 hold1203 (.A(\tholin_riscv.uart.dout[5] ),
    .Y(net1744));
 sky130_as_sc_hs__buff_2 hold1204 (.A(_14798_),
    .Y(net1745));
 sky130_as_sc_hs__buff_2 hold1205 (.A(_00976_),
    .Y(net1746));
 sky130_as_sc_hs__buff_2 hold1206 (.A(\tholin_riscv.uart.dout[3] ),
    .Y(net1747));
 sky130_as_sc_hs__buff_2 hold1207 (.A(_14792_),
    .Y(net1748));
 sky130_as_sc_hs__buff_2 hold1208 (.A(_00974_),
    .Y(net1749));
 sky130_as_sc_hs__buff_2 hold1209 (.A(\tholin_riscv.uart.dout[0] ),
    .Y(net1750));
 sky130_as_sc_hs__buff_2 hold121 (.A(_00567_),
    .Y(net662));
 sky130_as_sc_hs__buff_2 hold1210 (.A(_14783_),
    .Y(net1751));
 sky130_as_sc_hs__buff_2 hold1211 (.A(_00971_),
    .Y(net1752));
 sky130_as_sc_hs__buff_2 hold1212 (.A(\tholin_riscv.uart.dout[2] ),
    .Y(net1753));
 sky130_as_sc_hs__buff_2 hold1213 (.A(_14789_),
    .Y(net1754));
 sky130_as_sc_hs__buff_2 hold1214 (.A(_00973_),
    .Y(net1755));
 sky130_as_sc_hs__buff_2 hold1215 (.A(\tholin_riscv.uart.dout[6] ),
    .Y(net1756));
 sky130_as_sc_hs__buff_2 hold1216 (.A(_14801_),
    .Y(net1757));
 sky130_as_sc_hs__buff_2 hold1217 (.A(_00977_),
    .Y(net1758));
 sky130_as_sc_hs__buff_2 hold1218 (.A(\tholin_riscv.uart.dout[1] ),
    .Y(net1759));
 sky130_as_sc_hs__buff_2 hold1219 (.A(_14786_),
    .Y(net1760));
 sky130_as_sc_hs__buff_2 hold122 (.A(net1802),
    .Y(net663));
 sky130_as_sc_hs__buff_2 hold1220 (.A(_00972_),
    .Y(net1761));
 sky130_as_sc_hs__buff_2 hold1221 (.A(\tholin_riscv.spi.dout[4] ),
    .Y(net1762));
 sky130_as_sc_hs__buff_2 hold1222 (.A(_15116_),
    .Y(net1763));
 sky130_as_sc_hs__buff_2 hold1223 (.A(_01041_),
    .Y(net1764));
 sky130_as_sc_hs__buff_2 hold1224 (.A(\tholin_riscv.spi.dout[1] ),
    .Y(net1765));
 sky130_as_sc_hs__buff_2 hold1225 (.A(_15107_),
    .Y(net1766));
 sky130_as_sc_hs__buff_2 hold1226 (.A(_01038_),
    .Y(net1767));
 sky130_as_sc_hs__buff_2 hold1227 (.A(\tholin_riscv.spi.dout[6] ),
    .Y(net1768));
 sky130_as_sc_hs__buff_2 hold1228 (.A(_15122_),
    .Y(net1769));
 sky130_as_sc_hs__buff_2 hold1229 (.A(_01043_),
    .Y(net1770));
 sky130_as_sc_hs__buff_2 hold123 (.A(_14024_),
    .Y(net664));
 sky130_as_sc_hs__buff_2 hold1230 (.A(\tholin_riscv.tmr0_pre[8] ),
    .Y(net1771));
 sky130_as_sc_hs__buff_2 hold1231 (.A(_17923_),
    .Y(net1772));
 sky130_as_sc_hs__buff_2 hold1232 (.A(\tholin_riscv.uart.data_buff[9] ),
    .Y(net1773));
 sky130_as_sc_hs__buff_2 hold1233 (.A(\tholin_riscv.current_irq[0] ),
    .Y(net1774));
 sky130_as_sc_hs__buff_2 hold1234 (.A(\tholin_riscv.spi.busy ),
    .Y(net1775));
 sky130_as_sc_hs__buff_2 hold1235 (.A(\tholin_riscv.spi.divisor[1] ),
    .Y(net1776));
 sky130_as_sc_hs__buff_2 hold1236 (.A(\tholin_riscv.uart.counter[3] ),
    .Y(net1777));
 sky130_as_sc_hs__buff_2 hold1237 (.A(\tholin_riscv.spi.divisor[2] ),
    .Y(net1778));
 sky130_as_sc_hs__buff_2 hold1238 (.A(\tholin_riscv.Bimm[9] ),
    .Y(net1779));
 sky130_as_sc_hs__clkbuff_4 hold1239 (.A(\tholin_riscv.Bimm[2] ),
    .Y(net1780));
 sky130_as_sc_hs__buff_2 hold124 (.A(_00695_),
    .Y(net665));
 sky130_as_sc_hs__buff_2 hold1240 (.A(\tholin_riscv.Bimm[6] ),
    .Y(net1781));
 sky130_as_sc_hs__buff_2 hold1241 (.A(\tholin_riscv.mul_delay ),
    .Y(net1782));
 sky130_as_sc_hs__buff_2 hold1242 (.A(\tholin_riscv.spi.divisor[5] ),
    .Y(net1783));
 sky130_as_sc_hs__buff_2 hold1243 (.A(\tholin_riscv.load_dest[3] ),
    .Y(net1784));
 sky130_as_sc_hs__buff_2 hold1244 (.A(\tholin_riscv.load_funct ),
    .Y(net1785));
 sky130_as_sc_hs__buff_2 hold1245 (.A(\tholin_riscv.spi.divisor[0] ),
    .Y(net1786));
 sky130_as_sc_hs__buff_2 hold1246 (.A(\tholin_riscv.load_dest[4] ),
    .Y(net1787));
 sky130_as_sc_hs__buff_2 hold1247 (.A(\tholin_riscv.load_dest[1] ),
    .Y(net1788));
 sky130_as_sc_hs__buff_2 hold1248 (.A(\tholin_riscv.load_dest[2] ),
    .Y(net1789));
 sky130_as_sc_hs__buff_2 hold1249 (.A(\tholin_riscv.load_dest[0] ),
    .Y(net1790));
 sky130_as_sc_hs__buff_2 hold125 (.A(net1804),
    .Y(net666));
 sky130_as_sc_hs__buff_4 hold1250 (.A(\tholin_riscv.Bimm[3] ),
    .Y(net1791));
 sky130_as_sc_hs__clkbuff_4 hold1251 (.A(\tholin_riscv.Bimm[4] ),
    .Y(net1792));
 sky130_as_sc_hs__buff_2 hold1252 (.A(\tholin_riscv.Bimm[3] ),
    .Y(net1793));
 sky130_as_sc_hs__buff_2 hold1253 (.A(\tholin_riscv.Bimm[4] ),
    .Y(net1794));
 sky130_as_sc_hs__buff_2 hold1254 (.A(\tholin_riscv.irqs[0] ),
    .Y(net1795));
 sky130_as_sc_hs__buff_2 hold1255 (.A(\tholin_riscv.Jimm[14] ),
    .Y(net1796));
 sky130_as_sc_hs__buff_2 hold1256 (.A(\tholin_riscv.spi.divisor[4] ),
    .Y(net1797));
 sky130_as_sc_hs__buff_2 hold1257 (.A(\tholin_riscv.Jimm[14] ),
    .Y(net1798));
 sky130_as_sc_hs__buff_2 hold1258 (.A(\tholin_riscv.tmr1_pre_ctr[30] ),
    .Y(net1799));
 sky130_as_sc_hs__buff_2 hold1259 (.A(\tholin_riscv.regs[20][0] ),
    .Y(net1800));
 sky130_as_sc_hs__buff_2 hold126 (.A(_13150_),
    .Y(net667));
 sky130_as_sc_hs__buff_2 hold1260 (.A(\tholin_riscv.regs[13][0] ),
    .Y(net1801));
 sky130_as_sc_hs__buff_2 hold1261 (.A(\tholin_riscv.regs[24][0] ),
    .Y(net1802));
 sky130_as_sc_hs__buff_2 hold1262 (.A(\tholin_riscv.regs[30][0] ),
    .Y(net1803));
 sky130_as_sc_hs__buff_2 hold1263 (.A(\tholin_riscv.regs[17][0] ),
    .Y(net1804));
 sky130_as_sc_hs__buff_2 hold1264 (.A(\tholin_riscv.regs[28][0] ),
    .Y(net1805));
 sky130_as_sc_hs__buff_2 hold1265 (.A(\tholin_riscv.regs[7][0] ),
    .Y(net1806));
 sky130_as_sc_hs__buff_2 hold1266 (.A(\tholin_riscv.regs[29][0] ),
    .Y(net1807));
 sky130_as_sc_hs__buff_2 hold1267 (.A(\tholin_riscv.regs[3][0] ),
    .Y(net1808));
 sky130_as_sc_hs__buff_2 hold1268 (.A(\tholin_riscv.regs[9][0] ),
    .Y(net1809));
 sky130_as_sc_hs__buff_2 hold1269 (.A(\tholin_riscv.regs[12][0] ),
    .Y(net1810));
 sky130_as_sc_hs__buff_2 hold127 (.A(_00246_),
    .Y(net668));
 sky130_as_sc_hs__buff_2 hold1270 (.A(\tholin_riscv.regs[10][0] ),
    .Y(net1811));
 sky130_as_sc_hs__buff_2 hold1271 (.A(\tholin_riscv.regs[25][0] ),
    .Y(net1812));
 sky130_as_sc_hs__buff_2 hold1272 (.A(\tholin_riscv.regs[15][0] ),
    .Y(net1813));
 sky130_as_sc_hs__buff_2 hold1273 (.A(\tholin_riscv.regs[21][0] ),
    .Y(net1814));
 sky130_as_sc_hs__buff_2 hold1274 (.A(\tholin_riscv.regs[6][0] ),
    .Y(net1815));
 sky130_as_sc_hs__buff_2 hold1275 (.A(\tholin_riscv.regs[5][0] ),
    .Y(net1816));
 sky130_as_sc_hs__buff_2 hold1276 (.A(\tholin_riscv.regs[11][0] ),
    .Y(net1817));
 sky130_as_sc_hs__buff_2 hold1277 (.A(\tholin_riscv.regs[22][0] ),
    .Y(net1818));
 sky130_as_sc_hs__buff_2 hold1278 (.A(\tholin_riscv.regs[8][0] ),
    .Y(net1819));
 sky130_as_sc_hs__buff_2 hold1279 (.A(\tholin_riscv.regs[31][0] ),
    .Y(net1820));
 sky130_as_sc_hs__buff_2 hold128 (.A(net1807),
    .Y(net669));
 sky130_as_sc_hs__buff_2 hold1280 (.A(\tholin_riscv.regs[2][0] ),
    .Y(net1821));
 sky130_as_sc_hs__buff_2 hold1281 (.A(\tholin_riscv.regs[19][0] ),
    .Y(net1822));
 sky130_as_sc_hs__buff_2 hold1282 (.A(\tholin_riscv.regs[23][0] ),
    .Y(net1823));
 sky130_as_sc_hs__buff_2 hold1283 (.A(\tholin_riscv.regs[1][0] ),
    .Y(net1824));
 sky130_as_sc_hs__buff_2 hold1284 (.A(\tholin_riscv.regs[16][0] ),
    .Y(net1825));
 sky130_as_sc_hs__buff_2 hold1285 (.A(\tholin_riscv.regs[14][0] ),
    .Y(net1826));
 sky130_as_sc_hs__buff_2 hold1286 (.A(\tholin_riscv.regs[26][0] ),
    .Y(net1827));
 sky130_as_sc_hs__buff_2 hold1287 (.A(\tholin_riscv.regs[18][0] ),
    .Y(net1828));
 sky130_as_sc_hs__buff_2 hold1288 (.A(\tholin_riscv.regs[27][0] ),
    .Y(net1829));
 sky130_as_sc_hs__buff_2 hold1289 (.A(\tholin_riscv.uart.divisor[11] ),
    .Y(net1830));
 sky130_as_sc_hs__buff_2 hold129 (.A(_19408_),
    .Y(net670));
 sky130_as_sc_hs__buff_2 hold1290 (.A(\tholin_riscv.regs[4][0] ),
    .Y(net1831));
 sky130_as_sc_hs__buff_2 hold1291 (.A(\tholin_riscv.Bimm[9] ),
    .Y(net1832));
 sky130_as_sc_hs__buff_2 hold13 (.A(net1723),
    .Y(net554));
 sky130_as_sc_hs__buff_2 hold130 (.A(_01689_),
    .Y(net671));
 sky130_as_sc_hs__buff_2 hold131 (.A(net1814),
    .Y(net672));
 sky130_as_sc_hs__buff_2 hold132 (.A(_14222_),
    .Y(net673));
 sky130_as_sc_hs__buff_2 hold133 (.A(_00791_),
    .Y(net674));
 sky130_as_sc_hs__buff_2 hold134 (.A(net1808),
    .Y(net675));
 sky130_as_sc_hs__buff_2 hold135 (.A(_14486_),
    .Y(net676));
 sky130_as_sc_hs__buff_2 hold136 (.A(_00919_),
    .Y(net677));
 sky130_as_sc_hs__buff_2 hold137 (.A(net1809),
    .Y(net678));
 sky130_as_sc_hs__buff_2 hold138 (.A(_18638_),
    .Y(net679));
 sky130_as_sc_hs__buff_2 hold139 (.A(_01589_),
    .Y(net680));
 sky130_as_sc_hs__buff_2 hold14 (.A(_14796_),
    .Y(net555));
 sky130_as_sc_hs__buff_2 hold140 (.A(net1806),
    .Y(net681));
 sky130_as_sc_hs__buff_2 hold141 (.A(_13484_),
    .Y(net682));
 sky130_as_sc_hs__buff_2 hold142 (.A(_00438_),
    .Y(net683));
 sky130_as_sc_hs__buff_2 hold143 (.A(net1803),
    .Y(net684));
 sky130_as_sc_hs__buff_2 hold144 (.A(_13627_),
    .Y(net685));
 sky130_as_sc_hs__buff_2 hold145 (.A(_00503_),
    .Y(net686));
 sky130_as_sc_hs__buff_2 hold146 (.A(net1813),
    .Y(net687));
 sky130_as_sc_hs__buff_2 hold147 (.A(_13216_),
    .Y(net688));
 sky130_as_sc_hs__buff_2 hold148 (.A(_00278_),
    .Y(net689));
 sky130_as_sc_hs__buff_2 hold149 (.A(net1817),
    .Y(net690));
 sky130_as_sc_hs__buff_2 hold15 (.A(net1725),
    .Y(net556));
 sky130_as_sc_hs__buff_2 hold150 (.A(_12820_),
    .Y(net691));
 sky130_as_sc_hs__buff_2 hold151 (.A(_00117_),
    .Y(net692));
 sky130_as_sc_hs__buff_2 hold152 (.A(net1815),
    .Y(net693));
 sky130_as_sc_hs__buff_2 hold153 (.A(_13561_),
    .Y(net694));
 sky130_as_sc_hs__buff_2 hold154 (.A(_00471_),
    .Y(net695));
 sky130_as_sc_hs__buff_2 hold155 (.A(net1810),
    .Y(net696));
 sky130_as_sc_hs__buff_2 hold156 (.A(_13348_),
    .Y(net697));
 sky130_as_sc_hs__buff_2 hold157 (.A(_00342_),
    .Y(net698));
 sky130_as_sc_hs__buff_2 hold158 (.A(net1818),
    .Y(net699));
 sky130_as_sc_hs__buff_2 hold159 (.A(_14156_),
    .Y(net700));
 sky130_as_sc_hs__buff_2 hold16 (.A(net1727),
    .Y(net557));
 sky130_as_sc_hs__buff_2 hold160 (.A(_00759_),
    .Y(net701));
 sky130_as_sc_hs__buff_2 hold161 (.A(net1819),
    .Y(net702));
 sky130_as_sc_hs__buff_2 hold162 (.A(_12886_),
    .Y(net703));
 sky130_as_sc_hs__buff_2 hold163 (.A(_00149_),
    .Y(net704));
 sky130_as_sc_hs__buff_2 hold164 (.A(net1811),
    .Y(net705));
 sky130_as_sc_hs__buff_2 hold165 (.A(_13414_),
    .Y(net706));
 sky130_as_sc_hs__buff_2 hold166 (.A(_00374_),
    .Y(net707));
 sky130_as_sc_hs__buff_2 hold167 (.A(net1821),
    .Y(net708));
 sky130_as_sc_hs__buff_2 hold168 (.A(_13693_),
    .Y(net709));
 sky130_as_sc_hs__buff_2 hold169 (.A(_00535_),
    .Y(net710));
 sky130_as_sc_hs__buff_2 hold17 (.A(_15126_),
    .Y(net558));
 sky130_as_sc_hs__buff_2 hold170 (.A(net1825),
    .Y(net711));
 sky130_as_sc_hs__buff_2 hold171 (.A(_12684_),
    .Y(net712));
 sky130_as_sc_hs__buff_2 hold172 (.A(_00053_),
    .Y(net713));
 sky130_as_sc_hs__buff_2 hold173 (.A(net1823),
    .Y(net714));
 sky130_as_sc_hs__buff_2 hold174 (.A(_14090_),
    .Y(net715));
 sky130_as_sc_hs__buff_2 hold175 (.A(_00727_),
    .Y(net716));
 sky130_as_sc_hs__buff_2 hold176 (.A(\tholin_riscv.spi.counter[4] ),
    .Y(net717));
 sky130_as_sc_hs__buff_2 hold177 (.A(_19527_),
    .Y(net718));
 sky130_as_sc_hs__buff_2 hold178 (.A(_15160_),
    .Y(net719));
 sky130_as_sc_hs__buff_2 hold179 (.A(net1816),
    .Y(net720));
 sky130_as_sc_hs__buff_2 hold18 (.A(net1729),
    .Y(net559));
 sky130_as_sc_hs__buff_2 hold180 (.A(_14288_),
    .Y(net721));
 sky130_as_sc_hs__buff_2 hold181 (.A(_00823_),
    .Y(net722));
 sky130_as_sc_hs__buff_2 hold182 (.A(net1824),
    .Y(net723));
 sky130_as_sc_hs__buff_2 hold183 (.A(_18711_),
    .Y(net724));
 sky130_as_sc_hs__buff_2 hold184 (.A(_01622_),
    .Y(net725));
 sky130_as_sc_hs__buff_2 hold185 (.A(net1822),
    .Y(net726));
 sky130_as_sc_hs__buff_2 hold186 (.A(_14354_),
    .Y(net727));
 sky130_as_sc_hs__buff_2 hold187 (.A(_00855_),
    .Y(net728));
 sky130_as_sc_hs__buff_2 hold188 (.A(net1828),
    .Y(net729));
 sky130_as_sc_hs__buff_2 hold189 (.A(_13083_),
    .Y(net730));
 sky130_as_sc_hs__buff_2 hold19 (.A(net1731),
    .Y(net560));
 sky130_as_sc_hs__buff_2 hold190 (.A(_00214_),
    .Y(net731));
 sky130_as_sc_hs__buff_2 hold191 (.A(net1827),
    .Y(net732));
 sky130_as_sc_hs__buff_2 hold192 (.A(_13892_),
    .Y(net733));
 sky130_as_sc_hs__buff_2 hold193 (.A(_00631_),
    .Y(net734));
 sky130_as_sc_hs__buff_2 hold194 (.A(net1820),
    .Y(net735));
 sky130_as_sc_hs__buff_2 hold195 (.A(_06180_),
    .Y(net736));
 sky130_as_sc_hs__buff_2 hold196 (.A(_00021_),
    .Y(net737));
 sky130_as_sc_hs__buff_2 hold197 (.A(net1826),
    .Y(net738));
 sky130_as_sc_hs__buff_2 hold198 (.A(_12753_),
    .Y(net739));
 sky130_as_sc_hs__buff_2 hold199 (.A(_00085_),
    .Y(net740));
 sky130_as_sc_hs__buff_2 hold2 (.A(net1712),
    .Y(net543));
 sky130_as_sc_hs__buff_2 hold20 (.A(_15114_),
    .Y(net561));
 sky130_as_sc_hs__buff_2 hold200 (.A(net1829),
    .Y(net741));
 sky130_as_sc_hs__buff_2 hold201 (.A(_13826_),
    .Y(net742));
 sky130_as_sc_hs__buff_2 hold202 (.A(_00599_),
    .Y(net743));
 sky130_as_sc_hs__buff_2 hold203 (.A(net1831),
    .Y(net744));
 sky130_as_sc_hs__buff_2 hold204 (.A(_14420_),
    .Y(net745));
 sky130_as_sc_hs__buff_2 hold205 (.A(_00887_),
    .Y(net746));
 sky130_as_sc_hs__buff_2 hold206 (.A(\tholin_riscv.tmr0_pre_ctr[1] ),
    .Y(net747));
 sky130_as_sc_hs__buff_2 hold207 (.A(_17127_),
    .Y(net748));
 sky130_as_sc_hs__buff_2 hold208 (.A(_17128_),
    .Y(net749));
 sky130_as_sc_hs__buff_2 hold209 (.A(_01313_),
    .Y(net750));
 sky130_as_sc_hs__buff_2 hold21 (.A(net1733),
    .Y(net562));
 sky130_as_sc_hs__buff_2 hold210 (.A(\tholin_riscv.spi.divisor[6] ),
    .Y(net751));
 sky130_as_sc_hs__buff_2 hold211 (.A(_15268_),
    .Y(net752));
 sky130_as_sc_hs__buff_2 hold212 (.A(_01083_),
    .Y(net753));
 sky130_as_sc_hs__buff_2 hold213 (.A(net1709),
    .Y(net754));
 sky130_as_sc_hs__buff_2 hold214 (.A(_14927_),
    .Y(net755));
 sky130_as_sc_hs__buff_2 hold215 (.A(_01001_),
    .Y(net756));
 sky130_as_sc_hs__buff_2 hold216 (.A(\tholin_riscv.int_enabled ),
    .Y(net757));
 sky130_as_sc_hs__buff_2 hold217 (.A(_16417_),
    .Y(net758));
 sky130_as_sc_hs__buff_2 hold218 (.A(_01228_),
    .Y(net759));
 sky130_as_sc_hs__buff_2 hold219 (.A(\tholin_riscv.tmr0_pre_ctr[25] ),
    .Y(net760));
 sky130_as_sc_hs__buff_2 hold22 (.A(\tholin_riscv.spi.data_in_buff[5] ),
    .Y(net563));
 sky130_as_sc_hs__buff_2 hold220 (.A(_17224_),
    .Y(net761));
 sky130_as_sc_hs__buff_2 hold221 (.A(_17225_),
    .Y(net762));
 sky130_as_sc_hs__buff_2 hold222 (.A(_01337_),
    .Y(net763));
 sky130_as_sc_hs__buff_2 hold223 (.A(\tholin_riscv.tmr1_pre_ctr[25] ),
    .Y(net764));
 sky130_as_sc_hs__buff_2 hold224 (.A(_16334_),
    .Y(net765));
 sky130_as_sc_hs__buff_2 hold225 (.A(_16335_),
    .Y(net766));
 sky130_as_sc_hs__buff_2 hold226 (.A(_01217_),
    .Y(net767));
 sky130_as_sc_hs__buff_2 hold227 (.A(\tholin_riscv.tmr1_pre_ctr[1] ),
    .Y(net768));
 sky130_as_sc_hs__buff_2 hold228 (.A(_16237_),
    .Y(net769));
 sky130_as_sc_hs__buff_2 hold229 (.A(_16238_),
    .Y(net770));
 sky130_as_sc_hs__buff_2 hold23 (.A(_15120_),
    .Y(net564));
 sky130_as_sc_hs__buff_2 hold230 (.A(_01193_),
    .Y(net771));
 sky130_as_sc_hs__buff_2 hold231 (.A(\tholin_riscv.spi.divisor[3] ),
    .Y(net772));
 sky130_as_sc_hs__buff_2 hold232 (.A(_15259_),
    .Y(net773));
 sky130_as_sc_hs__buff_2 hold233 (.A(_01080_),
    .Y(net774));
 sky130_as_sc_hs__buff_2 hold234 (.A(\tholin_riscv.tmr0_pre_ctr[30] ),
    .Y(net775));
 sky130_as_sc_hs__buff_2 hold235 (.A(_17096_),
    .Y(net776));
 sky130_as_sc_hs__buff_2 hold236 (.A(_17253_),
    .Y(net777));
 sky130_as_sc_hs__buff_2 hold237 (.A(_01342_),
    .Y(net778));
 sky130_as_sc_hs__buff_2 hold238 (.A(\tholin_riscv.tmr0[0] ),
    .Y(net779));
 sky130_as_sc_hs__buff_2 hold239 (.A(_18136_),
    .Y(net780));
 sky130_as_sc_hs__buff_2 hold24 (.A(net1742),
    .Y(net565));
 sky130_as_sc_hs__buff_2 hold240 (.A(_18138_),
    .Y(net781));
 sky130_as_sc_hs__buff_2 hold241 (.A(_01505_),
    .Y(net782));
 sky130_as_sc_hs__buff_2 hold242 (.A(\tholin_riscv.tmr1[0] ),
    .Y(net783));
 sky130_as_sc_hs__buff_2 hold243 (.A(_17405_),
    .Y(net784));
 sky130_as_sc_hs__buff_2 hold244 (.A(_17407_),
    .Y(net785));
 sky130_as_sc_hs__buff_2 hold245 (.A(_01345_),
    .Y(net786));
 sky130_as_sc_hs__buff_2 hold246 (.A(net1799),
    .Y(net787));
 sky130_as_sc_hs__buff_2 hold247 (.A(_16206_),
    .Y(net788));
 sky130_as_sc_hs__buff_2 hold248 (.A(_16363_),
    .Y(net789));
 sky130_as_sc_hs__buff_2 hold249 (.A(\tholin_riscv.tmr0[7] ),
    .Y(net790));
 sky130_as_sc_hs__buff_2 hold25 (.A(net614),
    .Y(net566));
 sky130_as_sc_hs__buff_2 hold250 (.A(_19713_),
    .Y(net791));
 sky130_as_sc_hs__buff_2 hold251 (.A(_18188_),
    .Y(net792));
 sky130_as_sc_hs__buff_2 hold252 (.A(_18192_),
    .Y(net793));
 sky130_as_sc_hs__buff_2 hold253 (.A(\tholin_riscv.tmr0[13] ),
    .Y(net794));
 sky130_as_sc_hs__buff_2 hold254 (.A(_19707_),
    .Y(net795));
 sky130_as_sc_hs__buff_2 hold255 (.A(_18242_),
    .Y(net796));
 sky130_as_sc_hs__buff_2 hold256 (.A(_18246_),
    .Y(net797));
 sky130_as_sc_hs__buff_2 hold257 (.A(\tholin_riscv.tmr1[13] ),
    .Y(net798));
 sky130_as_sc_hs__buff_2 hold258 (.A(_19734_),
    .Y(net799));
 sky130_as_sc_hs__buff_2 hold259 (.A(_17511_),
    .Y(net800));
 sky130_as_sc_hs__buff_2 hold26 (.A(_14805_),
    .Y(net567));
 sky130_as_sc_hs__buff_2 hold260 (.A(_17515_),
    .Y(net801));
 sky130_as_sc_hs__buff_2 hold261 (.A(\tholin_riscv.tmr1[4] ),
    .Y(net802));
 sky130_as_sc_hs__buff_2 hold262 (.A(_19743_),
    .Y(net803));
 sky130_as_sc_hs__buff_2 hold263 (.A(_17430_),
    .Y(net804));
 sky130_as_sc_hs__buff_2 hold264 (.A(_17434_),
    .Y(net805));
 sky130_as_sc_hs__buff_2 hold265 (.A(\tholin_riscv.tmr0[4] ),
    .Y(net806));
 sky130_as_sc_hs__buff_2 hold266 (.A(_19716_),
    .Y(net807));
 sky130_as_sc_hs__buff_2 hold267 (.A(_18161_),
    .Y(net808));
 sky130_as_sc_hs__buff_2 hold268 (.A(_18165_),
    .Y(net809));
 sky130_as_sc_hs__buff_2 hold269 (.A(\tholin_riscv.tmr1_pre_ctr[23] ),
    .Y(net810));
 sky130_as_sc_hs__buff_2 hold27 (.A(_00978_),
    .Y(net568));
 sky130_as_sc_hs__buff_2 hold270 (.A(_16324_),
    .Y(net811));
 sky130_as_sc_hs__buff_2 hold271 (.A(_16325_),
    .Y(net812));
 sky130_as_sc_hs__buff_2 hold272 (.A(_01215_),
    .Y(net813));
 sky130_as_sc_hs__buff_2 hold273 (.A(\tholin_riscv.tmr1[10] ),
    .Y(net814));
 sky130_as_sc_hs__buff_2 hold274 (.A(_19737_),
    .Y(net815));
 sky130_as_sc_hs__buff_2 hold275 (.A(_17484_),
    .Y(net816));
 sky130_as_sc_hs__buff_2 hold276 (.A(_17488_),
    .Y(net817));
 sky130_as_sc_hs__buff_2 hold277 (.A(\tholin_riscv.tmr1[22] ),
    .Y(net818));
 sky130_as_sc_hs__buff_2 hold278 (.A(_19687_),
    .Y(net819));
 sky130_as_sc_hs__buff_2 hold279 (.A(_17591_),
    .Y(net820));
 sky130_as_sc_hs__buff_2 hold28 (.A(\tholin_riscv.spi.data_in_buff[1] ),
    .Y(net569));
 sky130_as_sc_hs__buff_2 hold280 (.A(_17595_),
    .Y(net821));
 sky130_as_sc_hs__buff_2 hold281 (.A(\tholin_riscv.tmr1_pre_ctr[4] ),
    .Y(net822));
 sky130_as_sc_hs__buff_2 hold282 (.A(_16226_),
    .Y(net823));
 sky130_as_sc_hs__buff_2 hold283 (.A(_16227_),
    .Y(net824));
 sky130_as_sc_hs__buff_2 hold284 (.A(_01196_),
    .Y(net825));
 sky130_as_sc_hs__buff_2 hold285 (.A(\tholin_riscv.tmr0[25] ),
    .Y(net826));
 sky130_as_sc_hs__buff_2 hold286 (.A(_19700_),
    .Y(net827));
 sky130_as_sc_hs__buff_2 hold287 (.A(_18347_),
    .Y(net828));
 sky130_as_sc_hs__buff_2 hold288 (.A(_18351_),
    .Y(net829));
 sky130_as_sc_hs__buff_2 hold289 (.A(\tholin_riscv.tmr1[16] ),
    .Y(net830));
 sky130_as_sc_hs__buff_2 hold29 (.A(_15108_),
    .Y(net570));
 sky130_as_sc_hs__buff_2 hold290 (.A(_19731_),
    .Y(net831));
 sky130_as_sc_hs__buff_2 hold291 (.A(_17538_),
    .Y(net832));
 sky130_as_sc_hs__buff_2 hold292 (.A(_17542_),
    .Y(net833));
 sky130_as_sc_hs__buff_2 hold293 (.A(_01360_),
    .Y(net834));
 sky130_as_sc_hs__buff_2 hold294 (.A(\tholin_riscv.tmr0[19] ),
    .Y(net835));
 sky130_as_sc_hs__buff_2 hold295 (.A(_19701_),
    .Y(net836));
 sky130_as_sc_hs__buff_2 hold296 (.A(_18296_),
    .Y(net837));
 sky130_as_sc_hs__buff_2 hold297 (.A(_18300_),
    .Y(net838));
 sky130_as_sc_hs__buff_2 hold298 (.A(\tholin_riscv.tmr1[19] ),
    .Y(net839));
 sky130_as_sc_hs__buff_2 hold299 (.A(_19728_),
    .Y(net840));
 sky130_as_sc_hs__buff_2 hold3 (.A(\tholin_riscv.tmr0_pre_ctr[0] ),
    .Y(net544));
 sky130_as_sc_hs__buff_2 hold30 (.A(net1767),
    .Y(net571));
 sky130_as_sc_hs__buff_2 hold300 (.A(_17565_),
    .Y(net841));
 sky130_as_sc_hs__buff_2 hold301 (.A(_17569_),
    .Y(net842));
 sky130_as_sc_hs__buff_2 hold302 (.A(\tholin_riscv.tmr1_pre_ctr[13] ),
    .Y(net843));
 sky130_as_sc_hs__buff_2 hold303 (.A(_16220_),
    .Y(net844));
 sky130_as_sc_hs__buff_2 hold304 (.A(_16221_),
    .Y(net845));
 sky130_as_sc_hs__buff_2 hold305 (.A(_01205_),
    .Y(net846));
 sky130_as_sc_hs__buff_2 hold306 (.A(\tholin_riscv.tmr0[10] ),
    .Y(net847));
 sky130_as_sc_hs__buff_2 hold307 (.A(_19710_),
    .Y(net848));
 sky130_as_sc_hs__buff_2 hold308 (.A(_18215_),
    .Y(net849));
 sky130_as_sc_hs__buff_2 hold309 (.A(_18219_),
    .Y(net850));
 sky130_as_sc_hs__buff_2 hold31 (.A(\tholin_riscv.spi.data_in_buff[2] ),
    .Y(net572));
 sky130_as_sc_hs__buff_2 hold310 (.A(\tholin_riscv.tmr1_pre_ctr[5] ),
    .Y(net851));
 sky130_as_sc_hs__buff_2 hold311 (.A(_16246_),
    .Y(net852));
 sky130_as_sc_hs__buff_2 hold312 (.A(_16247_),
    .Y(net853));
 sky130_as_sc_hs__buff_2 hold313 (.A(_01197_),
    .Y(net854));
 sky130_as_sc_hs__buff_2 hold314 (.A(\tholin_riscv.tmr1[7] ),
    .Y(net855));
 sky130_as_sc_hs__buff_2 hold315 (.A(_19740_),
    .Y(net856));
 sky130_as_sc_hs__buff_2 hold316 (.A(_17457_),
    .Y(net857));
 sky130_as_sc_hs__buff_2 hold317 (.A(_17461_),
    .Y(net858));
 sky130_as_sc_hs__buff_2 hold318 (.A(\tholin_riscv.tmr1_pre_ctr[16] ),
    .Y(net859));
 sky130_as_sc_hs__buff_2 hold319 (.A(_16295_),
    .Y(net860));
 sky130_as_sc_hs__buff_2 hold32 (.A(_15111_),
    .Y(net573));
 sky130_as_sc_hs__buff_2 hold320 (.A(_16296_),
    .Y(net861));
 sky130_as_sc_hs__buff_2 hold321 (.A(_01208_),
    .Y(net862));
 sky130_as_sc_hs__buff_2 hold322 (.A(\tholin_riscv.tmr1_pre_ctr[19] ),
    .Y(net863));
 sky130_as_sc_hs__buff_2 hold323 (.A(_16214_),
    .Y(net864));
 sky130_as_sc_hs__buff_2 hold324 (.A(_16215_),
    .Y(net865));
 sky130_as_sc_hs__buff_2 hold325 (.A(_01211_),
    .Y(net866));
 sky130_as_sc_hs__buff_2 hold326 (.A(\tholin_riscv.tmr1_pre_ctr[17] ),
    .Y(net867));
 sky130_as_sc_hs__buff_2 hold327 (.A(_16300_),
    .Y(net868));
 sky130_as_sc_hs__buff_2 hold328 (.A(_16301_),
    .Y(net869));
 sky130_as_sc_hs__buff_2 hold329 (.A(_01209_),
    .Y(net870));
 sky130_as_sc_hs__buff_2 hold33 (.A(net1739),
    .Y(net574));
 sky130_as_sc_hs__buff_2 hold330 (.A(\tholin_riscv.tmr1[25] ),
    .Y(net871));
 sky130_as_sc_hs__buff_2 hold331 (.A(_19727_),
    .Y(net872));
 sky130_as_sc_hs__buff_2 hold332 (.A(_17616_),
    .Y(net873));
 sky130_as_sc_hs__buff_2 hold333 (.A(_17620_),
    .Y(net874));
 sky130_as_sc_hs__buff_2 hold334 (.A(\tholin_riscv.tmr0[16] ),
    .Y(net875));
 sky130_as_sc_hs__buff_2 hold335 (.A(_19704_),
    .Y(net876));
 sky130_as_sc_hs__buff_2 hold336 (.A(_18269_),
    .Y(net877));
 sky130_as_sc_hs__buff_2 hold337 (.A(_18273_),
    .Y(net878));
 sky130_as_sc_hs__buff_2 hold338 (.A(_01520_),
    .Y(net879));
 sky130_as_sc_hs__buff_2 hold339 (.A(\tholin_riscv.tmr0_pre_ctr[5] ),
    .Y(net880));
 sky130_as_sc_hs__buff_2 hold34 (.A(\tholin_riscv.uart.receive_buff[3] ),
    .Y(net575));
 sky130_as_sc_hs__buff_2 hold340 (.A(_17136_),
    .Y(net881));
 sky130_as_sc_hs__buff_2 hold341 (.A(_17137_),
    .Y(net882));
 sky130_as_sc_hs__buff_2 hold342 (.A(_01317_),
    .Y(net883));
 sky130_as_sc_hs__buff_2 hold343 (.A(\tholin_riscv.tmr0_pre_ctr[2] ),
    .Y(net884));
 sky130_as_sc_hs__buff_2 hold344 (.A(_17123_),
    .Y(net885));
 sky130_as_sc_hs__buff_2 hold345 (.A(_17124_),
    .Y(net886));
 sky130_as_sc_hs__buff_2 hold346 (.A(_01314_),
    .Y(net887));
 sky130_as_sc_hs__buff_2 hold347 (.A(\tholin_riscv.tmr1[30] ),
    .Y(net888));
 sky130_as_sc_hs__buff_2 hold348 (.A(_19722_),
    .Y(net889));
 sky130_as_sc_hs__buff_2 hold349 (.A(_17658_),
    .Y(net890));
 sky130_as_sc_hs__buff_2 hold35 (.A(_14793_),
    .Y(net576));
 sky130_as_sc_hs__buff_2 hold350 (.A(\tholin_riscv.tmr0_pre_ctr[21] ),
    .Y(net891));
 sky130_as_sc_hs__buff_2 hold351 (.A(_17204_),
    .Y(net892));
 sky130_as_sc_hs__buff_2 hold352 (.A(_17205_),
    .Y(net893));
 sky130_as_sc_hs__buff_2 hold353 (.A(_01333_),
    .Y(net894));
 sky130_as_sc_hs__buff_2 hold354 (.A(\tholin_riscv.tmr1_pre_ctr[18] ),
    .Y(net895));
 sky130_as_sc_hs__buff_2 hold355 (.A(_16304_),
    .Y(net896));
 sky130_as_sc_hs__buff_2 hold356 (.A(_16305_),
    .Y(net897));
 sky130_as_sc_hs__buff_2 hold357 (.A(_01210_),
    .Y(net898));
 sky130_as_sc_hs__buff_2 hold358 (.A(\tholin_riscv.tmr0_pre_ctr[18] ),
    .Y(net899));
 sky130_as_sc_hs__buff_2 hold359 (.A(_17194_),
    .Y(net900));
 sky130_as_sc_hs__buff_2 hold36 (.A(net1749),
    .Y(net577));
 sky130_as_sc_hs__buff_2 hold360 (.A(_17195_),
    .Y(net901));
 sky130_as_sc_hs__buff_2 hold361 (.A(_01330_),
    .Y(net902));
 sky130_as_sc_hs__buff_2 hold362 (.A(\tholin_riscv.tmr1_pre_ctr[22] ),
    .Y(net903));
 sky130_as_sc_hs__buff_2 hold363 (.A(_16319_),
    .Y(net904));
 sky130_as_sc_hs__buff_2 hold364 (.A(_16320_),
    .Y(net905));
 sky130_as_sc_hs__buff_2 hold365 (.A(_01214_),
    .Y(net906));
 sky130_as_sc_hs__buff_2 hold366 (.A(\tholin_riscv.tmr1_pre_ctr[15] ),
    .Y(net907));
 sky130_as_sc_hs__buff_2 hold367 (.A(_16289_),
    .Y(net908));
 sky130_as_sc_hs__buff_2 hold368 (.A(_16290_),
    .Y(net909));
 sky130_as_sc_hs__buff_2 hold369 (.A(_01207_),
    .Y(net910));
 sky130_as_sc_hs__buff_2 hold37 (.A(\tholin_riscv.spi.data_in_buff[4] ),
    .Y(net578));
 sky130_as_sc_hs__buff_2 hold370 (.A(\tholin_riscv.tmr0_pre_ctr[20] ),
    .Y(net911));
 sky130_as_sc_hs__buff_2 hold371 (.A(_17101_),
    .Y(net912));
 sky130_as_sc_hs__buff_2 hold372 (.A(_17102_),
    .Y(net913));
 sky130_as_sc_hs__buff_2 hold373 (.A(_01332_),
    .Y(net914));
 sky130_as_sc_hs__buff_2 hold374 (.A(\tholin_riscv.tmr1_pre_ctr[24] ),
    .Y(net915));
 sky130_as_sc_hs__buff_2 hold375 (.A(_16329_),
    .Y(net916));
 sky130_as_sc_hs__buff_2 hold376 (.A(_16330_),
    .Y(net917));
 sky130_as_sc_hs__buff_2 hold377 (.A(_01216_),
    .Y(net918));
 sky130_as_sc_hs__buff_2 hold378 (.A(\tholin_riscv.tmr0_pre_ctr[13] ),
    .Y(net919));
 sky130_as_sc_hs__buff_2 hold379 (.A(_17110_),
    .Y(net920));
 sky130_as_sc_hs__buff_2 hold38 (.A(_15117_),
    .Y(net579));
 sky130_as_sc_hs__buff_2 hold380 (.A(_17111_),
    .Y(net921));
 sky130_as_sc_hs__buff_2 hold381 (.A(_01325_),
    .Y(net922));
 sky130_as_sc_hs__buff_2 hold382 (.A(\tholin_riscv.tmr0[28] ),
    .Y(net923));
 sky130_as_sc_hs__buff_2 hold383 (.A(_19697_),
    .Y(net924));
 sky130_as_sc_hs__buff_2 hold384 (.A(_18372_),
    .Y(net925));
 sky130_as_sc_hs__buff_2 hold385 (.A(_18376_),
    .Y(net926));
 sky130_as_sc_hs__buff_2 hold386 (.A(\tholin_riscv.tmr0_pre_ctr[7] ),
    .Y(net927));
 sky130_as_sc_hs__buff_2 hold387 (.A(_17147_),
    .Y(net928));
 sky130_as_sc_hs__buff_2 hold388 (.A(_17148_),
    .Y(net929));
 sky130_as_sc_hs__buff_2 hold389 (.A(_01319_),
    .Y(net930));
 sky130_as_sc_hs__buff_2 hold39 (.A(net1764),
    .Y(net580));
 sky130_as_sc_hs__buff_2 hold390 (.A(\tholin_riscv.tmr0_pre_ctr[22] ),
    .Y(net931));
 sky130_as_sc_hs__buff_2 hold391 (.A(_17209_),
    .Y(net932));
 sky130_as_sc_hs__buff_2 hold392 (.A(_17210_),
    .Y(net933));
 sky130_as_sc_hs__buff_2 hold393 (.A(_01334_),
    .Y(net934));
 sky130_as_sc_hs__buff_2 hold394 (.A(\tholin_riscv.tmr0_pre_ctr[17] ),
    .Y(net935));
 sky130_as_sc_hs__buff_2 hold395 (.A(_17190_),
    .Y(net936));
 sky130_as_sc_hs__buff_2 hold396 (.A(_17191_),
    .Y(net937));
 sky130_as_sc_hs__buff_2 hold397 (.A(_01329_),
    .Y(net938));
 sky130_as_sc_hs__buff_2 hold398 (.A(\tholin_riscv.tmr1_pre_ctr[26] ),
    .Y(net939));
 sky130_as_sc_hs__buff_2 hold399 (.A(_16336_),
    .Y(net940));
 sky130_as_sc_hs__buff_2 hold4 (.A(net1715),
    .Y(net545));
 sky130_as_sc_hs__buff_2 hold40 (.A(net1773),
    .Y(net581));
 sky130_as_sc_hs__buff_2 hold400 (.A(_16337_),
    .Y(net941));
 sky130_as_sc_hs__buff_2 hold401 (.A(_01218_),
    .Y(net942));
 sky130_as_sc_hs__buff_2 hold402 (.A(\tholin_riscv.tmr1_pre_ctr[14] ),
    .Y(net943));
 sky130_as_sc_hs__buff_2 hold403 (.A(_16217_),
    .Y(net944));
 sky130_as_sc_hs__buff_2 hold404 (.A(_16218_),
    .Y(net945));
 sky130_as_sc_hs__buff_2 hold405 (.A(_01206_),
    .Y(net946));
 sky130_as_sc_hs__buff_2 hold406 (.A(\tholin_riscv.tmr1_pre_ctr[9] ),
    .Y(net947));
 sky130_as_sc_hs__buff_2 hold407 (.A(_16267_),
    .Y(net948));
 sky130_as_sc_hs__buff_2 hold408 (.A(_16268_),
    .Y(net949));
 sky130_as_sc_hs__buff_2 hold409 (.A(_01201_),
    .Y(net950));
 sky130_as_sc_hs__buff_2 hold41 (.A(_14917_),
    .Y(net582));
 sky130_as_sc_hs__buff_2 hold410 (.A(\tholin_riscv.tmr1[28] ),
    .Y(net951));
 sky130_as_sc_hs__buff_2 hold411 (.A(_19724_),
    .Y(net952));
 sky130_as_sc_hs__buff_2 hold412 (.A(_17641_),
    .Y(net953));
 sky130_as_sc_hs__buff_2 hold413 (.A(_17645_),
    .Y(net954));
 sky130_as_sc_hs__buff_2 hold414 (.A(\tholin_riscv.tmr0_pre_ctr[29] ),
    .Y(net955));
 sky130_as_sc_hs__buff_2 hold415 (.A(_17247_),
    .Y(net956));
 sky130_as_sc_hs__buff_2 hold416 (.A(_17248_),
    .Y(net957));
 sky130_as_sc_hs__buff_2 hold417 (.A(_01341_),
    .Y(net958));
 sky130_as_sc_hs__buff_2 hold418 (.A(\tholin_riscv.tmr0_pre_ctr[26] ),
    .Y(net959));
 sky130_as_sc_hs__buff_2 hold419 (.A(_17226_),
    .Y(net960));
 sky130_as_sc_hs__buff_2 hold42 (.A(_00999_),
    .Y(net583));
 sky130_as_sc_hs__buff_2 hold420 (.A(_17227_),
    .Y(net961));
 sky130_as_sc_hs__buff_2 hold421 (.A(_01338_),
    .Y(net962));
 sky130_as_sc_hs__buff_2 hold422 (.A(\tholin_riscv.tmr0_pre_ctr[3] ),
    .Y(net963));
 sky130_as_sc_hs__buff_2 hold423 (.A(_17119_),
    .Y(net964));
 sky130_as_sc_hs__buff_2 hold424 (.A(_17120_),
    .Y(net965));
 sky130_as_sc_hs__buff_2 hold425 (.A(_01315_),
    .Y(net966));
 sky130_as_sc_hs__buff_2 hold426 (.A(\tholin_riscv.tmr1_pre_ctr[2] ),
    .Y(net967));
 sky130_as_sc_hs__buff_2 hold427 (.A(_16233_),
    .Y(net968));
 sky130_as_sc_hs__buff_2 hold428 (.A(_16234_),
    .Y(net969));
 sky130_as_sc_hs__buff_2 hold429 (.A(_01194_),
    .Y(net970));
 sky130_as_sc_hs__buff_2 hold43 (.A(\tholin_riscv.uart.receive_buff[6] ),
    .Y(net584));
 sky130_as_sc_hs__buff_2 hold430 (.A(\tholin_riscv.tmr0[22] ),
    .Y(net971));
 sky130_as_sc_hs__buff_2 hold431 (.A(_19688_),
    .Y(net972));
 sky130_as_sc_hs__buff_2 hold432 (.A(_18322_),
    .Y(net973));
 sky130_as_sc_hs__buff_2 hold433 (.A(_18326_),
    .Y(net974));
 sky130_as_sc_hs__buff_2 hold434 (.A(_01526_),
    .Y(net975));
 sky130_as_sc_hs__buff_2 hold435 (.A(\tholin_riscv.tmr0_pre_ctr[11] ),
    .Y(net976));
 sky130_as_sc_hs__buff_2 hold436 (.A(_17167_),
    .Y(net977));
 sky130_as_sc_hs__buff_2 hold437 (.A(_17168_),
    .Y(net978));
 sky130_as_sc_hs__buff_2 hold438 (.A(_01323_),
    .Y(net979));
 sky130_as_sc_hs__buff_2 hold439 (.A(\tholin_riscv.tmr0_pre_ctr[10] ),
    .Y(net980));
 sky130_as_sc_hs__buff_2 hold44 (.A(_14802_),
    .Y(net585));
 sky130_as_sc_hs__buff_2 hold440 (.A(_17162_),
    .Y(net981));
 sky130_as_sc_hs__buff_2 hold441 (.A(_17163_),
    .Y(net982));
 sky130_as_sc_hs__buff_2 hold442 (.A(_01322_),
    .Y(net983));
 sky130_as_sc_hs__buff_2 hold443 (.A(\tholin_riscv.tmr0_pre_ctr[4] ),
    .Y(net984));
 sky130_as_sc_hs__buff_2 hold444 (.A(_17116_),
    .Y(net985));
 sky130_as_sc_hs__buff_2 hold445 (.A(_17117_),
    .Y(net986));
 sky130_as_sc_hs__buff_2 hold446 (.A(_01316_),
    .Y(net987));
 sky130_as_sc_hs__buff_2 hold447 (.A(\tholin_riscv.tmr1_pre_ctr[27] ),
    .Y(net988));
 sky130_as_sc_hs__buff_2 hold448 (.A(_16339_),
    .Y(net989));
 sky130_as_sc_hs__buff_2 hold449 (.A(_16340_),
    .Y(net990));
 sky130_as_sc_hs__buff_2 hold45 (.A(net1758),
    .Y(net586));
 sky130_as_sc_hs__buff_2 hold450 (.A(_01219_),
    .Y(net991));
 sky130_as_sc_hs__buff_2 hold451 (.A(\tholin_riscv.tmr0_pre_ctr[24] ),
    .Y(net992));
 sky130_as_sc_hs__buff_2 hold452 (.A(_17219_),
    .Y(net993));
 sky130_as_sc_hs__buff_2 hold453 (.A(_17220_),
    .Y(net994));
 sky130_as_sc_hs__buff_2 hold454 (.A(_01336_),
    .Y(net995));
 sky130_as_sc_hs__buff_2 hold455 (.A(\tholin_riscv.tmr0_pre_ctr[14] ),
    .Y(net996));
 sky130_as_sc_hs__buff_2 hold456 (.A(_17107_),
    .Y(net997));
 sky130_as_sc_hs__buff_2 hold457 (.A(_17108_),
    .Y(net998));
 sky130_as_sc_hs__buff_2 hold458 (.A(_01326_),
    .Y(net999));
 sky130_as_sc_hs__buff_2 hold459 (.A(\tholin_riscv.tmr1_pre_ctr[6] ),
    .Y(net1000));
 sky130_as_sc_hs__buff_2 hold46 (.A(\tholin_riscv.uart.receive_buff[2] ),
    .Y(net587));
 sky130_as_sc_hs__buff_2 hold460 (.A(_16252_),
    .Y(net1001));
 sky130_as_sc_hs__buff_2 hold461 (.A(_16253_),
    .Y(net1002));
 sky130_as_sc_hs__buff_2 hold462 (.A(_01198_),
    .Y(net1003));
 sky130_as_sc_hs__buff_2 hold463 (.A(\tholin_riscv.tmr0_pre_ctr[8] ),
    .Y(net1004));
 sky130_as_sc_hs__buff_2 hold464 (.A(_17152_),
    .Y(net1005));
 sky130_as_sc_hs__buff_2 hold465 (.A(_17153_),
    .Y(net1006));
 sky130_as_sc_hs__buff_2 hold466 (.A(_01320_),
    .Y(net1007));
 sky130_as_sc_hs__buff_2 hold467 (.A(\tholin_riscv.tmr0_pre_ctr[9] ),
    .Y(net1008));
 sky130_as_sc_hs__buff_2 hold468 (.A(_17157_),
    .Y(net1009));
 sky130_as_sc_hs__buff_2 hold469 (.A(_17158_),
    .Y(net1010));
 sky130_as_sc_hs__buff_2 hold47 (.A(_14790_),
    .Y(net588));
 sky130_as_sc_hs__buff_2 hold470 (.A(_01321_),
    .Y(net1011));
 sky130_as_sc_hs__buff_2 hold471 (.A(\tholin_riscv.tmr1_pre_ctr[11] ),
    .Y(net1012));
 sky130_as_sc_hs__buff_2 hold472 (.A(_16277_),
    .Y(net1013));
 sky130_as_sc_hs__buff_2 hold473 (.A(_16278_),
    .Y(net1014));
 sky130_as_sc_hs__buff_2 hold474 (.A(_01203_),
    .Y(net1015));
 sky130_as_sc_hs__buff_2 hold475 (.A(\tholin_riscv.tmr1_pre_ctr[8] ),
    .Y(net1016));
 sky130_as_sc_hs__buff_2 hold476 (.A(_16262_),
    .Y(net1017));
 sky130_as_sc_hs__buff_2 hold477 (.A(_16263_),
    .Y(net1018));
 sky130_as_sc_hs__buff_2 hold478 (.A(_01200_),
    .Y(net1019));
 sky130_as_sc_hs__buff_2 hold479 (.A(\tholin_riscv.tmr1_pre_ctr[3] ),
    .Y(net1020));
 sky130_as_sc_hs__buff_2 hold48 (.A(net1755),
    .Y(net589));
 sky130_as_sc_hs__buff_2 hold480 (.A(_16229_),
    .Y(net1021));
 sky130_as_sc_hs__buff_2 hold481 (.A(_16230_),
    .Y(net1022));
 sky130_as_sc_hs__buff_2 hold482 (.A(_01195_),
    .Y(net1023));
 sky130_as_sc_hs__buff_2 hold483 (.A(\tholin_riscv.tmr1_pre_ctr[7] ),
    .Y(net1024));
 sky130_as_sc_hs__buff_2 hold484 (.A(_16257_),
    .Y(net1025));
 sky130_as_sc_hs__buff_2 hold485 (.A(_16258_),
    .Y(net1026));
 sky130_as_sc_hs__buff_2 hold486 (.A(_01199_),
    .Y(net1027));
 sky130_as_sc_hs__buff_2 hold487 (.A(\tholin_riscv.tmr0_pre_ctr[12] ),
    .Y(net1028));
 sky130_as_sc_hs__buff_2 hold488 (.A(_17113_),
    .Y(net1029));
 sky130_as_sc_hs__buff_2 hold489 (.A(_17114_),
    .Y(net1030));
 sky130_as_sc_hs__buff_2 hold49 (.A(\tholin_riscv.uart.receive_buff[5] ),
    .Y(net590));
 sky130_as_sc_hs__buff_2 hold490 (.A(_01324_),
    .Y(net1031));
 sky130_as_sc_hs__clkbuff_4 hold491 (.A(net1798),
    .Y(net1032));
 sky130_as_sc_hs__buff_2 hold492 (.A(_15243_),
    .Y(net1033));
 sky130_as_sc_hs__buff_2 hold493 (.A(\tholin_riscv.tmr0_pre_ctr[23] ),
    .Y(net1034));
 sky130_as_sc_hs__buff_2 hold494 (.A(_17214_),
    .Y(net1035));
 sky130_as_sc_hs__buff_2 hold495 (.A(_17215_),
    .Y(net1036));
 sky130_as_sc_hs__buff_2 hold496 (.A(_01335_),
    .Y(net1037));
 sky130_as_sc_hs__buff_2 hold497 (.A(\tholin_riscv.tmr0_pre_ctr[19] ),
    .Y(net1038));
 sky130_as_sc_hs__buff_2 hold498 (.A(_17104_),
    .Y(net1039));
 sky130_as_sc_hs__buff_2 hold499 (.A(_17105_),
    .Y(net1040));
 sky130_as_sc_hs__buff_2 hold5 (.A(net1717),
    .Y(net546));
 sky130_as_sc_hs__buff_2 hold50 (.A(_14799_),
    .Y(net591));
 sky130_as_sc_hs__buff_2 hold500 (.A(_01331_),
    .Y(net1041));
 sky130_as_sc_hs__buff_2 hold501 (.A(\tholin_riscv.tmr0[30] ),
    .Y(net1042));
 sky130_as_sc_hs__buff_2 hold502 (.A(_19695_),
    .Y(net1043));
 sky130_as_sc_hs__buff_2 hold503 (.A(_18389_),
    .Y(net1044));
 sky130_as_sc_hs__buff_2 hold504 (.A(\tholin_riscv.tmr1_pre_ctr[20] ),
    .Y(net1045));
 sky130_as_sc_hs__buff_2 hold505 (.A(_16211_),
    .Y(net1046));
 sky130_as_sc_hs__buff_2 hold506 (.A(_16212_),
    .Y(net1047));
 sky130_as_sc_hs__buff_2 hold507 (.A(_01212_),
    .Y(net1048));
 sky130_as_sc_hs__buff_2 hold508 (.A(\tholin_riscv.tmr1_pre_ctr[10] ),
    .Y(net1049));
 sky130_as_sc_hs__buff_2 hold509 (.A(_16272_),
    .Y(net1050));
 sky130_as_sc_hs__buff_2 hold51 (.A(net1746),
    .Y(net592));
 sky130_as_sc_hs__buff_2 hold510 (.A(_16273_),
    .Y(net1051));
 sky130_as_sc_hs__buff_2 hold511 (.A(_01202_),
    .Y(net1052));
 sky130_as_sc_hs__buff_2 hold512 (.A(\tholin_riscv.tmr0_pre_ctr[16] ),
    .Y(net1053));
 sky130_as_sc_hs__buff_2 hold513 (.A(_17185_),
    .Y(net1054));
 sky130_as_sc_hs__buff_2 hold514 (.A(_17186_),
    .Y(net1055));
 sky130_as_sc_hs__buff_2 hold515 (.A(_01328_),
    .Y(net1056));
 sky130_as_sc_hs__buff_2 hold516 (.A(\tholin_riscv.tmr0_pre_ctr[27] ),
    .Y(net1057));
 sky130_as_sc_hs__buff_2 hold517 (.A(_17229_),
    .Y(net1058));
 sky130_as_sc_hs__buff_2 hold518 (.A(_17230_),
    .Y(net1059));
 sky130_as_sc_hs__buff_2 hold519 (.A(_01339_),
    .Y(net1060));
 sky130_as_sc_hs__buff_2 hold52 (.A(\tholin_riscv.uart.receive_buff[1] ),
    .Y(net593));
 sky130_as_sc_hs__buff_2 hold520 (.A(\tholin_riscv.tmr1_pre_ctr[29] ),
    .Y(net1061));
 sky130_as_sc_hs__buff_2 hold521 (.A(_16357_),
    .Y(net1062));
 sky130_as_sc_hs__buff_2 hold522 (.A(_16358_),
    .Y(net1063));
 sky130_as_sc_hs__buff_2 hold523 (.A(_01221_),
    .Y(net1064));
 sky130_as_sc_hs__buff_2 hold524 (.A(\tholin_riscv.tmr0_pre_ctr[15] ),
    .Y(net1065));
 sky130_as_sc_hs__buff_2 hold525 (.A(_17179_),
    .Y(net1066));
 sky130_as_sc_hs__buff_2 hold526 (.A(_17180_),
    .Y(net1067));
 sky130_as_sc_hs__buff_2 hold527 (.A(_01327_),
    .Y(net1068));
 sky130_as_sc_hs__buff_2 hold528 (.A(\tholin_riscv.tmr1[9] ),
    .Y(net1069));
 sky130_as_sc_hs__buff_2 hold529 (.A(_19738_),
    .Y(net1070));
 sky130_as_sc_hs__buff_2 hold53 (.A(_14787_),
    .Y(net594));
 sky130_as_sc_hs__buff_2 hold530 (.A(_17475_),
    .Y(net1071));
 sky130_as_sc_hs__buff_2 hold531 (.A(_01353_),
    .Y(net1072));
 sky130_as_sc_hs__buff_2 hold532 (.A(\tholin_riscv.tmr0[3] ),
    .Y(net1073));
 sky130_as_sc_hs__buff_2 hold533 (.A(_19717_),
    .Y(net1074));
 sky130_as_sc_hs__buff_2 hold534 (.A(_18152_),
    .Y(net1075));
 sky130_as_sc_hs__buff_2 hold535 (.A(\tholin_riscv.intr_vec[16] ),
    .Y(net1076));
 sky130_as_sc_hs__buff_2 hold536 (.A(_17025_),
    .Y(net1077));
 sky130_as_sc_hs__buff_2 hold537 (.A(_17027_),
    .Y(net1078));
 sky130_as_sc_hs__buff_2 hold538 (.A(\tholin_riscv.div_shifter[16] ),
    .Y(net1079));
 sky130_as_sc_hs__buff_2 hold539 (.A(_15785_),
    .Y(net1080));
 sky130_as_sc_hs__buff_2 hold54 (.A(net1761),
    .Y(net595));
 sky130_as_sc_hs__buff_2 hold540 (.A(_15786_),
    .Y(net1081));
 sky130_as_sc_hs__buff_2 hold541 (.A(\tholin_riscv.tmr0[6] ),
    .Y(net1082));
 sky130_as_sc_hs__buff_2 hold542 (.A(_19714_),
    .Y(net1083));
 sky130_as_sc_hs__buff_2 hold543 (.A(_18179_),
    .Y(net1084));
 sky130_as_sc_hs__buff_2 hold544 (.A(_18183_),
    .Y(net1085));
 sky130_as_sc_hs__buff_2 hold545 (.A(\tholin_riscv.intr_vec[18] ),
    .Y(net1086));
 sky130_as_sc_hs__buff_2 hold546 (.A(_17031_),
    .Y(net1087));
 sky130_as_sc_hs__buff_2 hold547 (.A(_17033_),
    .Y(net1088));
 sky130_as_sc_hs__buff_2 hold548 (.A(\tholin_riscv.tmr1_pre_ctr[28] ),
    .Y(net1089));
 sky130_as_sc_hs__buff_2 hold549 (.A(_16352_),
    .Y(net1090));
 sky130_as_sc_hs__buff_2 hold55 (.A(net1782),
    .Y(net596));
 sky130_as_sc_hs__buff_2 hold550 (.A(_16353_),
    .Y(net1091));
 sky130_as_sc_hs__buff_2 hold551 (.A(_01220_),
    .Y(net1092));
 sky130_as_sc_hs__buff_2 hold552 (.A(\tholin_riscv.div_shifter[15] ),
    .Y(net1093));
 sky130_as_sc_hs__buff_2 hold553 (.A(_15778_),
    .Y(net1094));
 sky130_as_sc_hs__buff_2 hold554 (.A(_15779_),
    .Y(net1095));
 sky130_as_sc_hs__buff_2 hold555 (.A(\tholin_riscv.tmr0_pre_ctr[28] ),
    .Y(net1096));
 sky130_as_sc_hs__buff_2 hold556 (.A(_17242_),
    .Y(net1097));
 sky130_as_sc_hs__buff_2 hold557 (.A(_17243_),
    .Y(net1098));
 sky130_as_sc_hs__buff_2 hold558 (.A(_01340_),
    .Y(net1099));
 sky130_as_sc_hs__buff_2 hold559 (.A(\tholin_riscv.tmr0[9] ),
    .Y(net1100));
 sky130_as_sc_hs__buff_2 hold56 (.A(_18707_),
    .Y(net597));
 sky130_as_sc_hs__buff_2 hold560 (.A(_19711_),
    .Y(net1101));
 sky130_as_sc_hs__buff_2 hold561 (.A(_18206_),
    .Y(net1102));
 sky130_as_sc_hs__buff_2 hold562 (.A(\tholin_riscv.div_shifter[6] ),
    .Y(net1103));
 sky130_as_sc_hs__buff_2 hold563 (.A(_15714_),
    .Y(net1104));
 sky130_as_sc_hs__buff_2 hold564 (.A(_15715_),
    .Y(net1105));
 sky130_as_sc_hs__buff_2 hold565 (.A(\tholin_riscv.intr_vec[13] ),
    .Y(net1106));
 sky130_as_sc_hs__buff_2 hold566 (.A(_17016_),
    .Y(net1107));
 sky130_as_sc_hs__buff_2 hold567 (.A(_17018_),
    .Y(net1108));
 sky130_as_sc_hs__buff_2 hold568 (.A(\tholin_riscv.tmr0_pre_ctr[6] ),
    .Y(net1109));
 sky130_as_sc_hs__buff_2 hold569 (.A(_17142_),
    .Y(net1110));
 sky130_as_sc_hs__buff_2 hold57 (.A(_01621_),
    .Y(net598));
 sky130_as_sc_hs__buff_2 hold570 (.A(_17143_),
    .Y(net1111));
 sky130_as_sc_hs__buff_2 hold571 (.A(_01318_),
    .Y(net1112));
 sky130_as_sc_hs__buff_2 hold572 (.A(\tholin_riscv.intr_vec[21] ),
    .Y(net1113));
 sky130_as_sc_hs__buff_2 hold573 (.A(_17040_),
    .Y(net1114));
 sky130_as_sc_hs__buff_2 hold574 (.A(_17042_),
    .Y(net1115));
 sky130_as_sc_hs__buff_2 hold575 (.A(\tholin_riscv.intr_vec[29] ),
    .Y(net1116));
 sky130_as_sc_hs__buff_2 hold576 (.A(_17064_),
    .Y(net1117));
 sky130_as_sc_hs__buff_2 hold577 (.A(_17066_),
    .Y(net1118));
 sky130_as_sc_hs__buff_2 hold578 (.A(_01311_),
    .Y(net1119));
 sky130_as_sc_hs__buff_2 hold579 (.A(\tholin_riscv.intr_vec[12] ),
    .Y(net1120));
 sky130_as_sc_hs__buff_2 hold58 (.A(\tholin_riscv.spi.data_in_buff[6] ),
    .Y(net599));
 sky130_as_sc_hs__buff_2 hold580 (.A(_17013_),
    .Y(net1121));
 sky130_as_sc_hs__buff_2 hold581 (.A(_17015_),
    .Y(net1122));
 sky130_as_sc_hs__buff_2 hold582 (.A(\tholin_riscv.tmr1_pre_ctr[12] ),
    .Y(net1123));
 sky130_as_sc_hs__buff_2 hold583 (.A(_16223_),
    .Y(net1124));
 sky130_as_sc_hs__buff_2 hold584 (.A(_16224_),
    .Y(net1125));
 sky130_as_sc_hs__buff_2 hold585 (.A(_01204_),
    .Y(net1126));
 sky130_as_sc_hs__buff_2 hold586 (.A(\tholin_riscv.tmr1[3] ),
    .Y(net1127));
 sky130_as_sc_hs__buff_2 hold587 (.A(_19744_),
    .Y(net1128));
 sky130_as_sc_hs__buff_2 hold588 (.A(_17421_),
    .Y(net1129));
 sky130_as_sc_hs__buff_2 hold589 (.A(_17425_),
    .Y(net1130));
 sky130_as_sc_hs__buff_2 hold59 (.A(_15123_),
    .Y(net600));
 sky130_as_sc_hs__buff_2 hold590 (.A(\tholin_riscv.tmr0_pre[0] ),
    .Y(net1131));
 sky130_as_sc_hs__buff_2 hold591 (.A(_17899_),
    .Y(net1132));
 sky130_as_sc_hs__buff_2 hold592 (.A(_17901_),
    .Y(net1133));
 sky130_as_sc_hs__buff_2 hold593 (.A(_01472_),
    .Y(net1134));
 sky130_as_sc_hs__buff_2 hold594 (.A(\tholin_riscv.div_shifter[9] ),
    .Y(net1135));
 sky130_as_sc_hs__buff_2 hold595 (.A(_15736_),
    .Y(net1136));
 sky130_as_sc_hs__buff_2 hold596 (.A(_15737_),
    .Y(net1137));
 sky130_as_sc_hs__buff_2 hold597 (.A(\tholin_riscv.div_shifter[25] ),
    .Y(net1138));
 sky130_as_sc_hs__buff_2 hold598 (.A(_15848_),
    .Y(net1139));
 sky130_as_sc_hs__buff_2 hold599 (.A(_15849_),
    .Y(net1140));
 sky130_as_sc_hs__buff_2 hold6 (.A(net1719),
    .Y(net547));
 sky130_as_sc_hs__buff_2 hold60 (.A(net1770),
    .Y(net601));
 sky130_as_sc_hs__buff_2 hold600 (.A(\tholin_riscv.intr_vec[3] ),
    .Y(net1141));
 sky130_as_sc_hs__buff_2 hold601 (.A(_16986_),
    .Y(net1142));
 sky130_as_sc_hs__buff_2 hold602 (.A(_16988_),
    .Y(net1143));
 sky130_as_sc_hs__buff_2 hold603 (.A(\tholin_riscv.intr_vec[19] ),
    .Y(net1144));
 sky130_as_sc_hs__buff_2 hold604 (.A(_17034_),
    .Y(net1145));
 sky130_as_sc_hs__buff_2 hold605 (.A(_17036_),
    .Y(net1146));
 sky130_as_sc_hs__buff_2 hold606 (.A(\tholin_riscv.intr_vec[7] ),
    .Y(net1147));
 sky130_as_sc_hs__buff_2 hold607 (.A(_16998_),
    .Y(net1148));
 sky130_as_sc_hs__buff_2 hold608 (.A(_17000_),
    .Y(net1149));
 sky130_as_sc_hs__buff_2 hold609 (.A(_01289_),
    .Y(net1150));
 sky130_as_sc_hs__buff_2 hold61 (.A(net1774),
    .Y(net602));
 sky130_as_sc_hs__buff_2 hold610 (.A(\tholin_riscv.intr_vec[24] ),
    .Y(net1151));
 sky130_as_sc_hs__buff_2 hold611 (.A(_17049_),
    .Y(net1152));
 sky130_as_sc_hs__buff_2 hold612 (.A(_17051_),
    .Y(net1153));
 sky130_as_sc_hs__buff_2 hold613 (.A(_01306_),
    .Y(net1154));
 sky130_as_sc_hs__buff_2 hold614 (.A(\tholin_riscv.div_shifter[14] ),
    .Y(net1155));
 sky130_as_sc_hs__buff_2 hold615 (.A(_15771_),
    .Y(net1156));
 sky130_as_sc_hs__buff_2 hold616 (.A(_15772_),
    .Y(net1157));
 sky130_as_sc_hs__buff_2 hold617 (.A(\tholin_riscv.tmr1[6] ),
    .Y(net1158));
 sky130_as_sc_hs__buff_2 hold618 (.A(_19741_),
    .Y(net1159));
 sky130_as_sc_hs__buff_2 hold619 (.A(_17448_),
    .Y(net1160));
 sky130_as_sc_hs__buff_2 hold62 (.A(_18570_),
    .Y(net603));
 sky130_as_sc_hs__buff_2 hold620 (.A(_17452_),
    .Y(net1161));
 sky130_as_sc_hs__buff_2 hold621 (.A(\tholin_riscv.tmr1[27] ),
    .Y(net1162));
 sky130_as_sc_hs__buff_2 hold622 (.A(_19725_),
    .Y(net1163));
 sky130_as_sc_hs__buff_2 hold623 (.A(_17633_),
    .Y(net1164));
 sky130_as_sc_hs__buff_2 hold624 (.A(\tholin_riscv.div_shifter[23] ),
    .Y(net1165));
 sky130_as_sc_hs__buff_2 hold625 (.A(_15834_),
    .Y(net1166));
 sky130_as_sc_hs__buff_2 hold626 (.A(_15835_),
    .Y(net1167));
 sky130_as_sc_hs__clkbuff_4 hold627 (.A(\tholin_riscv.Bimm[2] ),
    .Y(net1168));
 sky130_as_sc_hs__buff_2 hold628 (.A(_15228_),
    .Y(net1169));
 sky130_as_sc_hs__buff_2 hold629 (.A(\tholin_riscv.tmr0[12] ),
    .Y(net1170));
 sky130_as_sc_hs__buff_2 hold63 (.A(_01569_),
    .Y(net604));
 sky130_as_sc_hs__buff_2 hold630 (.A(_19708_),
    .Y(net1171));
 sky130_as_sc_hs__buff_2 hold631 (.A(_18233_),
    .Y(net1172));
 sky130_as_sc_hs__buff_2 hold632 (.A(\tholin_riscv.ret_cycle[0] ),
    .Y(net1173));
 sky130_as_sc_hs__buff_2 hold633 (.A(_16430_),
    .Y(net1174));
 sky130_as_sc_hs__buff_2 hold634 (.A(_16431_),
    .Y(net1175));
 sky130_as_sc_hs__buff_2 hold635 (.A(\tholin_riscv.div_shifter[17] ),
    .Y(net1176));
 sky130_as_sc_hs__buff_2 hold636 (.A(_15792_),
    .Y(net1177));
 sky130_as_sc_hs__buff_2 hold637 (.A(_15793_),
    .Y(net1178));
 sky130_as_sc_hs__buff_2 hold638 (.A(\tholin_riscv.div_shifter[8] ),
    .Y(net1179));
 sky130_as_sc_hs__buff_2 hold639 (.A(_15729_),
    .Y(net1180));
 sky130_as_sc_hs__buff_2 hold64 (.A(\tholin_riscv.uart.receive_buff[0] ),
    .Y(net605));
 sky130_as_sc_hs__buff_2 hold640 (.A(_15730_),
    .Y(net1181));
 sky130_as_sc_hs__buff_2 hold641 (.A(\tholin_riscv.intr_vec[25] ),
    .Y(net1182));
 sky130_as_sc_hs__buff_2 hold642 (.A(_17052_),
    .Y(net1183));
 sky130_as_sc_hs__buff_2 hold643 (.A(_17054_),
    .Y(net1184));
 sky130_as_sc_hs__buff_2 hold644 (.A(\tholin_riscv.tmr1_pre[0] ),
    .Y(net1185));
 sky130_as_sc_hs__buff_2 hold645 (.A(_17802_),
    .Y(net1186));
 sky130_as_sc_hs__buff_2 hold646 (.A(_17804_),
    .Y(net1187));
 sky130_as_sc_hs__buff_2 hold647 (.A(_01440_),
    .Y(net1188));
 sky130_as_sc_hs__buff_2 hold648 (.A(\tholin_riscv.div_shifter[21] ),
    .Y(net1189));
 sky130_as_sc_hs__buff_2 hold649 (.A(_15820_),
    .Y(net1190));
 sky130_as_sc_hs__buff_2 hold65 (.A(_14784_),
    .Y(net606));
 sky130_as_sc_hs__buff_2 hold650 (.A(_15821_),
    .Y(net1191));
 sky130_as_sc_hs__buff_2 hold651 (.A(\tholin_riscv.div_shifter[12] ),
    .Y(net1192));
 sky130_as_sc_hs__buff_2 hold652 (.A(_15757_),
    .Y(net1193));
 sky130_as_sc_hs__buff_2 hold653 (.A(_15758_),
    .Y(net1194));
 sky130_as_sc_hs__buff_2 hold654 (.A(\tholin_riscv.intr_vec[22] ),
    .Y(net1195));
 sky130_as_sc_hs__buff_2 hold655 (.A(_17043_),
    .Y(net1196));
 sky130_as_sc_hs__buff_2 hold656 (.A(_17045_),
    .Y(net1197));
 sky130_as_sc_hs__buff_2 hold657 (.A(\tholin_riscv.tmr0[27] ),
    .Y(net1198));
 sky130_as_sc_hs__buff_2 hold658 (.A(_19698_),
    .Y(net1199));
 sky130_as_sc_hs__buff_2 hold659 (.A(_18364_),
    .Y(net1200));
 sky130_as_sc_hs__buff_2 hold66 (.A(net1752),
    .Y(net607));
 sky130_as_sc_hs__buff_2 hold660 (.A(\tholin_riscv.div_shifter[13] ),
    .Y(net1201));
 sky130_as_sc_hs__buff_2 hold661 (.A(_15764_),
    .Y(net1202));
 sky130_as_sc_hs__buff_2 hold662 (.A(_15765_),
    .Y(net1203));
 sky130_as_sc_hs__buff_2 hold663 (.A(\tholin_riscv.tmr1_pre_ctr[21] ),
    .Y(net1204));
 sky130_as_sc_hs__buff_2 hold664 (.A(_16314_),
    .Y(net1205));
 sky130_as_sc_hs__buff_2 hold665 (.A(_16315_),
    .Y(net1206));
 sky130_as_sc_hs__buff_2 hold666 (.A(_01213_),
    .Y(net1207));
 sky130_as_sc_hs__buff_2 hold667 (.A(\tholin_riscv.div_shifter[28] ),
    .Y(net1208));
 sky130_as_sc_hs__buff_2 hold668 (.A(_15869_),
    .Y(net1209));
 sky130_as_sc_hs__buff_2 hold669 (.A(_15870_),
    .Y(net1210));
 sky130_as_sc_hs__buff_2 hold67 (.A(net1775),
    .Y(net608));
 sky130_as_sc_hs__buff_2 hold670 (.A(\tholin_riscv.tmr0[15] ),
    .Y(net1211));
 sky130_as_sc_hs__buff_2 hold671 (.A(_19705_),
    .Y(net1212));
 sky130_as_sc_hs__buff_2 hold672 (.A(_18260_),
    .Y(net1213));
 sky130_as_sc_hs__buff_2 hold673 (.A(\tholin_riscv.div_shifter[1] ),
    .Y(net1214));
 sky130_as_sc_hs__buff_2 hold674 (.A(_15678_),
    .Y(net1215));
 sky130_as_sc_hs__buff_2 hold675 (.A(_15679_),
    .Y(net1216));
 sky130_as_sc_hs__buff_2 hold676 (.A(\tholin_riscv.intr_vec[2] ),
    .Y(net1217));
 sky130_as_sc_hs__buff_2 hold677 (.A(_16983_),
    .Y(net1218));
 sky130_as_sc_hs__buff_2 hold678 (.A(_16985_),
    .Y(net1219));
 sky130_as_sc_hs__buff_2 hold679 (.A(\tholin_riscv.intr_vec[1] ),
    .Y(net1220));
 sky130_as_sc_hs__buff_2 hold68 (.A(_15139_),
    .Y(net609));
 sky130_as_sc_hs__buff_2 hold680 (.A(_16980_),
    .Y(net1221));
 sky130_as_sc_hs__buff_2 hold681 (.A(_16982_),
    .Y(net1222));
 sky130_as_sc_hs__buff_2 hold682 (.A(\tholin_riscv.div_shifter[26] ),
    .Y(net1223));
 sky130_as_sc_hs__buff_2 hold683 (.A(_15855_),
    .Y(net1224));
 sky130_as_sc_hs__buff_2 hold684 (.A(_15856_),
    .Y(net1225));
 sky130_as_sc_hs__buff_2 hold685 (.A(\tholin_riscv.div_shifter[20] ),
    .Y(net1226));
 sky130_as_sc_hs__buff_2 hold686 (.A(_15813_),
    .Y(net1227));
 sky130_as_sc_hs__buff_2 hold687 (.A(_15814_),
    .Y(net1228));
 sky130_as_sc_hs__buff_2 hold688 (.A(\tholin_riscv.intr_vec[27] ),
    .Y(net1229));
 sky130_as_sc_hs__buff_2 hold689 (.A(_17058_),
    .Y(net1230));
 sky130_as_sc_hs__buff_2 hold69 (.A(_01047_),
    .Y(net610));
 sky130_as_sc_hs__buff_2 hold690 (.A(_17060_),
    .Y(net1231));
 sky130_as_sc_hs__buff_2 hold691 (.A(\tholin_riscv.div_shifter[7] ),
    .Y(net1232));
 sky130_as_sc_hs__buff_2 hold692 (.A(_15722_),
    .Y(net1233));
 sky130_as_sc_hs__buff_2 hold693 (.A(_15723_),
    .Y(net1234));
 sky130_as_sc_hs__buff_2 hold694 (.A(\tholin_riscv.div_shifter[27] ),
    .Y(net1235));
 sky130_as_sc_hs__buff_2 hold695 (.A(_15862_),
    .Y(net1236));
 sky130_as_sc_hs__buff_2 hold696 (.A(_15863_),
    .Y(net1237));
 sky130_as_sc_hs__buff_2 hold697 (.A(\tholin_riscv.spi.dout[0] ),
    .Y(net1238));
 sky130_as_sc_hs__buff_2 hold698 (.A(_15104_),
    .Y(net1239));
 sky130_as_sc_hs__buff_2 hold699 (.A(_15106_),
    .Y(net1240));
 sky130_as_sc_hs__buff_2 hold7 (.A(net1602),
    .Y(net548));
 sky130_as_sc_hs__buff_2 hold70 (.A(net1776),
    .Y(net611));
 sky130_as_sc_hs__buff_2 hold700 (.A(\tholin_riscv.intr_vec[8] ),
    .Y(net1241));
 sky130_as_sc_hs__buff_2 hold701 (.A(_17001_),
    .Y(net1242));
 sky130_as_sc_hs__buff_2 hold702 (.A(_17003_),
    .Y(net1243));
 sky130_as_sc_hs__buff_2 hold703 (.A(_01290_),
    .Y(net1244));
 sky130_as_sc_hs__buff_2 hold704 (.A(\tholin_riscv.intr_vec[11] ),
    .Y(net1245));
 sky130_as_sc_hs__buff_2 hold705 (.A(_17010_),
    .Y(net1246));
 sky130_as_sc_hs__buff_2 hold706 (.A(_17012_),
    .Y(net1247));
 sky130_as_sc_hs__buff_2 hold707 (.A(\tholin_riscv.div_shifter[4] ),
    .Y(net1248));
 sky130_as_sc_hs__buff_2 hold708 (.A(_15700_),
    .Y(net1249));
 sky130_as_sc_hs__buff_2 hold709 (.A(_15701_),
    .Y(net1250));
 sky130_as_sc_hs__buff_2 hold71 (.A(_15253_),
    .Y(net612));
 sky130_as_sc_hs__buff_2 hold710 (.A(\tholin_riscv.tmr1[15] ),
    .Y(net1251));
 sky130_as_sc_hs__buff_2 hold711 (.A(_19732_),
    .Y(net1252));
 sky130_as_sc_hs__buff_2 hold712 (.A(_17529_),
    .Y(net1253));
 sky130_as_sc_hs__buff_2 hold713 (.A(\tholin_riscv.div_shifter[30] ),
    .Y(net1254));
 sky130_as_sc_hs__buff_2 hold714 (.A(_15883_),
    .Y(net1255));
 sky130_as_sc_hs__buff_2 hold715 (.A(_15884_),
    .Y(net1256));
 sky130_as_sc_hs__buff_2 hold716 (.A(\tholin_riscv.tmr1[21] ),
    .Y(net1257));
 sky130_as_sc_hs__buff_2 hold717 (.A(_19685_),
    .Y(net1258));
 sky130_as_sc_hs__buff_2 hold718 (.A(_17583_),
    .Y(net1259));
 sky130_as_sc_hs__buff_4 hold719 (.A(\tholin_riscv.Bimm[1] ),
    .Y(net1260));
 sky130_as_sc_hs__buff_2 hold72 (.A(_01078_),
    .Y(net613));
 sky130_as_sc_hs__buff_2 hold720 (.A(_17924_),
    .Y(net1261));
 sky130_as_sc_hs__buff_2 hold721 (.A(_01480_),
    .Y(net1262));
 sky130_as_sc_hs__buff_2 hold722 (.A(\tholin_riscv.intr_vec[10] ),
    .Y(net1263));
 sky130_as_sc_hs__buff_2 hold723 (.A(_17007_),
    .Y(net1264));
 sky130_as_sc_hs__buff_2 hold724 (.A(_17009_),
    .Y(net1265));
 sky130_as_sc_hs__buff_2 hold725 (.A(\tholin_riscv.intr_vec[5] ),
    .Y(net1266));
 sky130_as_sc_hs__buff_2 hold726 (.A(_16992_),
    .Y(net1267));
 sky130_as_sc_hs__buff_2 hold727 (.A(_16994_),
    .Y(net1268));
 sky130_as_sc_hs__buff_2 hold728 (.A(_01287_),
    .Y(net1269));
 sky130_as_sc_hs__buff_2 hold729 (.A(\tholin_riscv.intr_vec[9] ),
    .Y(net1270));
 sky130_as_sc_hs__buff_2 hold73 (.A(\tholin_riscv.uart.receive_buff[7] ),
    .Y(net614));
 sky130_as_sc_hs__buff_2 hold730 (.A(_17004_),
    .Y(net1271));
 sky130_as_sc_hs__buff_2 hold731 (.A(_17006_),
    .Y(net1272));
 sky130_as_sc_hs__buff_2 hold732 (.A(_01291_),
    .Y(net1273));
 sky130_as_sc_hs__buff_2 hold733 (.A(\tholin_riscv.div_shifter[3] ),
    .Y(net1274));
 sky130_as_sc_hs__buff_2 hold734 (.A(_15693_),
    .Y(net1275));
 sky130_as_sc_hs__buff_2 hold735 (.A(_15694_),
    .Y(net1276));
 sky130_as_sc_hs__buff_2 hold736 (.A(\tholin_riscv.intr_vec[6] ),
    .Y(net1277));
 sky130_as_sc_hs__buff_2 hold737 (.A(_16995_),
    .Y(net1278));
 sky130_as_sc_hs__buff_2 hold738 (.A(_16997_),
    .Y(net1279));
 sky130_as_sc_hs__buff_2 hold739 (.A(\tholin_riscv.div_shifter[29] ),
    .Y(net1280));
 sky130_as_sc_hs__buff_2 hold74 (.A(net566),
    .Y(net615));
 sky130_as_sc_hs__buff_2 hold740 (.A(_15876_),
    .Y(net1281));
 sky130_as_sc_hs__buff_2 hold741 (.A(_15877_),
    .Y(net1282));
 sky130_as_sc_hs__buff_2 hold742 (.A(\tholin_riscv.div_shifter[10] ),
    .Y(net1283));
 sky130_as_sc_hs__buff_2 hold743 (.A(_15743_),
    .Y(net1284));
 sky130_as_sc_hs__buff_2 hold744 (.A(_15744_),
    .Y(net1285));
 sky130_as_sc_hs__buff_2 hold745 (.A(\tholin_riscv.tmr0[21] ),
    .Y(net1286));
 sky130_as_sc_hs__buff_2 hold746 (.A(_19686_),
    .Y(net1287));
 sky130_as_sc_hs__buff_2 hold747 (.A(_18314_),
    .Y(net1288));
 sky130_as_sc_hs__buff_2 hold748 (.A(\tholin_riscv.div_shifter[2] ),
    .Y(net1289));
 sky130_as_sc_hs__buff_2 hold749 (.A(_15686_),
    .Y(net1290));
 sky130_as_sc_hs__buff_2 hold75 (.A(_14967_),
    .Y(net616));
 sky130_as_sc_hs__buff_2 hold750 (.A(_15687_),
    .Y(net1291));
 sky130_as_sc_hs__buff_2 hold751 (.A(\tholin_riscv.div_shifter[19] ),
    .Y(net1292));
 sky130_as_sc_hs__buff_2 hold752 (.A(_15806_),
    .Y(net1293));
 sky130_as_sc_hs__buff_2 hold753 (.A(_15807_),
    .Y(net1294));
 sky130_as_sc_hs__buff_2 hold754 (.A(\tholin_riscv.intr_vec[4] ),
    .Y(net1295));
 sky130_as_sc_hs__buff_2 hold755 (.A(_16989_),
    .Y(net1296));
 sky130_as_sc_hs__buff_2 hold756 (.A(_16991_),
    .Y(net1297));
 sky130_as_sc_hs__buff_2 hold757 (.A(\tholin_riscv.div_shifter[22] ),
    .Y(net1298));
 sky130_as_sc_hs__buff_2 hold758 (.A(_15827_),
    .Y(net1299));
 sky130_as_sc_hs__buff_2 hold759 (.A(_15828_),
    .Y(net1300));
 sky130_as_sc_hs__buff_2 hold76 (.A(_01012_),
    .Y(net617));
 sky130_as_sc_hs__buff_2 hold760 (.A(\tholin_riscv.tmr1[24] ),
    .Y(net1301));
 sky130_as_sc_hs__buff_2 hold761 (.A(_19691_),
    .Y(net1302));
 sky130_as_sc_hs__buff_2 hold762 (.A(_17608_),
    .Y(net1303));
 sky130_as_sc_hs__buff_2 hold763 (.A(\tholin_riscv.div_shifter[24] ),
    .Y(net1304));
 sky130_as_sc_hs__buff_2 hold764 (.A(_15841_),
    .Y(net1305));
 sky130_as_sc_hs__buff_2 hold765 (.A(_15842_),
    .Y(net1306));
 sky130_as_sc_hs__buff_2 hold766 (.A(\tholin_riscv.div_shifter[18] ),
    .Y(net1307));
 sky130_as_sc_hs__buff_2 hold767 (.A(_15799_),
    .Y(net1308));
 sky130_as_sc_hs__buff_2 hold768 (.A(_15800_),
    .Y(net1309));
 sky130_as_sc_hs__buff_2 hold769 (.A(\tholin_riscv.tmr1[12] ),
    .Y(net1310));
 sky130_as_sc_hs__buff_2 hold77 (.A(net1778),
    .Y(net618));
 sky130_as_sc_hs__buff_2 hold770 (.A(_19735_),
    .Y(net1311));
 sky130_as_sc_hs__buff_2 hold771 (.A(_17502_),
    .Y(net1312));
 sky130_as_sc_hs__buff_2 hold772 (.A(\tholin_riscv.div_shifter[11] ),
    .Y(net1313));
 sky130_as_sc_hs__buff_2 hold773 (.A(_15750_),
    .Y(net1314));
 sky130_as_sc_hs__buff_2 hold774 (.A(_15751_),
    .Y(net1315));
 sky130_as_sc_hs__buff_2 hold775 (.A(\tholin_riscv.intr_vec[0] ),
    .Y(net1316));
 sky130_as_sc_hs__buff_2 hold776 (.A(_16977_),
    .Y(net1317));
 sky130_as_sc_hs__buff_2 hold777 (.A(_16979_),
    .Y(net1318));
 sky130_as_sc_hs__buff_2 hold778 (.A(\tholin_riscv.spi.data_out_buff[0] ),
    .Y(net1319));
 sky130_as_sc_hs__buff_2 hold779 (.A(_15162_),
    .Y(net1320));
 sky130_as_sc_hs__buff_2 hold78 (.A(_15256_),
    .Y(net619));
 sky130_as_sc_hs__buff_2 hold780 (.A(_15164_),
    .Y(net1321));
 sky130_as_sc_hs__buff_2 hold781 (.A(_01053_),
    .Y(net1322));
 sky130_as_sc_hs__buff_2 hold782 (.A(\tholin_riscv.tmr0[24] ),
    .Y(net1323));
 sky130_as_sc_hs__buff_2 hold783 (.A(_19692_),
    .Y(net1324));
 sky130_as_sc_hs__buff_2 hold784 (.A(_18339_),
    .Y(net1325));
 sky130_as_sc_hs__buff_2 hold785 (.A(\tholin_riscv.tmr0[18] ),
    .Y(net1326));
 sky130_as_sc_hs__buff_2 hold786 (.A(_19702_),
    .Y(net1327));
 sky130_as_sc_hs__buff_2 hold787 (.A(_18287_),
    .Y(net1328));
 sky130_as_sc_hs__buff_2 hold788 (.A(_18291_),
    .Y(net1329));
 sky130_as_sc_hs__buff_2 hold789 (.A(\tholin_riscv.tmr0_pre[9] ),
    .Y(net1330));
 sky130_as_sc_hs__buff_2 hold79 (.A(_01079_),
    .Y(net620));
 sky130_as_sc_hs__buff_2 hold790 (.A(_17926_),
    .Y(net1331));
 sky130_as_sc_hs__buff_2 hold791 (.A(_17928_),
    .Y(net1332));
 sky130_as_sc_hs__buff_2 hold792 (.A(_01481_),
    .Y(net1333));
 sky130_as_sc_hs__buff_2 hold793 (.A(\tholin_riscv.tmr1[18] ),
    .Y(net1334));
 sky130_as_sc_hs__buff_2 hold794 (.A(_19729_),
    .Y(net1335));
 sky130_as_sc_hs__buff_2 hold795 (.A(_17556_),
    .Y(net1336));
 sky130_as_sc_hs__buff_2 hold796 (.A(\tholin_riscv.intr_vec[15] ),
    .Y(net1337));
 sky130_as_sc_hs__buff_2 hold797 (.A(_17022_),
    .Y(net1338));
 sky130_as_sc_hs__buff_2 hold798 (.A(_17024_),
    .Y(net1339));
 sky130_as_sc_hs__buff_2 hold799 (.A(\tholin_riscv.div_shifter[5] ),
    .Y(net1340));
 sky130_as_sc_hs__buff_2 hold8 (.A(_18579_),
    .Y(net549));
 sky130_as_sc_hs__buff_2 hold80 (.A(net1777),
    .Y(net621));
 sky130_as_sc_hs__buff_2 hold800 (.A(_15707_),
    .Y(net1341));
 sky130_as_sc_hs__buff_2 hold801 (.A(_15708_),
    .Y(net1342));
 sky130_as_sc_hs__buff_2 hold802 (.A(net1794),
    .Y(net1343));
 sky130_as_sc_hs__buff_2 hold803 (.A(_15234_),
    .Y(net1344));
 sky130_as_sc_hs__buff_2 hold804 (.A(_01072_),
    .Y(net1345));
 sky130_as_sc_hs__buff_2 hold805 (.A(\tholin_riscv.tmr0_pre[16] ),
    .Y(net1346));
 sky130_as_sc_hs__buff_2 hold806 (.A(_17946_),
    .Y(net1347));
 sky130_as_sc_hs__buff_2 hold807 (.A(_17948_),
    .Y(net1348));
 sky130_as_sc_hs__buff_2 hold808 (.A(\tholin_riscv.tmr1_pre[17] ),
    .Y(net1349));
 sky130_as_sc_hs__buff_2 hold809 (.A(_17852_),
    .Y(net1350));
 sky130_as_sc_hs__buff_2 hold81 (.A(_14936_),
    .Y(net622));
 sky130_as_sc_hs__buff_2 hold810 (.A(_17854_),
    .Y(net1351));
 sky130_as_sc_hs__buff_2 hold811 (.A(\tholin_riscv.tmr0_pre[24] ),
    .Y(net1352));
 sky130_as_sc_hs__buff_2 hold812 (.A(_17970_),
    .Y(net1353));
 sky130_as_sc_hs__buff_2 hold813 (.A(_17972_),
    .Y(net1354));
 sky130_as_sc_hs__buff_2 hold814 (.A(\tholin_riscv.tmr0_pre[3] ),
    .Y(net1355));
 sky130_as_sc_hs__buff_2 hold815 (.A(_17908_),
    .Y(net1356));
 sky130_as_sc_hs__buff_2 hold816 (.A(_17910_),
    .Y(net1357));
 sky130_as_sc_hs__buff_2 hold817 (.A(\tholin_riscv.requested_addr[31] ),
    .Y(net1358));
 sky130_as_sc_hs__buff_2 hold818 (.A(_16975_),
    .Y(net1359));
 sky130_as_sc_hs__buff_2 hold819 (.A(_16976_),
    .Y(net1360));
 sky130_as_sc_hs__buff_2 hold82 (.A(_01003_),
    .Y(net623));
 sky130_as_sc_hs__buff_2 hold820 (.A(\tholin_riscv.tmr1_pre[22] ),
    .Y(net1361));
 sky130_as_sc_hs__buff_2 hold821 (.A(_17867_),
    .Y(net1362));
 sky130_as_sc_hs__buff_2 hold822 (.A(_17869_),
    .Y(net1363));
 sky130_as_sc_hs__buff_2 hold823 (.A(\tholin_riscv.tmr0_pre[25] ),
    .Y(net1364));
 sky130_as_sc_hs__buff_2 hold824 (.A(_17973_),
    .Y(net1365));
 sky130_as_sc_hs__buff_2 hold825 (.A(_17975_),
    .Y(net1366));
 sky130_as_sc_hs__buff_2 hold826 (.A(_01497_),
    .Y(net1367));
 sky130_as_sc_hs__buff_2 hold827 (.A(\tholin_riscv.tmr0_pre[28] ),
    .Y(net1368));
 sky130_as_sc_hs__buff_2 hold828 (.A(_17982_),
    .Y(net1369));
 sky130_as_sc_hs__buff_2 hold829 (.A(_17984_),
    .Y(net1370));
 sky130_as_sc_hs__buff_2 hold83 (.A(net1783),
    .Y(net624));
 sky130_as_sc_hs__buff_2 hold830 (.A(\tholin_riscv.tmr0_pre[17] ),
    .Y(net1371));
 sky130_as_sc_hs__buff_2 hold831 (.A(_17949_),
    .Y(net1372));
 sky130_as_sc_hs__buff_2 hold832 (.A(_17951_),
    .Y(net1373));
 sky130_as_sc_hs__clkbuff_4 hold833 (.A(net1793),
    .Y(net1374));
 sky130_as_sc_hs__buff_2 hold834 (.A(_15231_),
    .Y(net1375));
 sky130_as_sc_hs__buff_2 hold835 (.A(\tholin_riscv.tmr1_pre[1] ),
    .Y(net1376));
 sky130_as_sc_hs__buff_2 hold836 (.A(_17805_),
    .Y(net1377));
 sky130_as_sc_hs__buff_2 hold837 (.A(_17807_),
    .Y(net1378));
 sky130_as_sc_hs__buff_2 hold838 (.A(_01441_),
    .Y(net1379));
 sky130_as_sc_hs__buff_2 hold839 (.A(\tholin_riscv.tmr1_pre[18] ),
    .Y(net1380));
 sky130_as_sc_hs__buff_2 hold84 (.A(_15265_),
    .Y(net625));
 sky130_as_sc_hs__buff_2 hold840 (.A(_17855_),
    .Y(net1381));
 sky130_as_sc_hs__buff_2 hold841 (.A(_17857_),
    .Y(net1382));
 sky130_as_sc_hs__buff_2 hold842 (.A(\tholin_riscv.tmr1_pre[14] ),
    .Y(net1383));
 sky130_as_sc_hs__buff_2 hold843 (.A(_17843_),
    .Y(net1384));
 sky130_as_sc_hs__buff_2 hold844 (.A(_17845_),
    .Y(net1385));
 sky130_as_sc_hs__buff_2 hold845 (.A(\tholin_riscv.requested_addr[27] ),
    .Y(net1386));
 sky130_as_sc_hs__buff_2 hold846 (.A(_16951_),
    .Y(net1387));
 sky130_as_sc_hs__buff_2 hold847 (.A(_16952_),
    .Y(net1388));
 sky130_as_sc_hs__buff_2 hold848 (.A(\tholin_riscv.tmr0_pre[23] ),
    .Y(net1389));
 sky130_as_sc_hs__buff_2 hold849 (.A(_17967_),
    .Y(net1390));
 sky130_as_sc_hs__buff_2 hold85 (.A(_01082_),
    .Y(net626));
 sky130_as_sc_hs__buff_2 hold850 (.A(_17969_),
    .Y(net1391));
 sky130_as_sc_hs__buff_2 hold851 (.A(\tholin_riscv.tmr1_pre[2] ),
    .Y(net1392));
 sky130_as_sc_hs__buff_2 hold852 (.A(_17808_),
    .Y(net1393));
 sky130_as_sc_hs__buff_2 hold853 (.A(_17810_),
    .Y(net1394));
 sky130_as_sc_hs__buff_2 hold854 (.A(\tholin_riscv.tmr1_pre[5] ),
    .Y(net1395));
 sky130_as_sc_hs__buff_2 hold855 (.A(_17817_),
    .Y(net1396));
 sky130_as_sc_hs__buff_2 hold856 (.A(_17819_),
    .Y(net1397));
 sky130_as_sc_hs__buff_2 hold857 (.A(\tholin_riscv.requested_addr[11] ),
    .Y(net1398));
 sky130_as_sc_hs__buff_2 hold858 (.A(_16855_),
    .Y(net1399));
 sky130_as_sc_hs__buff_2 hold859 (.A(_16856_),
    .Y(net1400));
 sky130_as_sc_hs__buff_2 hold86 (.A(net1786),
    .Y(net627));
 sky130_as_sc_hs__buff_2 hold860 (.A(\tholin_riscv.requested_addr[18] ),
    .Y(net1401));
 sky130_as_sc_hs__buff_2 hold861 (.A(_16897_),
    .Y(net1402));
 sky130_as_sc_hs__buff_2 hold862 (.A(_16898_),
    .Y(net1403));
 sky130_as_sc_hs__buff_2 hold863 (.A(\tholin_riscv.tmr0_pre[7] ),
    .Y(net1404));
 sky130_as_sc_hs__buff_2 hold864 (.A(_17920_),
    .Y(net1405));
 sky130_as_sc_hs__buff_2 hold865 (.A(_17922_),
    .Y(net1406));
 sky130_as_sc_hs__buff_2 hold866 (.A(_01479_),
    .Y(net1407));
 sky130_as_sc_hs__buff_2 hold867 (.A(\tholin_riscv.intr_vec[23] ),
    .Y(net1408));
 sky130_as_sc_hs__buff_2 hold868 (.A(_17046_),
    .Y(net1409));
 sky130_as_sc_hs__buff_2 hold869 (.A(_17048_),
    .Y(net1410));
 sky130_as_sc_hs__buff_2 hold87 (.A(_15250_),
    .Y(net628));
 sky130_as_sc_hs__buff_2 hold870 (.A(\tholin_riscv.tmr0_pre[10] ),
    .Y(net1411));
 sky130_as_sc_hs__buff_2 hold871 (.A(_17929_),
    .Y(net1412));
 sky130_as_sc_hs__buff_2 hold872 (.A(_17931_),
    .Y(net1413));
 sky130_as_sc_hs__buff_2 hold873 (.A(_01482_),
    .Y(net1414));
 sky130_as_sc_hs__buff_2 hold874 (.A(\tholin_riscv.tmr1_pre[25] ),
    .Y(net1415));
 sky130_as_sc_hs__buff_2 hold875 (.A(_17876_),
    .Y(net1416));
 sky130_as_sc_hs__buff_2 hold876 (.A(_17878_),
    .Y(net1417));
 sky130_as_sc_hs__buff_2 hold877 (.A(_01465_),
    .Y(net1418));
 sky130_as_sc_hs__buff_2 hold878 (.A(\tholin_riscv.tmr1_pre[19] ),
    .Y(net1419));
 sky130_as_sc_hs__buff_2 hold879 (.A(_17858_),
    .Y(net1420));
 sky130_as_sc_hs__buff_2 hold88 (.A(_01077_),
    .Y(net629));
 sky130_as_sc_hs__buff_2 hold880 (.A(_17860_),
    .Y(net1421));
 sky130_as_sc_hs__buff_2 hold881 (.A(\tholin_riscv.tmr0_pre[12] ),
    .Y(net1422));
 sky130_as_sc_hs__buff_2 hold882 (.A(_17935_),
    .Y(net1423));
 sky130_as_sc_hs__buff_2 hold883 (.A(_17937_),
    .Y(net1424));
 sky130_as_sc_hs__buff_2 hold884 (.A(\tholin_riscv.intr_vec[28] ),
    .Y(net1425));
 sky130_as_sc_hs__buff_2 hold885 (.A(_17061_),
    .Y(net1426));
 sky130_as_sc_hs__buff_2 hold886 (.A(_17063_),
    .Y(net1427));
 sky130_as_sc_hs__buff_2 hold887 (.A(\tholin_riscv.instr[6] ),
    .Y(net1428));
 sky130_as_sc_hs__buff_2 hold888 (.A(_21447_),
    .Y(net1429));
 sky130_as_sc_hs__buff_2 hold889 (.A(_00019_),
    .Y(net1430));
 sky130_as_sc_hs__buff_2 hold89 (.A(net1788),
    .Y(net630));
 sky130_as_sc_hs__buff_2 hold890 (.A(\tholin_riscv.tmr1_pre[15] ),
    .Y(net1431));
 sky130_as_sc_hs__buff_2 hold891 (.A(_17846_),
    .Y(net1432));
 sky130_as_sc_hs__buff_2 hold892 (.A(_17848_),
    .Y(net1433));
 sky130_as_sc_hs__buff_2 hold893 (.A(\tholin_riscv.tmr0_pre[30] ),
    .Y(net1434));
 sky130_as_sc_hs__buff_2 hold894 (.A(_17988_),
    .Y(net1435));
 sky130_as_sc_hs__buff_2 hold895 (.A(_17990_),
    .Y(net1436));
 sky130_as_sc_hs__buff_2 hold896 (.A(_01502_),
    .Y(net1437));
 sky130_as_sc_hs__buff_2 hold897 (.A(\tholin_riscv.tmr0_pre[13] ),
    .Y(net1438));
 sky130_as_sc_hs__buff_2 hold898 (.A(_17938_),
    .Y(net1439));
 sky130_as_sc_hs__buff_2 hold899 (.A(_17940_),
    .Y(net1440));
 sky130_as_sc_hs__buff_2 hold9 (.A(_01571_),
    .Y(net550));
 sky130_as_sc_hs__buff_2 hold90 (.A(_15280_),
    .Y(net631));
 sky130_as_sc_hs__buff_2 hold900 (.A(\tholin_riscv.tmr1_pre[27] ),
    .Y(net1441));
 sky130_as_sc_hs__buff_2 hold901 (.A(_17882_),
    .Y(net1442));
 sky130_as_sc_hs__buff_2 hold902 (.A(_17884_),
    .Y(net1443));
 sky130_as_sc_hs__buff_2 hold903 (.A(\tholin_riscv.tmr0_pre[6] ),
    .Y(net1444));
 sky130_as_sc_hs__buff_2 hold904 (.A(_17917_),
    .Y(net1445));
 sky130_as_sc_hs__buff_2 hold905 (.A(_17919_),
    .Y(net1446));
 sky130_as_sc_hs__buff_2 hold906 (.A(\tholin_riscv.tmr0_pre[19] ),
    .Y(net1447));
 sky130_as_sc_hs__buff_2 hold907 (.A(_17955_),
    .Y(net1448));
 sky130_as_sc_hs__buff_2 hold908 (.A(_17957_),
    .Y(net1449));
 sky130_as_sc_hs__buff_2 hold909 (.A(\tholin_riscv.tmr0_pre[4] ),
    .Y(net1450));
 sky130_as_sc_hs__buff_2 hold91 (.A(_01086_),
    .Y(net632));
 sky130_as_sc_hs__buff_2 hold910 (.A(_17911_),
    .Y(net1451));
 sky130_as_sc_hs__buff_2 hold911 (.A(_17913_),
    .Y(net1452));
 sky130_as_sc_hs__buff_2 hold912 (.A(\tholin_riscv.tmr1_pre[24] ),
    .Y(net1453));
 sky130_as_sc_hs__buff_2 hold913 (.A(_17873_),
    .Y(net1454));
 sky130_as_sc_hs__buff_2 hold914 (.A(_17875_),
    .Y(net1455));
 sky130_as_sc_hs__buff_2 hold915 (.A(\tholin_riscv.tmr0_pre[31] ),
    .Y(net1456));
 sky130_as_sc_hs__buff_2 hold916 (.A(_17991_),
    .Y(net1457));
 sky130_as_sc_hs__buff_2 hold917 (.A(_17993_),
    .Y(net1458));
 sky130_as_sc_hs__buff_2 hold918 (.A(\tholin_riscv.tmr1_pre[21] ),
    .Y(net1459));
 sky130_as_sc_hs__buff_2 hold919 (.A(_17864_),
    .Y(net1460));
 sky130_as_sc_hs__buff_2 hold92 (.A(net1787),
    .Y(net633));
 sky130_as_sc_hs__buff_2 hold920 (.A(_17866_),
    .Y(net1461));
 sky130_as_sc_hs__buff_2 hold921 (.A(\tholin_riscv.tmr0_pre[1] ),
    .Y(net1462));
 sky130_as_sc_hs__buff_2 hold922 (.A(_17902_),
    .Y(net1463));
 sky130_as_sc_hs__buff_2 hold923 (.A(_17904_),
    .Y(net1464));
 sky130_as_sc_hs__buff_2 hold924 (.A(_01473_),
    .Y(net1465));
 sky130_as_sc_hs__buff_2 hold925 (.A(\tholin_riscv.tmr0_pre[18] ),
    .Y(net1466));
 sky130_as_sc_hs__buff_2 hold926 (.A(_17952_),
    .Y(net1467));
 sky130_as_sc_hs__buff_2 hold927 (.A(_17954_),
    .Y(net1468));
 sky130_as_sc_hs__buff_2 hold928 (.A(\tholin_riscv.tmr1_pre[30] ),
    .Y(net1469));
 sky130_as_sc_hs__buff_2 hold929 (.A(_17891_),
    .Y(net1470));
 sky130_as_sc_hs__buff_2 hold93 (.A(_15286_),
    .Y(net634));
 sky130_as_sc_hs__buff_2 hold930 (.A(_17893_),
    .Y(net1471));
 sky130_as_sc_hs__buff_2 hold931 (.A(_01470_),
    .Y(net1472));
 sky130_as_sc_hs__buff_2 hold932 (.A(\tholin_riscv.tmr1_pre[3] ),
    .Y(net1473));
 sky130_as_sc_hs__buff_2 hold933 (.A(_17811_),
    .Y(net1474));
 sky130_as_sc_hs__buff_2 hold934 (.A(_17813_),
    .Y(net1475));
 sky130_as_sc_hs__buff_2 hold935 (.A(\tholin_riscv.tmr1_pre[16] ),
    .Y(net1476));
 sky130_as_sc_hs__buff_2 hold936 (.A(_17849_),
    .Y(net1477));
 sky130_as_sc_hs__buff_2 hold937 (.A(_17851_),
    .Y(net1478));
 sky130_as_sc_hs__buff_2 hold938 (.A(\tholin_riscv.tmr1_pre[8] ),
    .Y(net1479));
 sky130_as_sc_hs__buff_2 hold939 (.A(_17826_),
    .Y(net1480));
 sky130_as_sc_hs__buff_2 hold94 (.A(_01089_),
    .Y(net635));
 sky130_as_sc_hs__buff_2 hold940 (.A(_17828_),
    .Y(net1481));
 sky130_as_sc_hs__buff_2 hold941 (.A(_01448_),
    .Y(net1482));
 sky130_as_sc_hs__buff_2 hold942 (.A(\tholin_riscv.requested_addr[14] ),
    .Y(net1483));
 sky130_as_sc_hs__buff_2 hold943 (.A(_16873_),
    .Y(net1484));
 sky130_as_sc_hs__buff_2 hold944 (.A(_16874_),
    .Y(net1485));
 sky130_as_sc_hs__buff_2 hold945 (.A(\tholin_riscv.tmr0_pre[11] ),
    .Y(net1486));
 sky130_as_sc_hs__buff_2 hold946 (.A(_17932_),
    .Y(net1487));
 sky130_as_sc_hs__buff_2 hold947 (.A(_17934_),
    .Y(net1488));
 sky130_as_sc_hs__buff_2 hold948 (.A(_01483_),
    .Y(net1489));
 sky130_as_sc_hs__buff_2 hold949 (.A(\tholin_riscv.tmr1_pre[6] ),
    .Y(net1490));
 sky130_as_sc_hs__buff_2 hold95 (.A(net1784),
    .Y(net636));
 sky130_as_sc_hs__buff_2 hold950 (.A(_17820_),
    .Y(net1491));
 sky130_as_sc_hs__buff_2 hold951 (.A(_17822_),
    .Y(net1492));
 sky130_as_sc_hs__buff_2 hold952 (.A(\tholin_riscv.tmr1_pre[11] ),
    .Y(net1493));
 sky130_as_sc_hs__buff_2 hold953 (.A(_17835_),
    .Y(net1494));
 sky130_as_sc_hs__buff_2 hold954 (.A(_17837_),
    .Y(net1495));
 sky130_as_sc_hs__buff_2 hold955 (.A(\tholin_riscv.uart_int_enable ),
    .Y(net1496));
 sky130_as_sc_hs__buff_2 hold956 (.A(_18589_),
    .Y(net1497));
 sky130_as_sc_hs__buff_2 hold957 (.A(_18591_),
    .Y(net1498));
 sky130_as_sc_hs__buff_2 hold958 (.A(\tholin_riscv.tmr0_pre[2] ),
    .Y(net1499));
 sky130_as_sc_hs__buff_2 hold959 (.A(_17905_),
    .Y(net1500));
 sky130_as_sc_hs__buff_2 hold96 (.A(_15284_),
    .Y(net637));
 sky130_as_sc_hs__buff_2 hold960 (.A(_17907_),
    .Y(net1501));
 sky130_as_sc_hs__buff_2 hold961 (.A(\tholin_riscv.tmr1_pre[31] ),
    .Y(net1502));
 sky130_as_sc_hs__buff_2 hold962 (.A(_17894_),
    .Y(net1503));
 sky130_as_sc_hs__buff_2 hold963 (.A(_17896_),
    .Y(net1504));
 sky130_as_sc_hs__buff_2 hold964 (.A(_01471_),
    .Y(net1505));
 sky130_as_sc_hs__buff_2 hold965 (.A(\tholin_riscv.tmr1_pre[4] ),
    .Y(net1506));
 sky130_as_sc_hs__buff_2 hold966 (.A(_17814_),
    .Y(net1507));
 sky130_as_sc_hs__buff_2 hold967 (.A(_17816_),
    .Y(net1508));
 sky130_as_sc_hs__buff_2 hold968 (.A(\tholin_riscv.tmr1_pre[23] ),
    .Y(net1509));
 sky130_as_sc_hs__buff_2 hold969 (.A(_17870_),
    .Y(net1510));
 sky130_as_sc_hs__buff_2 hold97 (.A(_01088_),
    .Y(net638));
 sky130_as_sc_hs__buff_2 hold970 (.A(_17872_),
    .Y(net1511));
 sky130_as_sc_hs__buff_2 hold971 (.A(\tholin_riscv.requested_addr[23] ),
    .Y(net1512));
 sky130_as_sc_hs__buff_2 hold972 (.A(_16927_),
    .Y(net1513));
 sky130_as_sc_hs__buff_2 hold973 (.A(_16928_),
    .Y(net1514));
 sky130_as_sc_hs__buff_2 hold974 (.A(\tholin_riscv.tmr0_pre[21] ),
    .Y(net1515));
 sky130_as_sc_hs__buff_2 hold975 (.A(_17961_),
    .Y(net1516));
 sky130_as_sc_hs__buff_2 hold976 (.A(_17963_),
    .Y(net1517));
 sky130_as_sc_hs__buff_2 hold977 (.A(\tholin_riscv.requested_addr[22] ),
    .Y(net1518));
 sky130_as_sc_hs__buff_2 hold978 (.A(_16921_),
    .Y(net1519));
 sky130_as_sc_hs__buff_2 hold979 (.A(_16922_),
    .Y(net1520));
 sky130_as_sc_hs__buff_2 hold98 (.A(net1785),
    .Y(net639));
 sky130_as_sc_hs__buff_2 hold980 (.A(\tholin_riscv.tmr0_pre[20] ),
    .Y(net1521));
 sky130_as_sc_hs__buff_2 hold981 (.A(_17958_),
    .Y(net1522));
 sky130_as_sc_hs__buff_2 hold982 (.A(_17960_),
    .Y(net1523));
 sky130_as_sc_hs__buff_2 hold983 (.A(\tholin_riscv.intr_vec[20] ),
    .Y(net1524));
 sky130_as_sc_hs__buff_2 hold984 (.A(_17037_),
    .Y(net1525));
 sky130_as_sc_hs__buff_2 hold985 (.A(\tholin_riscv.tmr1_pre[13] ),
    .Y(net1526));
 sky130_as_sc_hs__buff_2 hold986 (.A(_17840_),
    .Y(net1527));
 sky130_as_sc_hs__buff_2 hold987 (.A(_17842_),
    .Y(net1528));
 sky130_as_sc_hs__buff_2 hold988 (.A(\tholin_riscv.tmr0_pre[14] ),
    .Y(net1529));
 sky130_as_sc_hs__buff_2 hold989 (.A(_17941_),
    .Y(net1530));
 sky130_as_sc_hs__buff_2 hold99 (.A(_16176_),
    .Y(net640));
 sky130_as_sc_hs__buff_2 hold990 (.A(_17943_),
    .Y(net1531));
 sky130_as_sc_hs__buff_2 hold991 (.A(_01486_),
    .Y(net1532));
 sky130_as_sc_hs__buff_2 hold992 (.A(\tholin_riscv.tmr0_pre[27] ),
    .Y(net1533));
 sky130_as_sc_hs__buff_2 hold993 (.A(_17979_),
    .Y(net1534));
 sky130_as_sc_hs__buff_2 hold994 (.A(_17981_),
    .Y(net1535));
 sky130_as_sc_hs__buff_2 hold995 (.A(\tholin_riscv.tmr1_pre[7] ),
    .Y(net1536));
 sky130_as_sc_hs__buff_2 hold996 (.A(_17823_),
    .Y(net1537));
 sky130_as_sc_hs__buff_2 hold997 (.A(_17825_),
    .Y(net1538));
 sky130_as_sc_hs__buff_2 hold998 (.A(\tholin_riscv.intr_vec[14] ),
    .Y(net1539));
 sky130_as_sc_hs__buff_2 hold999 (.A(_17019_),
    .Y(net1540));
 sky130_as_sc_hs__buff_2 input1 (.A(custom_settings[0]),
    .Y(net1));
 sky130_as_sc_hs__buff_2 input10 (.A(io_in[1]),
    .Y(net10));
 sky130_as_sc_hs__buff_2 input11 (.A(io_in[23]),
    .Y(net11));
 sky130_as_sc_hs__clkbuff_8 input12 (.Y(net12),
    .A(io_in[26]));
 sky130_as_sc_hs__buff_2 input13 (.A(io_in[2]),
    .Y(net13));
 sky130_as_sc_hs__clkbuff_8 input14 (.Y(net14),
    .A(io_in[32]));
 sky130_as_sc_hs__buff_2 input15 (.A(io_in[3]),
    .Y(net15));
 sky130_as_sc_hs__buff_2 input16 (.A(io_in[4]),
    .Y(net16));
 sky130_as_sc_hs__buff_2 input17 (.A(io_in[5]),
    .Y(net17));
 sky130_as_sc_hs__buff_2 input18 (.A(io_in[6]),
    .Y(net18));
 sky130_as_sc_hs__buff_2 input19 (.A(io_in[7]),
    .Y(net19));
 sky130_as_sc_hs__buff_2 input2 (.A(custom_settings[1]),
    .Y(net2));
 sky130_as_sc_hs__buff_2 input20 (.A(io_in[8]),
    .Y(net20));
 sky130_as_sc_hs__buff_2 input21 (.A(io_in[9]),
    .Y(net21));
 sky130_as_sc_hs__buff_11 input22 (.A(rst_n),
    .Y(net22));
 sky130_as_sc_hs__buff_2 input3 (.A(io_in[0]),
    .Y(net3));
 sky130_as_sc_hs__buff_2 input4 (.A(io_in[10]),
    .Y(net4));
 sky130_as_sc_hs__clkbuff_4 input5 (.A(io_in[11]),
    .Y(net5));
 sky130_as_sc_hs__buff_2 input6 (.A(io_in[12]),
    .Y(net6));
 sky130_as_sc_hs__buff_2 input7 (.A(io_in[13]),
    .Y(net7));
 sky130_as_sc_hs__clkbuff_4 input8 (.A(io_in[14]),
    .Y(net8));
 sky130_as_sc_hs__clkbuff_4 input9 (.A(io_in[15]),
    .Y(net9));
 sky130_as_sc_hs__clkbuff_11 output23 (.A(net23),
    .Y(io_oeb[0]));
 sky130_as_sc_hs__clkbuff_11 output24 (.A(net24),
    .Y(io_oeb[10]));
 sky130_as_sc_hs__clkbuff_11 output25 (.A(net25),
    .Y(io_oeb[11]));
 sky130_as_sc_hs__clkbuff_11 output26 (.A(net26),
    .Y(io_oeb[12]));
 sky130_as_sc_hs__clkbuff_11 output27 (.A(net27),
    .Y(io_oeb[13]));
 sky130_as_sc_hs__clkbuff_11 output28 (.A(net28),
    .Y(io_oeb[14]));
 sky130_as_sc_hs__clkbuff_11 output29 (.A(net29),
    .Y(io_oeb[15]));
 sky130_as_sc_hs__clkbuff_11 output30 (.A(net30),
    .Y(io_oeb[1]));
 sky130_as_sc_hs__clkbuff_11 output31 (.A(net31),
    .Y(io_oeb[27]));
 sky130_as_sc_hs__clkbuff_11 output32 (.A(net32),
    .Y(io_oeb[28]));
 sky130_as_sc_hs__clkbuff_11 output33 (.A(net33),
    .Y(io_oeb[29]));
 sky130_as_sc_hs__clkbuff_11 output34 (.A(net34),
    .Y(io_oeb[2]));
 sky130_as_sc_hs__clkbuff_11 output35 (.A(net35),
    .Y(io_oeb[30]));
 sky130_as_sc_hs__clkbuff_11 output36 (.A(net36),
    .Y(io_oeb[31]));
 sky130_as_sc_hs__clkbuff_11 output37 (.A(net37),
    .Y(io_oeb[32]));
 sky130_as_sc_hs__clkbuff_11 output38 (.A(net38),
    .Y(io_oeb[3]));
 sky130_as_sc_hs__clkbuff_11 output39 (.A(net39),
    .Y(io_oeb[4]));
 sky130_as_sc_hs__clkbuff_11 output40 (.A(net40),
    .Y(io_oeb[5]));
 sky130_as_sc_hs__clkbuff_11 output41 (.A(net41),
    .Y(io_oeb[6]));
 sky130_as_sc_hs__clkbuff_11 output42 (.A(net42),
    .Y(io_oeb[7]));
 sky130_as_sc_hs__clkbuff_11 output43 (.A(net43),
    .Y(io_oeb[8]));
 sky130_as_sc_hs__clkbuff_11 output44 (.A(net44),
    .Y(io_oeb[9]));
 sky130_as_sc_hs__clkbuff_11 output45 (.A(net45),
    .Y(io_out[0]));
 sky130_as_sc_hs__clkbuff_11 output46 (.A(net46),
    .Y(io_out[10]));
 sky130_as_sc_hs__clkbuff_11 output47 (.A(net47),
    .Y(io_out[11]));
 sky130_as_sc_hs__clkbuff_11 output48 (.A(net48),
    .Y(io_out[12]));
 sky130_as_sc_hs__clkbuff_11 output49 (.A(net49),
    .Y(io_out[13]));
 sky130_as_sc_hs__clkbuff_11 output50 (.A(net50),
    .Y(io_out[14]));
 sky130_as_sc_hs__clkbuff_11 output51 (.A(net51),
    .Y(io_out[15]));
 sky130_as_sc_hs__buff_2 output52 (.A(net52),
    .Y(io_out[16]));
 sky130_as_sc_hs__buff_2 output53 (.A(net53),
    .Y(io_out[17]));
 sky130_as_sc_hs__clkbuff_11 output54 (.A(net54),
    .Y(io_out[18]));
 sky130_as_sc_hs__clkbuff_11 output55 (.A(net55),
    .Y(io_out[19]));
 sky130_as_sc_hs__clkbuff_11 output56 (.A(net56),
    .Y(io_out[1]));
 sky130_as_sc_hs__clkbuff_11 output57 (.A(net57),
    .Y(io_out[22]));
 sky130_as_sc_hs__clkbuff_11 output58 (.A(net58),
    .Y(io_out[24]));
 sky130_as_sc_hs__clkbuff_11 output59 (.A(net59),
    .Y(io_out[25]));
 sky130_as_sc_hs__clkbuff_11 output60 (.A(net60),
    .Y(io_out[27]));
 sky130_as_sc_hs__clkbuff_11 output61 (.A(net61),
    .Y(io_out[28]));
 sky130_as_sc_hs__clkbuff_11 output62 (.A(net62),
    .Y(io_out[29]));
 sky130_as_sc_hs__clkbuff_11 output63 (.A(net63),
    .Y(io_out[2]));
 sky130_as_sc_hs__clkbuff_11 output64 (.A(net64),
    .Y(io_out[30]));
 sky130_as_sc_hs__clkbuff_11 output65 (.A(net65),
    .Y(io_out[31]));
 sky130_as_sc_hs__clkbuff_11 output66 (.A(net66),
    .Y(io_out[32]));
 sky130_as_sc_hs__clkbuff_11 output67 (.A(net67),
    .Y(io_out[3]));
 sky130_as_sc_hs__clkbuff_11 output68 (.A(net68),
    .Y(io_out[4]));
 sky130_as_sc_hs__clkbuff_11 output69 (.A(net69),
    .Y(io_out[5]));
 sky130_as_sc_hs__clkbuff_11 output70 (.A(net70),
    .Y(io_out[6]));
 sky130_as_sc_hs__clkbuff_11 output71 (.A(net71),
    .Y(io_out[7]));
 sky130_as_sc_hs__clkbuff_11 output72 (.A(net72),
    .Y(io_out[8]));
 sky130_as_sc_hs__clkbuff_11 output73 (.A(net73),
    .Y(io_out[9]));
 sky130_as_sc_hs__tiel wrapped_tholin_riscv_528 (.ZERO(net528));
 sky130_as_sc_hs__tiel wrapped_tholin_riscv_529 (.ZERO(net529));
 sky130_as_sc_hs__tiel wrapped_tholin_riscv_530 (.ZERO(net530));
 sky130_as_sc_hs__tiel wrapped_tholin_riscv_531 (.ZERO(net531));
 sky130_as_sc_hs__tiel wrapped_tholin_riscv_532 (.ZERO(net532));
 sky130_as_sc_hs__tiel wrapped_tholin_riscv_533 (.ZERO(net533));
 sky130_as_sc_hs__tiel wrapped_tholin_riscv_534 (.ZERO(net534));
 sky130_as_sc_hs__tiel wrapped_tholin_riscv_535 (.ZERO(net535));
 sky130_as_sc_hs__tiel wrapped_tholin_riscv_536 (.ZERO(net536));
 sky130_as_sc_hs__tiel wrapped_tholin_riscv_537 (.ZERO(net537));
 sky130_as_sc_hs__tiel wrapped_tholin_riscv_538 (.ZERO(net538));
 sky130_as_sc_hs__tieh wrapped_tholin_riscv_539 (.ONE(net539));
 sky130_as_sc_hs__tieh wrapped_tholin_riscv_540 (.ONE(net540));
 sky130_as_sc_hs__tieh wrapped_tholin_riscv_541 (.ONE(net541));
 assign io_oeb[16] = net528;
 assign io_oeb[17] = net529;
 assign io_oeb[18] = net530;
 assign io_oeb[19] = net531;
 assign io_oeb[20] = net532;
 assign io_oeb[21] = net533;
 assign io_oeb[22] = net534;
 assign io_oeb[23] = net539;
 assign io_oeb[24] = net535;
 assign io_oeb[25] = net536;
 assign io_oeb[26] = net540;
 assign io_oeb[33] = net541;
 assign io_out[23] = net537;
 assign io_out[26] = net538;
endmodule

